
// 	Thu Dec 22 20:07:40 2022
//	vlsi
//	192.168.126.129

module datapath__0_131 (opt_ipoPP_0, opt_ipoPP_2, B_in, p_0);

output [31:0] p_0;
input [31:0] B_in;
input opt_ipoPP_0;
input opt_ipoPP_2;
wire n_0;
wire n_4;
wire n_1;
wire n_2;
wire n_3;
wire n_7;
wire n_137;
wire n_138;
wire n_5;
wire n_6;
wire n_136;
wire n_110;
wire n_8;
wire n_9;
wire n_17;
wire n_133;
wire n_10;
wire n_14;
wire n_11;
wire n_16;
wire n_13;
wire n_12;
wire n_15;
wire n_134;
wire n_18;
wire n_130;
wire n_126;
wire n_19;
wire n_20;
wire n_22;
wire n_21;
wire n_124;
wire n_127;
wire n_23;
wire n_24;
wire n_120;
wire n_25;
wire n_27;
wire n_26;
wire n_30;
wire n_84;
wire n_121;
wire CLOCK_slo__n776;
wire n_28;
wire n_87;
wire n_86;
wire n_31;
wire n_81;
wire n_129;
wire n_33;
wire n_34;
wire n_36;
wire n_80;
wire n_106;
wire n_35;
wire n_40;
wire n_107;
wire n_37;
wire n_116;
wire n_38;
wire slo__n517;
wire n_39;
wire n_46;
wire n_42;
wire n_43;
wire n_44;
wire n_109;
wire n_108;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_105;
wire n_51;
wire n_113;
wire opt_ipo_n562;
wire n_52;
wire n_55;
wire n_53;
wire n_54;
wire n_114;
wire n_56;
wire n_62;
wire n_112;
wire n_57;
wire n_59;
wire n_58;
wire n_63;
wire n_60;
wire n_100;
wire n_76;
wire n_61;
wire n_65;
wire n_67;
wire n_74;
wire n_64;
wire n_66;
wire n_102;
wire n_68;
wire n_101;
wire n_69;
wire n_70;
wire n_94;
wire n_96;
wire n_71;
wire n_73;
wire n_72;
wire n_91;
wire n_93;
wire n_75;
wire n_98;
wire n_77;
wire n_115;
wire n_78;
wire n_89;
wire n_79;
wire n_88;
wire slo__mro_n111;
wire n_123;
wire n_85;
wire n_122;
wire n_131;
wire n_90;
wire n_92;
wire n_95;
wire n_97;
wire n_99;
wire n_103;
wire n_117;
wire n_119;
wire CLOCK_slo__n1165;
wire n_128;
wire n_132;
wire n_111;
wire slo__mro_n109;
wire CLOCK_slo__n753;
wire sgo__sro_n10;
wire slo__mro_n110;
wire sgo__sro_n35;
wire sgo__sro_n36;
wire slo__xsl_n355;
wire slo__n341;
wire opt_ipo_n613;
wire slo__n207;
wire slo__n168;
wire CLOCK_slo__sro_n764;
wire slo__n422;
wire slo__n326;
wire slo__n549;
wire slo__xsl_n489;
wire slo__sro_n433;
wire slo__sro_n434;
wire opt_ipo_n596;
wire opt_ipo_n599;
wire opt_ipo_n575;
wire CLOCK_slo__xsl_n931;


INV_X1 i_169 (.ZN (n_114), .A (opt_ipoPP_0));
INV_X1 i_168 (.ZN (n_113), .A (B_in[20]));
NOR3_X2 i_167 (.ZN (n_112), .A1 (B_in[22]), .A2 (B_in[20]), .A3 (B_in[21]));
INV_X2 i_166 (.ZN (n_111), .A (B_in[3]));
INV_X4 i_165 (.ZN (n_110), .A (B_in[2]));
INV_X1 i_164 (.ZN (n_138), .A (B_in[1]));
INV_X1 i_163 (.ZN (n_137), .A (B_in[0]));
NAND2_X2 CLOCK_slo__c1304 (.ZN (CLOCK_slo__n1165), .A1 (opt_ipo_n575), .A2 (slo__n207));
NAND3_X4 CLOCK_slo__sro_c848 (.ZN (CLOCK_slo__sro_n764), .A1 (n_128), .A2 (slo__n326), .A3 (n_127));
INV_X2 i_160 (.ZN (n_134), .A (B_in[6]));
INV_X2 i_159 (.ZN (n_133), .A (B_in[5]));
INV_X4 i_158 (.ZN (n_132), .A (B_in[4]));
INV_X4 slo__mro_c165 (.ZN (slo__mro_n111), .A (n_136));
INV_X2 i_155 (.ZN (n_129), .A (B_in[15]));
INV_X1 i_154 (.ZN (n_128), .A (B_in[10]));
INV_X2 i_153 (.ZN (n_127), .A (B_in[9]));
INV_X1 i_152 (.ZN (n_126), .A (B_in[8]));
INV_X4 i_150 (.ZN (n_124), .A (CLOCK_slo__sro_n764));
INV_X2 i_149 (.ZN (n_123), .A (B_in[14]));
INV_X2 i_148 (.ZN (n_122), .A (B_in[13]));
INV_X4 i_147 (.ZN (n_121), .A (B_in[12]));
INV_X2 i_146 (.ZN (n_120), .A (B_in[11]));
INV_X2 CLOCK_slo__c863 (.ZN (CLOCK_slo__n776), .A (n_117));
INV_X2 opt_ipo_c642 (.ZN (opt_ipo_n562), .A (n_33));
NAND3_X4 i_143 (.ZN (n_117), .A1 (n_119), .A2 (n_129), .A3 (CLOCK_slo__n753));
INV_X4 i_142 (.ZN (n_116), .A (n_117));
INV_X1 i_141 (.ZN (n_115), .A (B_in[23]));
INV_X1 i_140 (.ZN (n_109), .A (B_in[19]));
INV_X1 i_139 (.ZN (n_108), .A (B_in[18]));
INV_X1 i_138 (.ZN (n_107), .A (B_in[17]));
INV_X1 i_137 (.ZN (n_106), .A (B_in[16]));
INV_X1 opt_ipo_c673 (.ZN (opt_ipo_n599), .A (n_42));
INV_X1 opt_ipo_c671 (.ZN (opt_ipo_n596), .A (opt_ipoPP_2));
INV_X1 i_134 (.ZN (n_103), .A (B_in[27]));
INV_X1 i_133 (.ZN (n_102), .A (B_in[26]));
INV_X1 i_132 (.ZN (n_101), .A (B_in[25]));
INV_X1 i_131 (.ZN (n_100), .A (B_in[24]));
NAND4_X1 i_130 (.ZN (n_99), .A1 (n_103), .A2 (n_102), .A3 (n_101), .A4 (n_100));
INV_X1 i_129 (.ZN (n_98), .A (n_99));
NAND4_X1 i_128 (.ZN (n_97), .A1 (n_105), .A2 (n_98), .A3 (n_115), .A4 (n_112));
INV_X1 i_127 (.ZN (n_96), .A (n_97));
INV_X1 i_126 (.ZN (n_95), .A (B_in[29]));
INV_X1 i_125 (.ZN (n_94), .A (B_in[28]));
NAND2_X1 i_124 (.ZN (n_93), .A1 (n_95), .A2 (n_94));
OR2_X1 i_123 (.ZN (n_92), .A1 (n_93), .A2 (B_in[30]));
INV_X1 i_122 (.ZN (n_91), .A (n_92));
NAND4_X1 i_121 (.ZN (n_90), .A1 (n_96), .A2 (n_130), .A3 (n_116), .A4 (n_91));
NAND2_X1 i_120 (.ZN (n_89), .A1 (n_90), .A2 (B_in[31]));
INV_X1 i_119 (.ZN (n_88), .A (B_in[31]));
INV_X4 i_118 (.ZN (n_87), .A (CLOCK_slo__n1165));
INV_X4 i_117 (.ZN (n_86), .A (n_131));
NAND2_X2 i_116 (.ZN (n_85), .A1 (n_122), .A2 (n_121));
INV_X4 i_115 (.ZN (n_84), .A (n_85));
AND4_X4 slo__xsl_c576 (.ZN (n_105), .A1 (n_108), .A2 (n_109), .A3 (slo__n517), .A4 (n_107));
NAND4_X4 i_112 (.ZN (n_81), .A1 (sgo__sro_n35), .A2 (n_87), .A3 (n_86), .A4 (n_124));
INV_X4 i_111 (.ZN (n_80), .A (n_81));
NAND4_X1 i_110 (.ZN (n_79), .A1 (n_80), .A2 (n_88), .A3 (n_96), .A4 (n_91));
NAND2_X1 i_109 (.ZN (n_78), .A1 (n_89), .A2 (n_79));
INV_X1 i_108 (.ZN (p_0[31]), .A (n_78));
NAND3_X4 i_107 (.ZN (n_77), .A1 (n_105), .A2 (n_115), .A3 (slo__n549));
INV_X4 i_106 (.ZN (n_76), .A (n_77));
NAND4_X1 i_105 (.ZN (n_75), .A1 (n_130), .A2 (n_116), .A3 (n_76), .A4 (n_98));
INV_X2 i_104 (.ZN (n_74), .A (n_75));
INV_X1 i_103 (.ZN (n_73), .A (n_93));
NAND4_X1 i_102 (.ZN (n_72), .A1 (n_96), .A2 (n_130), .A3 (n_116), .A4 (n_73));
AOI22_X1 i_101 (.ZN (p_0[30]), .A1 (n_72), .A2 (B_in[30]), .B1 (n_74), .B2 (n_91));
NAND4_X1 i_100 (.ZN (n_71), .A1 (n_96), .A2 (n_130), .A3 (n_94), .A4 (n_116));
AOI22_X1 i_99 (.ZN (p_0[29]), .A1 (n_71), .A2 (B_in[29]), .B1 (n_74), .B2 (n_73));
INV_X1 i_98 (.ZN (n_70), .A (n_71));
AND4_X4 slo__c539 (.ZN (n_119), .A1 (n_123), .A2 (n_121), .A3 (n_122), .A4 (slo__n341));
NOR2_X1 i_96 (.ZN (p_0[28]), .A1 (n_69), .A2 (n_70));
NAND2_X1 i_95 (.ZN (n_68), .A1 (n_101), .A2 (n_100));
INV_X1 i_94 (.ZN (n_67), .A (n_68));
NAND2_X1 i_93 (.ZN (n_66), .A1 (n_67), .A2 (n_102));
INV_X1 i_92 (.ZN (n_65), .A (n_66));
NAND3_X1 i_91 (.ZN (n_64), .A1 (n_80), .A2 (n_76), .A3 (n_65));
AOI21_X1 i_90 (.ZN (p_0[27]), .A (n_74), .B1 (n_64), .B2 (B_in[27]));
NAND3_X1 i_89 (.ZN (n_63), .A1 (n_130), .A2 (n_116), .A3 (n_76));
INV_X1 i_88 (.ZN (n_62), .A (n_63));
NAND4_X1 i_87 (.ZN (n_61), .A1 (n_130), .A2 (n_116), .A3 (n_76), .A4 (n_67));
AOI22_X1 i_86 (.ZN (p_0[26]), .A1 (n_61), .A2 (B_in[26]), .B1 (n_65), .B2 (n_62));
INV_X1 i_85 (.ZN (n_60), .A (n_61));
NAND3_X2 i_84 (.ZN (n_59), .A1 (n_80), .A2 (n_100), .A3 (n_76));
AOI21_X2 i_83 (.ZN (p_0[25]), .A (n_60), .B1 (n_59), .B2 (B_in[25]));
NAND2_X1 i_82 (.ZN (n_58), .A1 (n_63), .A2 (B_in[24]));
NAND2_X1 i_81 (.ZN (n_57), .A1 (n_59), .A2 (n_58));
INV_X1 i_80 (.ZN (p_0[24]), .A (n_57));
NAND3_X1 i_79 (.ZN (n_56), .A1 (n_80), .A2 (n_112), .A3 (n_105));
AOI21_X1 i_78 (.ZN (p_0[23]), .A (n_62), .B1 (n_56), .B2 (B_in[23]));
INV_X1 i_77 (.ZN (n_55), .A (n_56));
NAND2_X1 i_76 (.ZN (n_54), .A1 (n_114), .A2 (n_113));
INV_X1 i_75 (.ZN (n_53), .A (n_54));
NAND4_X2 i_74 (.ZN (n_52), .A1 (n_130), .A2 (CLOCK_slo__n776), .A3 (n_53), .A4 (n_105));
AOI21_X1 i_73 (.ZN (p_0[22]), .A (n_55), .B1 (B_in[22]), .B2 (n_52));
INV_X1 i_72 (.ZN (n_51), .A (n_52));
NAND3_X2 i_71 (.ZN (n_50), .A1 (n_80), .A2 (n_113), .A3 (n_105));
AOI21_X2 i_70 (.ZN (p_0[21]), .A (n_51), .B1 (n_50), .B2 (opt_ipoPP_0));
OAI21_X1 i_69 (.ZN (n_49), .A (B_in[20]), .B1 (opt_ipo_n613), .B2 (slo__xsl_n489));
NAND2_X1 i_68 (.ZN (n_48), .A1 (n_49), .A2 (n_50));
INV_X1 i_67 (.ZN (p_0[20]), .A (n_48));
NAND2_X1 i_66 (.ZN (n_47), .A1 (n_107), .A2 (n_106));
INV_X1 i_65 (.ZN (n_46), .A (n_47));
INV_X1 slo__xsl_c573 (.ZN (slo__xsl_n489), .A (n_105));
NAND2_X1 i_63 (.ZN (n_44), .A1 (n_109), .A2 (n_108));
INV_X1 i_62 (.ZN (n_43), .A (n_44));
NAND4_X4 i_61 (.ZN (n_42), .A1 (n_130), .A2 (n_116), .A3 (n_46), .A4 (n_43));
AOI21_X1 i_59 (.ZN (p_0[19]), .A (opt_ipo_n599), .B1 (slo__sro_n433), .B2 (B_in[19]));
NAND3_X1 i_58 (.ZN (n_40), .A1 (n_130), .A2 (CLOCK_slo__n776), .A3 (n_46));
NAND2_X1 i_57 (.ZN (n_39), .A1 (n_40), .A2 (B_in[18]));
NAND2_X1 i_56 (.ZN (n_38), .A1 (n_39), .A2 (slo__sro_n433));
INV_X1 i_55 (.ZN (p_0[18]), .A (n_38));
NAND3_X1 i_54 (.ZN (n_37), .A1 (n_130), .A2 (n_106), .A3 (CLOCK_slo__n776));
INV_X1 i_53 (.ZN (n_36), .A (n_37));
OAI21_X1 i_52 (.ZN (n_35), .A (n_40), .B1 (n_36), .B2 (n_107));
INV_X1 i_51 (.ZN (p_0[17]), .A (n_35));
NOR2_X1 i_50 (.ZN (n_34), .A1 (n_80), .A2 (n_106));
NOR2_X1 i_49 (.ZN (p_0[16]), .A1 (n_34), .A2 (n_36));
NAND3_X2 i_48 (.ZN (n_33), .A1 (n_130), .A2 (n_124), .A3 (n_119));
AND3_X4 CLOCK_slo__c1109 (.ZN (sgo__sro_n35), .A1 (n_84), .A2 (sgo__sro_n36), .A3 (n_129));
OAI21_X1 i_46 (.ZN (n_31), .A (opt_ipo_n613), .B1 (opt_ipo_n562), .B2 (n_129));
INV_X1 i_45 (.ZN (p_0[15]), .A (n_31));
NAND2_X1 i_42 (.ZN (n_28), .A1 (n_30), .A2 (n_84));
AOI21_X1 i_41 (.ZN (p_0[14]), .A (opt_ipo_n562), .B1 (n_28), .B2 (B_in[14]));
NAND2_X2 i_40 (.ZN (n_27), .A1 (n_30), .A2 (n_121));
AOI22_X1 i_39 (.ZN (p_0[13]), .A1 (n_27), .A2 (B_in[13]), .B1 (n_84), .B2 (n_30));
NAND2_X1 i_38 (.ZN (n_26), .A1 (CLOCK_slo__xsl_n931), .A2 (B_in[12]));
NAND2_X1 i_37 (.ZN (n_25), .A1 (n_27), .A2 (n_26));
INV_X1 i_36 (.ZN (p_0[12]), .A (n_25));
AOI21_X1 i_35 (.ZN (n_24), .A (n_120), .B1 (n_130), .B2 (n_124));
OR2_X1 i_34 (.ZN (n_23), .A1 (n_24), .A2 (n_30));
INV_X1 i_33 (.ZN (p_0[11]), .A (n_23));
NAND3_X2 i_32 (.ZN (n_22), .A1 (n_130), .A2 (n_127), .A3 (n_126));
AOI22_X2 i_31 (.ZN (p_0[10]), .A1 (n_22), .A2 (B_in[10]), .B1 (n_130), .B2 (n_124));
NAND2_X1 i_30 (.ZN (n_21), .A1 (n_130), .A2 (n_126));
NAND2_X1 i_29 (.ZN (n_20), .A1 (n_21), .A2 (B_in[9]));
NAND2_X1 i_28 (.ZN (n_19), .A1 (n_20), .A2 (n_22));
INV_X1 i_27 (.ZN (p_0[9]), .A (n_19));
XNOR2_X1 i_26 (.ZN (n_18), .A (n_130), .B (n_126));
INV_X1 i_25 (.ZN (p_0[8]), .A (n_18));
NOR2_X2 i_24 (.ZN (n_17), .A1 (n_136), .A2 (B_in[4]));
NAND2_X1 i_23 (.ZN (n_16), .A1 (n_17), .A2 (n_133));
INV_X1 i_22 (.ZN (n_15), .A (n_16));
NAND2_X1 i_21 (.ZN (n_14), .A1 (n_15), .A2 (n_134));
NAND2_X1 i_20 (.ZN (n_13), .A1 (n_14), .A2 (opt_ipo_n596));
NAND3_X1 i_19 (.ZN (n_12), .A1 (n_15), .A2 (opt_ipoPP_2), .A3 (n_134));
NAND2_X1 i_18 (.ZN (p_0[7]), .A1 (n_13), .A2 (n_12));
NAND2_X1 i_17 (.ZN (n_11), .A1 (n_16), .A2 (B_in[6]));
NAND2_X1 i_16 (.ZN (n_10), .A1 (n_14), .A2 (n_11));
INV_X1 i_15 (.ZN (p_0[6]), .A (n_10));
XNOR2_X1 i_14 (.ZN (n_9), .A (n_17), .B (n_133));
INV_X1 i_13 (.ZN (p_0[5]), .A (n_9));
XNOR2_X1 i_12 (.ZN (n_8), .A (n_136), .B (B_in[4]));
INV_X1 i_11 (.ZN (p_0[4]), .A (n_8));
NAND3_X1 i_10 (.ZN (n_7), .A1 (n_137), .A2 (n_110), .A3 (n_138));
NAND2_X1 i_9 (.ZN (n_6), .A1 (n_7), .A2 (B_in[3]));
NAND2_X1 i_8 (.ZN (n_5), .A1 (n_6), .A2 (n_136));
INV_X1 i_7 (.ZN (p_0[3]), .A (n_5));
NAND2_X1 i_6 (.ZN (n_4), .A1 (n_137), .A2 (n_138));
NAND2_X1 i_5 (.ZN (n_3), .A1 (n_4), .A2 (B_in[2]));
NAND2_X1 i_4 (.ZN (n_2), .A1 (n_3), .A2 (n_7));
INV_X1 i_3 (.ZN (p_0[2]), .A (n_2));
NAND2_X1 i_2 (.ZN (n_1), .A1 (B_in[0]), .A2 (B_in[1]));
NAND2_X1 i_1 (.ZN (n_0), .A1 (n_4), .A2 (n_1));
INV_X1 i_0 (.ZN (p_0[1]), .A (n_0));
INV_X1 slo__xsl_c406 (.ZN (slo__xsl_n355), .A (n_81));
INV_X8 sgo__c5 (.ZN (n_130), .A (slo__mro_n109));
INV_X2 slo__mro_c166 (.ZN (slo__mro_n110), .A (n_131));
NAND2_X4 slo__mro_c167 (.ZN (slo__mro_n109), .A1 (slo__mro_n111), .A2 (slo__mro_n110));
NAND3_X4 sgo__sro_c16 (.ZN (sgo__sro_n10), .A1 (slo__n168), .A2 (n_110), .A3 (n_111));
INV_X2 CLOCK_slo__c834 (.ZN (CLOCK_slo__n753), .A (CLOCK_slo__sro_n764));
NAND2_X4 sgo__sro_c18 (.ZN (n_136), .A1 (opt_ipo_n575), .A2 (slo__n207));
INV_X1 slo__c386 (.ZN (slo__n341), .A (B_in[11]));
AND2_X2 sgo__sro_c64 (.ZN (sgo__sro_n36), .A1 (n_123), .A2 (n_120));
AOI21_X1 slo__sro_c391 (.ZN (n_69), .A (n_94), .B1 (slo__n422), .B2 (n_96));
INV_X4 slo__c230 (.ZN (slo__n168), .A (B_in[1]));
INV_X1 slo__c273 (.ZN (slo__n207), .A (B_in[0]));
NOR3_X2 slo__c634 (.ZN (slo__n549), .A1 (B_in[22]), .A2 (B_in[20]), .A3 (B_in[21]));
INV_X2 slo__c484 (.ZN (slo__n422), .A (n_81));
INV_X1 slo__c370 (.ZN (slo__n326), .A (B_in[8]));
INV_X1 opt_ipo_c684 (.ZN (opt_ipo_n613), .A (slo__xsl_n355));
INV_X1 slo__c611 (.ZN (slo__n517), .A (B_in[16]));
AND2_X1 slo__sro_c498 (.ZN (slo__sro_n434), .A1 (n_46), .A2 (n_108));
NAND2_X2 slo__sro_c499 (.ZN (slo__sro_n433), .A1 (slo__n422), .A2 (slo__sro_n434));
NAND4_X4 CLOCK_slo__sro_c888 (.ZN (n_131), .A1 (n_134), .A2 (n_132), .A3 (B_in[7]), .A4 (n_133));
INV_X4 opt_ipo_c655 (.ZN (opt_ipo_n575), .A (sgo__sro_n10));
INV_X1 CLOCK_slo__xsl_c1022 (.ZN (CLOCK_slo__xsl_n931), .A (n_30));
AND4_X4 CLOCK_slo__xsl_c1025 (.ZN (n_30), .A1 (n_87), .A2 (n_124), .A3 (n_86), .A4 (n_120));

endmodule //datapath__0_131

module datapath__0_129 (opt_ipoPP_2, A_in, p_0);

output [31:0] p_0;
input [31:0] A_in;
input opt_ipoPP_2;
wire CLOCK_slo__sro_n2198;
wire CLOCK_slo__sro_n1730;
wire CLOCK_sgo__sro_n1460;
wire CLOCK_slo__sro_n2502;
wire CLOCK_slo__n2461;
wire n_0;
wire n_4;
wire n_1;
wire n_2;
wire n_3;
wire n_7;
wire n_74;
wire n_87;
wire n_5;
wire n_6;
wire n_73;
wire n_88;
wire n_9;
wire n_17;
wire n_130;
wire n_10;
wire n_14;
wire n_11;
wire n_16;
wire n_13;
wire n_12;
wire n_15;
wire n_131;
wire n_71;
wire n_28;
wire n_123;
wire n_18;
wire n_19;
wire n_26;
wire n_24;
wire n_21;
wire CLOCK_slo__sro_n2199;
wire n_22;
wire n_25;
wire n_125;
wire n_126;
wire n_27;
wire n_124;
wire n_72;
wire n_127;
wire n_29;
wire n_36;
wire n_30;
wire n_63;
wire n_31;
wire n_33;
wire n_32;
wire n_35;
wire n_118;
wire n_34;
wire n_38;
wire n_119;
wire n_117;
wire n_37;
wire n_39;
wire slo__n960;
wire n_120;
wire CLOCK_slo__sro_n2263;
wire n_45;
wire CLOCK_slo__sro_n1977;
wire n_114;
wire CLOCK_slo__n1960;
wire n_44;
wire n_111;
wire n_109;
wire n_113;
wire n_110;
wire n_46;
wire n_49;
wire n_48;
wire n_47;
wire n_106;
wire slo__n660;
wire n_107;
wire n_50;
wire CLOCK_slo__n2408;
wire n_103;
wire n_52;
wire n_99;
wire n_102;
wire n_53;
wire n_57;
wire n_54;
wire n_55;
wire n_100;
wire n_56;
wire n_58;
wire n_59;
wire n_112;
wire sgo__sro_n151;
wire CLOCK_slo__sro_n2072;
wire n_61;
wire n_98;
wire n_121;
wire n_64;
wire n_65;
wire n_94;
wire sgo__sro_n195;
wire n_66;
wire n_93;
wire n_67;
wire n_92;
wire n_69;
wire n_81;
wire n_70;
wire n_76;
wire n_105;
wire n_77;
wire n_78;
wire n_80;
wire n_89;
wire n_97;
wire n_90;
wire n_82;
wire n_85;
wire n_83;
wire n_84;
wire n_86;
wire n_101;
wire n_116;
wire n_122;
wire slo__n428;
wire n_129;
wire n_91;
wire n_95;
wire n_96;
wire n_104;
wire slo__n602;
wire sgo__sro_n150;
wire sgo__sro_n196;
wire sgo__sro_n197;
wire CLOCK_sgo__sro_n1461;
wire slo__xsl_n580;
wire slo__n900;
wire slo__n967;
wire slo__n554;
wire slo__n648;
wire slo__n1020;
wire CLOCK_slo__sro_n1932;
wire opt_ipo_n1163;
wire CLOCK_sgo__sro_n1459;
wire slo__sro_n1043;
wire CLOCK_slo__sro_n1729;
wire CLOCK_slo__mro_n1619;
wire slo__n760;
wire opt_ipo_n1185;
wire CLOCK_slo__n1914;
wire CLOCK_slo__mro_n2257;
wire CLOCK_slo__sro_n2264;
wire CLOCK_slo__sro_n2265;
wire CLOCK_slo__n2694;
wire CLOCK_slo__sro_n2595;


INV_X1 i_161 (.ZN (n_107), .A (A_in[19]));
INV_X1 i_160 (.ZN (n_106), .A (A_in[18]));
NOR2_X4 i_159 (.ZN (n_105), .A1 (A_in[19]), .A2 (A_in[18]));
INV_X1 i_158 (.ZN (n_104), .A (A_in[27]));
NAND3_X1 CLOCK_slo__sro_c3127 (.ZN (n_67), .A1 (n_113), .A2 (n_76), .A3 (n_93));
INV_X1 i_156 (.ZN (n_100), .A (A_in[21]));
INV_X1 i_155 (.ZN (n_99), .A (A_in[20]));
NOR3_X4 i_154 (.ZN (n_98), .A1 (A_in[22]), .A2 (A_in[20]), .A3 (A_in[21]));
NOR2_X1 i_153 (.ZN (n_97), .A1 (A_in[29]), .A2 (A_in[28]));
INV_X1 i_152 (.ZN (n_96), .A (A_in[26]));
INV_X1 i_151 (.ZN (n_95), .A (A_in[25]));
INV_X1 i_150 (.ZN (n_94), .A (A_in[24]));
NOR2_X1 i_149 (.ZN (n_93), .A1 (A_in[25]), .A2 (A_in[24]));
NOR3_X1 i_148 (.ZN (n_92), .A1 (A_in[25]), .A2 (A_in[24]), .A3 (A_in[26]));
INV_X4 i_147 (.ZN (n_91), .A (A_in[3]));
INV_X4 i_146 (.ZN (n_88), .A (A_in[2]));
INV_X1 i_145 (.ZN (n_87), .A (A_in[1]));
INV_X4 i_144 (.ZN (n_74), .A (A_in[0]));
AOI21_X2 CLOCK_slo__sro_c2276 (.ZN (p_0[21]), .A (n_52), .B1 (CLOCK_slo__sro_n2263), .B2 (A_in[21]));
INV_X4 i_142 (.ZN (n_72), .A (n_73));
INV_X4 i_141 (.ZN (n_71), .A (A_in[7]));
INV_X1 i_140 (.ZN (n_131), .A (A_in[6]));
INV_X2 i_139 (.ZN (n_130), .A (A_in[5]));
INV_X4 i_138 (.ZN (n_129), .A (A_in[4]));
INV_X2 slo__c588 (.ZN (slo__n428), .A (A_in[6]));
INV_X4 i_136 (.ZN (n_127), .A (CLOCK_slo__sro_n1977));
INV_X1 i_135 (.ZN (n_126), .A (A_in[11]));
INV_X1 i_134 (.ZN (n_125), .A (opt_ipoPP_2));
INV_X1 i_133 (.ZN (n_124), .A (A_in[9]));
INV_X1 i_132 (.ZN (n_123), .A (A_in[8]));
NAND4_X4 i_131 (.ZN (n_122), .A1 (A_in[10]), .A2 (slo__n900), .A3 (slo__n760), .A4 (slo__n554));
INV_X4 i_130 (.ZN (n_121), .A (n_122));
INV_X1 i_129 (.ZN (n_120), .A (A_in[15]));
INV_X2 i_128 (.ZN (n_119), .A (A_in[14]));
INV_X1 i_127 (.ZN (n_118), .A (A_in[13]));
INV_X4 i_126 (.ZN (n_117), .A (A_in[12]));
NOR2_X1 sgo__sro_c247 (.ZN (n_116), .A1 (sgo__sro_n151), .A2 (sgo__sro_n150));
NAND2_X4 CLOCK_slo__sro_c2535 (.ZN (CLOCK_slo__sro_n2199), .A1 (n_102), .A2 (n_54));
NAND4_X4 i_123 (.ZN (n_114), .A1 (n_72), .A2 (n_127), .A3 (n_121), .A4 (slo__n960));
INV_X8 i_122 (.ZN (n_113), .A (n_114));
INV_X1 i_121 (.ZN (n_112), .A (A_in[23]));
INV_X4 i_120 (.ZN (n_111), .A (A_in[17]));
INV_X1 i_119 (.ZN (n_110), .A (A_in[16]));
INV_X4 slo__c822 (.ZN (slo__n648), .A (A_in[1]));
NAND3_X1 slo__c837 (.ZN (slo__n660), .A1 (n_72), .A2 (n_127), .A3 (n_121));
NAND2_X4 i_116 (.ZN (n_103), .A1 (n_105), .A2 (n_109));
INV_X4 i_115 (.ZN (n_102), .A (n_103));
INV_X4 CLOCK_slo__sro_c2536 (.ZN (CLOCK_slo__sro_n2198), .A (CLOCK_slo__sro_n2199));
INV_X4 i_113 (.ZN (n_89), .A (n_90));
NAND3_X1 i_112 (.ZN (n_86), .A1 (n_113), .A2 (n_89), .A3 (n_97));
NAND2_X1 i_111 (.ZN (n_85), .A1 (n_86), .A2 (A_in[30]));
INV_X1 i_110 (.ZN (n_84), .A (A_in[30]));
NAND4_X1 i_109 (.ZN (n_83), .A1 (n_113), .A2 (n_89), .A3 (n_84), .A4 (n_97));
NAND2_X1 i_108 (.ZN (n_82), .A1 (n_85), .A2 (n_83));
INV_X1 i_107 (.ZN (p_0[30]), .A (n_82));
NOR2_X1 i_106 (.ZN (n_81), .A1 (n_114), .A2 (n_90));
INV_X1 i_105 (.ZN (n_80), .A (A_in[28]));
AOI22_X1 i_103 (.ZN (p_0[29]), .A1 (CLOCK_slo__sro_n2595), .A2 (A_in[29]), .B1 (n_81), .B2 (n_97));
INV_X1 i_102 (.ZN (n_78), .A (CLOCK_slo__sro_n2595));
AOI21_X1 i_101 (.ZN (n_77), .A (n_80), .B1 (n_113), .B2 (n_89));
NOR2_X1 i_100 (.ZN (p_0[28]), .A1 (n_77), .A2 (n_78));
NAND3_X1 sgo__sro_c307 (.ZN (sgo__sro_n197), .A1 (n_118), .A2 (n_117), .A3 (n_119));
INV_X1 sgo__sro_c308 (.ZN (sgo__sro_n196), .A (sgo__sro_n197));
NAND3_X2 i_97 (.ZN (n_70), .A1 (n_113), .A2 (n_76), .A3 (n_92));
AOI21_X1 i_96 (.ZN (p_0[27]), .A (n_81), .B1 (n_70), .B2 (A_in[27]));
NAND4_X4 CLOCK_slo__sro_c2259 (.ZN (CLOCK_slo__sro_n1977), .A1 (n_130), .A2 (n_129)
    , .A3 (slo__n428), .A4 (n_71));
NAND3_X2 i_91 (.ZN (n_66), .A1 (n_113), .A2 (n_94), .A3 (n_76));
AOI22_X2 i_90 (.ZN (p_0[25]), .A1 (n_66), .A2 (A_in[25]), .B1 (n_93), .B2 (n_69));
INV_X1 i_89 (.ZN (n_65), .A (n_66));
AOI21_X1 i_88 (.ZN (n_64), .A (n_94), .B1 (n_113), .B2 (n_76));
NOR2_X1 i_87 (.ZN (p_0[24]), .A1 (n_64), .A2 (n_65));
NAND3_X2 i_86 (.ZN (n_63), .A1 (n_72), .A2 (n_127), .A3 (n_121));
INV_X1 CLOCK_sgo__sro_c1666 (.ZN (CLOCK_sgo__sro_n1461), .A (n_114));
NAND2_X1 i_84 (.ZN (n_61), .A1 (CLOCK_slo__n2408), .A2 (n_98));
NAND4_X4 CLOCK_slo__sro_c1979 (.ZN (n_73), .A1 (n_88), .A2 (slo__n648), .A3 (n_74), .A4 (n_91));
NAND2_X1 i_81 (.ZN (n_58), .A1 (n_59), .A2 (n_112));
INV_X1 i_80 (.ZN (n_57), .A (n_59));
NAND2_X1 i_79 (.ZN (n_56), .A1 (n_57), .A2 (A_in[23]));
NAND2_X1 i_78 (.ZN (p_0[23]), .A1 (n_56), .A2 (n_58));
NAND2_X1 i_77 (.ZN (n_55), .A1 (n_100), .A2 (n_99));
INV_X1 i_76 (.ZN (n_54), .A (n_55));
NAND2_X2 CLOCK_slo__mro_c2610 (.ZN (CLOCK_slo__mro_n2257), .A1 (CLOCK_slo__n2694), .A2 (CLOCK_slo__mro_n1619));
AOI21_X2 i_74 (.ZN (p_0[22]), .A (CLOCK_slo__n2461), .B1 (n_53), .B2 (A_in[22]));
INV_X1 i_73 (.ZN (n_52), .A (n_53));
INV_X2 CLOCK_slo__c2751 (.ZN (CLOCK_slo__n2408), .A (n_103));
OAI21_X1 i_70 (.ZN (n_50), .A (A_in[20]), .B1 (n_114), .B2 (n_103));
AND2_X2 i_69 (.ZN (p_0[20]), .A1 (n_50), .A2 (CLOCK_slo__sro_n2263));
NAND3_X1 i_68 (.ZN (n_49), .A1 (n_113), .A2 (n_106), .A3 (n_109));
NAND2_X1 i_67 (.ZN (n_48), .A1 (n_49), .A2 (n_107));
NAND4_X2 i_66 (.ZN (n_47), .A1 (n_113), .A2 (A_in[19]), .A3 (n_106), .A4 (n_109));
NAND2_X1 i_65 (.ZN (p_0[19]), .A1 (n_48), .A2 (n_47));
OAI21_X1 i_64 (.ZN (n_46), .A (A_in[18]), .B1 (n_114), .B2 (slo__xsl_n580));
AND2_X2 i_63 (.ZN (p_0[18]), .A1 (n_46), .A2 (n_49));
NAND2_X4 i_62 (.ZN (n_45), .A1 (n_113), .A2 (n_110));
INV_X2 i_61 (.ZN (n_44), .A (n_45));
NAND4_X1 CLOCK_slo__c2230 (.ZN (CLOCK_slo__n1960), .A1 (n_95), .A2 (n_94), .A3 (n_96), .A4 (n_104));
OAI21_X2 CLOCK_sgo__sro_c1669 (.ZN (p_0[17]), .A (CLOCK_sgo__sro_n1459), .B1 (n_44), .B2 (n_111));
AND2_X4 CLOCK_slo__sro_c2212 (.ZN (CLOCK_slo__sro_n1932), .A1 (n_98), .A2 (n_112));
NAND2_X4 CLOCK_slo__sro_c2619 (.ZN (CLOCK_slo__sro_n2265), .A1 (n_102), .A2 (n_99));
INV_X2 i_56 (.ZN (p_0[16]), .A (CLOCK_slo__mro_n2257));
NOR2_X4 slo__c1156 (.ZN (slo__n960), .A1 (sgo__sro_n150), .A2 (sgo__sro_n151));
NAND2_X1 i_54 (.ZN (n_39), .A1 (sgo__sro_n195), .A2 (n_120));
INV_X2 i_53 (.ZN (n_38), .A (sgo__sro_n195));
NAND2_X2 i_52 (.ZN (n_37), .A1 (n_38), .A2 (A_in[15]));
INV_X2 CLOCK_slo__c2232 (.ZN (n_101), .A (CLOCK_slo__n1960));
NAND2_X4 i_50 (.ZN (n_36), .A1 (opt_ipo_n1163), .A2 (n_117));
INV_X4 i_49 (.ZN (n_35), .A (n_36));
AOI21_X2 i_48 (.ZN (n_34), .A (n_119), .B1 (n_35), .B2 (n_118));
NOR2_X2 i_47 (.ZN (p_0[14]), .A1 (n_34), .A2 (n_38));
NAND2_X1 i_46 (.ZN (n_33), .A1 (n_35), .A2 (n_118));
NAND2_X2 i_45 (.ZN (n_32), .A1 (n_36), .A2 (A_in[13]));
NAND2_X1 i_44 (.ZN (n_31), .A1 (n_33), .A2 (n_32));
INV_X2 i_43 (.ZN (p_0[13]), .A (n_31));
NAND2_X1 i_42 (.ZN (n_30), .A1 (slo__n660), .A2 (A_in[12]));
NAND2_X1 i_41 (.ZN (n_29), .A1 (n_36), .A2 (n_30));
INV_X1 i_40 (.ZN (p_0[12]), .A (n_29));
NAND2_X2 i_39 (.ZN (n_28), .A1 (n_72), .A2 (CLOCK_slo__n1914));
INV_X2 i_38 (.ZN (n_27), .A (n_28));
NAND2_X2 slo__sro_c1272 (.ZN (p_0[15]), .A1 (n_37), .A2 (n_39));
INV_X2 i_36 (.ZN (n_25), .A (CLOCK_slo__sro_n1729));
NAND2_X2 i_35 (.ZN (n_24), .A1 (n_25), .A2 (n_125));
NAND2_X1 CLOCK_slo__sro_c2537 (.ZN (n_53), .A1 (CLOCK_slo__sro_n2198), .A2 (n_113));
NAND3_X1 i_33 (.ZN (n_22), .A1 (n_25), .A2 (A_in[11]), .A3 (n_125));
NAND2_X1 i_32 (.ZN (p_0[11]), .A1 (CLOCK_slo__sro_n2072), .A2 (n_22));
NAND2_X1 i_31 (.ZN (n_21), .A1 (n_26), .A2 (opt_ipoPP_2));
NAND2_X1 i_30 (.ZN (p_0[10]), .A1 (n_24), .A2 (n_21));
NAND2_X1 CLOCK_slo__sro_c2621 (.ZN (CLOCK_slo__sro_n2263), .A1 (CLOCK_slo__sro_n2264), .A2 (n_113));
OAI21_X1 i_28 (.ZN (n_19), .A (A_in[9]), .B1 (n_28), .B2 (A_in[8]));
NAND2_X1 i_27 (.ZN (n_18), .A1 (n_19), .A2 (n_26));
INV_X1 i_26 (.ZN (p_0[9]), .A (n_18));
XNOR2_X1 i_25 (.ZN (p_0[8]), .A (n_28), .B (n_123));
NOR2_X2 i_24 (.ZN (n_17), .A1 (n_73), .A2 (A_in[4]));
NAND2_X2 i_23 (.ZN (n_16), .A1 (n_17), .A2 (n_130));
INV_X2 i_22 (.ZN (n_15), .A (n_16));
NAND2_X2 i_21 (.ZN (n_14), .A1 (n_15), .A2 (n_131));
NAND2_X1 i_20 (.ZN (n_13), .A1 (n_14), .A2 (n_71));
NAND3_X1 i_19 (.ZN (n_12), .A1 (n_15), .A2 (A_in[7]), .A3 (n_131));
NAND2_X1 i_18 (.ZN (p_0[7]), .A1 (n_13), .A2 (n_12));
NAND2_X1 i_17 (.ZN (n_11), .A1 (n_16), .A2 (A_in[6]));
NAND2_X1 i_16 (.ZN (n_10), .A1 (n_14), .A2 (n_11));
INV_X1 i_15 (.ZN (p_0[6]), .A (n_10));
XNOR2_X1 i_14 (.ZN (n_9), .A (n_17), .B (n_130));
INV_X1 i_13 (.ZN (p_0[5]), .A (n_9));
XNOR2_X1 i_12 (.ZN (p_0[4]), .A (n_73), .B (A_in[4]));
INV_X4 CLOCK_slo__sro_c2620 (.ZN (CLOCK_slo__sro_n2264), .A (CLOCK_slo__sro_n2265));
NAND3_X1 i_10 (.ZN (n_7), .A1 (n_74), .A2 (n_88), .A3 (n_87));
NAND2_X1 i_9 (.ZN (n_6), .A1 (n_7), .A2 (A_in[3]));
NAND2_X1 i_8 (.ZN (n_5), .A1 (n_6), .A2 (n_73));
INV_X1 i_7 (.ZN (p_0[3]), .A (n_5));
NAND2_X1 i_6 (.ZN (n_4), .A1 (n_74), .A2 (n_87));
NAND2_X1 i_5 (.ZN (n_3), .A1 (n_4), .A2 (A_in[2]));
NAND2_X1 i_4 (.ZN (n_2), .A1 (n_3), .A2 (n_7));
INV_X1 i_3 (.ZN (p_0[2]), .A (n_2));
NAND2_X1 i_2 (.ZN (n_1), .A1 (A_in[0]), .A2 (A_in[1]));
NAND2_X1 i_1 (.ZN (n_0), .A1 (n_4), .A2 (n_1));
INV_X1 i_0 (.ZN (p_0[1]), .A (n_0));
INV_X2 slo__c784 (.ZN (slo__n602), .A (A_in[16]));
INV_X2 opt_ipo_c1426 (.ZN (opt_ipo_n1185), .A (n_61));
AND4_X2 sgo__c268 (.ZN (n_76), .A1 (n_98), .A2 (n_109), .A3 (n_105), .A4 (n_112));
NAND2_X2 sgo__sro_c245 (.ZN (sgo__sro_n151), .A1 (n_119), .A2 (slo__n967));
NAND2_X2 sgo__sro_c246 (.ZN (sgo__sro_n150), .A1 (slo__n1020), .A2 (n_117));
NAND2_X2 sgo__sro_c309 (.ZN (sgo__sro_n195), .A1 (opt_ipo_n1163), .A2 (sgo__sro_n196));
INV_X1 slo__xsl_c750 (.ZN (slo__xsl_n580), .A (n_109));
AOI22_X2 slo__sro_c1048 (.ZN (p_0[26]), .A1 (n_67), .A2 (A_in[26]), .B1 (n_69), .B2 (n_92));
NAND2_X2 CLOCK_slo__sro_c2027 (.ZN (CLOCK_slo__sro_n1729), .A1 (n_27), .A2 (CLOCK_slo__sro_n1730));
INV_X4 opt_ipo_c1412 (.ZN (opt_ipo_n1163), .A (n_63));
INV_X2 slo__c1109 (.ZN (slo__n900), .A (A_in[11]));
AND2_X4 slo__xsl_c753 (.ZN (n_109), .A1 (slo__n602), .A2 (n_111));
INV_X1 slo__c1227 (.ZN (slo__n1020), .A (A_in[13]));
INV_X2 slo__c717 (.ZN (slo__n554), .A (A_in[8]));
AND2_X1 CLOCK_slo__sro_c2026 (.ZN (CLOCK_slo__sro_n1730), .A1 (n_123), .A2 (n_124));
INV_X1 CLOCK_sgo__sro_c1667 (.ZN (CLOCK_sgo__sro_n1460), .A (slo__xsl_n580));
INV_X1 slo__c1166 (.ZN (slo__n967), .A (A_in[15]));
AND2_X1 slo__sro_c1259 (.ZN (slo__sro_n1043), .A1 (n_124), .A2 (n_123));
NAND2_X1 CLOCK_sgo__sro_c1668 (.ZN (CLOCK_sgo__sro_n1459), .A1 (CLOCK_sgo__sro_n1460), .A2 (CLOCK_sgo__sro_n1461));
NAND2_X1 slo__sro_c1260 (.ZN (n_26), .A1 (n_27), .A2 (slo__sro_n1043));
INV_X1 CLOCK_slo__c2188 (.ZN (CLOCK_slo__n1914), .A (CLOCK_slo__sro_n1977));
NAND2_X1 CLOCK_slo__mro_c1899 (.ZN (CLOCK_slo__mro_n1619), .A1 (n_114), .A2 (A_in[16]));
INV_X4 slo__c941 (.ZN (slo__n760), .A (A_in[9]));
NAND3_X4 CLOCK_slo__sro_c2213 (.ZN (n_90), .A1 (CLOCK_slo__sro_n1932), .A2 (n_101), .A3 (n_102));
NAND2_X2 CLOCK_slo__sro_c2374 (.ZN (CLOCK_slo__sro_n2072), .A1 (n_24), .A2 (n_126));
AND2_X2 CLOCK_slo__c3181 (.ZN (n_69), .A1 (n_113), .A2 (n_76));
INV_X2 CLOCK_slo__c2825 (.ZN (CLOCK_slo__n2461), .A (n_59));
NAND2_X2 CLOCK_slo__c3116 (.ZN (CLOCK_slo__n2694), .A1 (n_113), .A2 (n_110));
NAND3_X2 CLOCK_slo__sro_c2996 (.ZN (CLOCK_slo__sro_n2595), .A1 (n_113), .A2 (n_89), .A3 (n_80));
BUF_X2 CLOCK_slo__sro_c2884 (.Z (CLOCK_slo__sro_n2502), .A (n_116));
NAND3_X2 CLOCK_slo__sro_c2885 (.ZN (n_59), .A1 (opt_ipo_n1163), .A2 (opt_ipo_n1185), .A3 (CLOCK_slo__sro_n2502));

endmodule //datapath__0_129

module datapath__0_119 (opt_ipoPP_0, opt_ipoPP_3, Res_imm, p_0);

output [63:0] p_0;
input [63:0] Res_imm;
input opt_ipoPP_0;
input opt_ipoPP_3;
wire CLOCK_slo_n763;
wire CLOCK_slo__sro_n716;
wire CLOCK_slo__n859;
wire slo__sro_n463;
wire CLOCK_slo__sro_n764;
wire slo__xsl_n335;
wire n_14;
wire n_11;
wire n_13;
wire n_9;
wire n_10;
wire n_5;
wire n_8;
wire n_3;
wire n_4;
wire n_7;
wire n_2;
wire n_19;
wire n_22;
wire n_16;
wire n_18;
wire n_30;
wire n_24;
wire n_28;
wire n_29;
wire n_36;
wire n_12;
wire n_26;
wire n_41;
wire n_35;
wire n_50;
wire n_47;
wire n_62;
wire n_55;
wire n_70;
wire n_65;
wire n_79;
wire n_73;
wire n_94;
wire n_89;
wire n_104;
wire n_97;
wire n_103;
wire n_105;
wire n_212;
wire n_0;
wire n_203;
wire n_223;
wire n_1;
wire n_6;
wire n_15;
wire n_17;
wire n_20;
wire n_21;
wire n_23;
wire n_25;
wire n_27;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_39;
wire n_37;
wire n_38;
wire n_43;
wire n_40;
wire n_42;
wire n_45;
wire n_44;
wire n_46;
wire n_48;
wire n_49;
wire n_51;
wire n_53;
wire n_52;
wire n_54;
wire n_58;
wire n_56;
wire n_57;
wire n_59;
wire n_60;
wire n_61;
wire n_63;
wire n_64;
wire n_66;
wire sgo__sro_n189;
wire n_68;
wire n_69;
wire sgo__n70;
wire n_72;
wire n_76;
wire n_74;
wire sgo__sro_n188;
wire n_77;
wire n_78;
wire n_82;
wire n_80;
wire n_81;
wire slo__n432;
wire n_84;
wire slo__sro_n325;
wire sgo__sro_n238;
wire n_86;
wire n_87;
wire sgo__sro_n166;
wire n_90;
wire n_92;
wire n_93;
wire n_95;
wire n_96;
wire n_98;
wire sgo__n76;
wire n_99;
wire n_101;
wire n_102;
wire n_108;
wire n_106;
wire n_107;
wire n_110;
wire n_109;
wire n_115;
wire n_112;
wire n_111;
wire n_113;
wire slo__xsl_n363;
wire n_116;
wire sgo__sro_n187;
wire n_118;
wire n_119;
wire n_120;
wire n_122;
wire n_121;
wire n_124;
wire n_123;
wire n_125;
wire n_126;
wire n_127;
wire n_129;
wire n_128;
wire n_131;
wire n_130;
wire n_132;
wire n_133;
wire n_139;
wire n_138;
wire n_135;
wire n_137;
wire n_136;
wire n_141;
wire n_140;
wire n_145;
wire n_142;
wire n_144;
wire n_143;
wire n_146;
wire n_147;
wire n_149;
wire n_150;
wire n_152;
wire n_151;
wire n_153;
wire n_154;
wire n_155;
wire sgo__sro_n239;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_164;
wire n_163;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_175;
wire n_174;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_188;
wire n_186;
wire n_187;
wire n_189;
wire slo__xsl_n263;
wire n_191;
wire n_192;
wire n_193;
wire slo__n307;
wire n_195;
wire n_196;
wire n_197;
wire sgo__n11;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_204;
wire n_205;
wire n_206;
wire n_209;
wire n_207;
wire n_208;
wire n_210;
wire n_213;
wire n_211;
wire n_215;
wire n_214;
wire n_216;
wire n_220;
wire n_218;
wire n_217;
wire n_219;
wire n_222;
wire n_221;
wire n_224;
wire sgo__sro_n167;
wire sgo__sro_n168;
wire sgo__sro_n169;
wire sgo__sro_n170;
wire slo__n437;
wire CLOCK_slo__sro_n729;
wire CLOCK_slo__sro_n765;
wire CLOCK_slo__sro_n766;
wire CLOCK_slo__n781;
wire CLOCK_slo__n877;


INV_X1 i_287 (.ZN (n_224), .A (Res_imm[62]));
NAND3_X1 i_286 (.ZN (n_223), .A1 (n_216), .A2 (n_210), .A3 (n_224));
NAND2_X1 i_285 (.ZN (n_222), .A1 (n_199), .A2 (n_200));
NAND4_X1 i_284 (.ZN (n_221), .A1 (n_178), .A2 (n_157), .A3 (n_180), .A4 (slo__n432));
AND2_X1 slo__sro_c486 (.ZN (slo__sro_n325), .A1 (n_167), .A2 (Res_imm[53]));
NAND4_X2 i_282 (.ZN (n_219), .A1 (n_216), .A2 (CLOCK_slo__n859), .A3 (n_164), .A4 (n_163));
NOR4_X2 i_281 (.ZN (n_218), .A1 (n_208), .A2 (Res_imm[62]), .A3 (n_219), .A4 (Res_imm[63]));
AND3_X1 i_280 (.ZN (n_217), .A1 (n_84), .A2 (n_143), .A3 (n_181));
AOI22_X1 i_279 (.ZN (p_0[63]), .A1 (Res_imm[63]), .A2 (n_220), .B1 (n_218), .B2 (n_217));
INV_X1 i_278 (.ZN (n_216), .A (Res_imm[61]));
NAND4_X1 i_277 (.ZN (n_215), .A1 (n_216), .A2 (n_210), .A3 (n_199), .A4 (n_200));
NOR3_X2 i_275 (.ZN (n_213), .A1 (n_215), .A2 (n_214), .A3 (n_177));
INV_X1 i_274 (.ZN (n_212), .A (n_213));
NAND2_X1 i_273 (.ZN (n_211), .A1 (n_209), .A2 (n_207));
AOI21_X1 i_272 (.ZN (p_0[61]), .A (n_213), .B1 (Res_imm[61]), .B2 (n_211));
INV_X1 i_271 (.ZN (n_210), .A (Res_imm[60]));
AND4_X2 i_270 (.ZN (n_209), .A1 (n_73), .A2 (n_86), .A3 (n_143), .A4 (n_181));
NAND3_X2 i_269 (.ZN (n_208), .A1 (n_199), .A2 (n_200), .A3 (n_210));
NOR2_X2 i_268 (.ZN (n_207), .A1 (n_208), .A2 (n_177));
NAND3_X4 CLOCK_slo__sro_c840 (.ZN (n_201), .A1 (n_199), .A2 (n_180), .A3 (n_200));
AOI21_X1 i_266 (.ZN (p_0[59]), .A (n_203), .B1 (Res_imm[59]), .B2 (n_206));
NAND2_X1 i_265 (.ZN (n_206), .A1 (n_205), .A2 (n_157));
AND3_X1 i_264 (.ZN (n_205), .A1 (n_196), .A2 (n_178), .A3 (slo__n432));
INV_X1 i_263 (.ZN (n_204), .A (n_203));
NOR3_X4 i_262 (.ZN (n_203), .A1 (n_202), .A2 (n_177), .A3 (n_201));
NAND3_X4 i_261 (.ZN (n_202), .A1 (sgo__n70), .A2 (n_73), .A3 (n_80));
NOR2_X4 CLOCK_slo__c884 (.ZN (CLOCK_slo__n859), .A1 (n_176), .A2 (Res_imm[54]));
AND2_X1 i_259 (.ZN (n_200), .A1 (n_193), .A2 (n_189));
AND2_X1 sgo__sro_c301 (.ZN (sgo__sro_n189), .A1 (n_86), .A2 (n_74));
BUF_X4 sgo__c11 (.Z (n_147), .A (sgo__n11));
INV_X1 i_256 (.ZN (n_197), .A (Res_imm[58]));
AND4_X1 i_255 (.ZN (n_196), .A1 (n_197), .A2 (n_189), .A3 (n_193), .A4 (n_180));
NOR2_X2 slo__sro_c617 (.ZN (p_0[57]), .A1 (n_192), .A2 (slo__sro_n463));
CLKBUF_X1 CLOCK_slo___L1_c2_c786 (.Z (CLOCK_slo_n763), .A (Res_imm[28]));
NAND4_X1 i_252 (.ZN (n_195), .A1 (n_157), .A2 (n_188), .A3 (n_178), .A4 (slo__n432));
NOR3_X1 slo__c461 (.ZN (slo__n307), .A1 (n_221), .A2 (n_223), .A3 (n_222));
INV_X1 i_250 (.ZN (n_193), .A (Res_imm[57]));
NOR2_X1 slo__sro_c487 (.ZN (p_0[53]), .A1 (n_170), .A2 (slo__sro_n325));
NOR3_X4 i_248 (.ZN (n_191), .A1 (n_177), .A2 (Res_imm[56]), .A3 (Res_imm[57]));
INV_X1 slo__c463 (.ZN (n_220), .A (slo__n307));
INV_X1 i_246 (.ZN (n_189), .A (Res_imm[56]));
AND2_X1 i_245 (.ZN (n_188), .A1 (n_189), .A2 (n_180));
AND2_X1 i_244 (.ZN (n_187), .A1 (n_73), .A2 (n_86));
AND4_X1 i_243 (.ZN (n_186), .A1 (n_143), .A2 (n_187), .A3 (n_135), .A4 (slo__n437));
INV_X1 CLOCK_slo__sro_c789 (.ZN (CLOCK_slo__sro_n766), .A (Res_imm[27]));
AOI21_X1 i_241 (.ZN (p_0[55]), .A (n_183), .B1 (Res_imm[55]), .B2 (n_185));
NAND4_X1 i_240 (.ZN (n_185), .A1 (n_184), .A2 (n_157), .A3 (n_144), .A4 (slo__n432));
AND2_X1 i_239 (.ZN (n_184), .A1 (n_175), .A2 (CLOCK_slo__n877));
INV_X1 i_238 (.ZN (n_183), .A (n_182));
NAND4_X1 i_237 (.ZN (n_182), .A1 (n_181), .A2 (n_84), .A3 (slo__n437), .A4 (n_143));
AND2_X2 i_236 (.ZN (n_181), .A1 (n_180), .A2 (n_135));
AND3_X4 i_235 (.ZN (n_180), .A1 (n_179), .A2 (n_146), .A3 (n_145));
INV_X1 i_234 (.ZN (n_179), .A (Res_imm[55]));
INV_X1 i_233 (.ZN (n_178), .A (n_177));
AOI22_X2 CLOCK_slo__sro_c736 (.ZN (p_0[62]), .A1 (n_203), .A2 (n_0), .B1 (n_212), .B2 (Res_imm[62]));
NAND2_X4 i_231 (.ZN (n_176), .A1 (n_173), .A2 (n_169));
NOR2_X1 i_230 (.ZN (n_175), .A1 (n_176), .A2 (Res_imm[54]));
AND4_X1 i_229 (.ZN (n_174), .A1 (n_157), .A2 (n_162), .A3 (n_144), .A4 (slo__n432));
AOI22_X1 i_228 (.ZN (p_0[54]), .A1 (n_175), .A2 (n_174), .B1 (Res_imm[54]), .B2 (n_171));
INV_X1 i_227 (.ZN (n_173), .A (Res_imm[53]));
AND4_X4 i_226 (.ZN (n_172), .A1 (n_173), .A2 (n_144), .A3 (n_169), .A4 (n_157));
NAND3_X2 i_225 (.ZN (n_171), .A1 (n_172), .A2 (n_162), .A3 (slo__n432));
INV_X1 i_224 (.ZN (n_170), .A (n_171));
INV_X1 slo__xsl_c534 (.ZN (slo__xsl_n363), .A (n_73));
INV_X4 i_222 (.ZN (n_169), .A (Res_imm[52]));
AND2_X1 i_221 (.ZN (n_168), .A1 (n_169), .A2 (n_144));
NAND4_X1 i_220 (.ZN (n_167), .A1 (n_157), .A2 (n_168), .A3 (n_162), .A4 (slo__n432));
INV_X1 i_219 (.ZN (n_166), .A (n_167));
AOI21_X1 i_218 (.ZN (p_0[52]), .A (n_166), .B1 (Res_imm[52]), .B2 (n_161));
INV_X1 slo__xsl_c408 (.ZN (slo__xsl_n263), .A (n_192));
NOR2_X4 i_216 (.ZN (n_164), .A1 (Res_imm[51]), .A2 (Res_imm[50]));
AND2_X4 i_215 (.ZN (n_163), .A1 (n_153), .A2 (n_150));
AND2_X1 i_214 (.ZN (n_162), .A1 (n_164), .A2 (n_163));
NAND4_X1 i_213 (.ZN (n_161), .A1 (n_157), .A2 (n_144), .A3 (CLOCK_slo__n877), .A4 (n_135));
INV_X1 i_212 (.ZN (n_160), .A (n_161));
AOI21_X1 i_211 (.ZN (p_0[51]), .A (n_160), .B1 (Res_imm[51]), .B2 (sgo__sro_n166));
AOI21_X1 i_210 (.ZN (p_0[50]), .A (n_158), .B1 (n_159), .B2 (opt_ipoPP_0));
NAND4_X1 i_209 (.ZN (n_159), .A1 (n_157), .A2 (n_152), .A3 (n_144), .A4 (slo__n432));
INV_X2 i_208 (.ZN (n_158), .A (sgo__sro_n166));
OR2_X1 sgo__c129 (.ZN (sgo__n76), .A1 (Res_imm[59]), .A2 (Res_imm[58]));
AND2_X1 CLOCK_slo__sro_c758 (.ZN (CLOCK_slo__sro_n729), .A1 (n_182), .A2 (Res_imm[56]));
AND2_X1 i_205 (.ZN (n_155), .A1 (n_73), .A2 (n_86));
INV_X1 i_204 (.ZN (n_154), .A (opt_ipoPP_0));
INV_X2 i_203 (.ZN (n_153), .A (Res_imm[49]));
AND2_X1 i_202 (.ZN (n_152), .A1 (n_153), .A2 (n_150));
NAND3_X1 i_201 (.ZN (n_151), .A1 (n_73), .A2 (n_86), .A3 (n_147));
AOI22_X1 i_200 (.ZN (p_0[49]), .A1 (n_141), .A2 (n_152), .B1 (Res_imm[49]), .B2 (n_151));
INV_X1 i_199 (.ZN (n_150), .A (Res_imm[48]));
INV_X2 i_198 (.ZN (n_149), .A (n_144));
NAND3_X4 CLOCK_slo__sro_c776 (.ZN (n_177), .A1 (CLOCK_slo__n859), .A2 (n_163), .A3 (n_164));
NOR3_X2 i_196 (.ZN (sgo__n11), .A1 (CLOCK_slo__sro_n716), .A2 (opt_ipoPP_3), .A3 (n_149));
AOI22_X1 i_195 (.ZN (p_0[48]), .A1 (opt_ipoPP_3), .A2 (n_142), .B1 (n_84), .B2 (n_147));
INV_X2 i_194 (.ZN (n_146), .A (Res_imm[47]));
INV_X1 i_193 (.ZN (n_145), .A (Res_imm[46]));
NOR2_X4 i_192 (.ZN (n_144), .A1 (Res_imm[47]), .A2 (Res_imm[46]));
AND3_X4 i_191 (.ZN (n_143), .A1 (n_115), .A2 (n_128), .A3 (n_129));
NAND4_X1 i_190 (.ZN (n_142), .A1 (n_84), .A2 (n_135), .A3 (n_144), .A4 (n_143));
INV_X1 i_189 (.ZN (n_141), .A (n_142));
NAND2_X1 i_188 (.ZN (n_140), .A1 (n_145), .A2 (n_132));
AOI21_X2 i_187 (.ZN (p_0[47]), .A (n_141), .B1 (Res_imm[47]), .B2 (n_140));
XOR2_X1 i_186 (.Z (p_0[46]), .A (n_133), .B (Res_imm[46]));
AND2_X4 i_185 (.ZN (n_139), .A1 (n_128), .A2 (n_129));
AND2_X2 i_184 (.ZN (n_138), .A1 (n_116), .A2 (n_99));
AND2_X4 i_183 (.ZN (n_137), .A1 (n_107), .A2 (n_106));
NOR2_X2 i_182 (.ZN (n_136), .A1 (Res_imm[44]), .A2 (Res_imm[45]));
AND2_X4 i_181 (.ZN (n_135), .A1 (n_137), .A2 (n_136));
INV_X1 slo__xsl_c496 (.ZN (slo__xsl_n335), .A (n_115));
NAND3_X1 i_179 (.ZN (n_133), .A1 (n_73), .A2 (n_80), .A3 (sgo__n70));
INV_X1 i_178 (.ZN (n_132), .A (n_133));
AOI21_X1 i_177 (.ZN (p_0[45]), .A (n_132), .B1 (Res_imm[45]), .B2 (n_130));
INV_X1 i_176 (.ZN (n_131), .A (Res_imm[44]));
NAND2_X1 i_175 (.ZN (n_130), .A1 (n_131), .A2 (n_126));
AOI22_X1 i_174 (.ZN (p_0[44]), .A1 (n_131), .A2 (n_126), .B1 (Res_imm[44]), .B2 (n_127));
NOR2_X4 i_173 (.ZN (n_129), .A1 (Res_imm[43]), .A2 (Res_imm[42]));
NOR2_X4 i_172 (.ZN (n_128), .A1 (Res_imm[40]), .A2 (Res_imm[41]));
NAND3_X1 i_171 (.ZN (n_127), .A1 (n_129), .A2 (n_128), .A3 (n_110));
INV_X1 i_170 (.ZN (n_126), .A (n_127));
AOI21_X1 i_169 (.ZN (p_0[43]), .A (n_126), .B1 (Res_imm[43]), .B2 (n_123));
NAND3_X1 i_168 (.ZN (n_125), .A1 (n_84), .A2 (n_113), .A3 (n_120));
NOR3_X1 i_167 (.ZN (n_124), .A1 (n_125), .A2 (Res_imm[41]), .A3 (Res_imm[42]));
INV_X1 i_166 (.ZN (n_123), .A (n_124));
AOI21_X1 i_165 (.ZN (p_0[42]), .A (n_124), .B1 (n_121), .B2 (Res_imm[42]));
INV_X1 i_164 (.ZN (n_122), .A (Res_imm[41]));
NAND2_X1 i_163 (.ZN (n_121), .A1 (n_122), .A2 (n_118));
AOI22_X1 i_162 (.ZN (p_0[41]), .A1 (n_122), .A2 (n_118), .B1 (Res_imm[41]), .B2 (n_119));
NOR2_X1 i_161 (.ZN (n_120), .A1 (slo__xsl_n335), .A2 (Res_imm[40]));
NAND2_X1 i_160 (.ZN (n_119), .A1 (n_111), .A2 (n_120));
INV_X1 i_159 (.ZN (n_118), .A (n_119));
AOI21_X1 i_158 (.ZN (p_0[40]), .A (n_118), .B1 (Res_imm[40]), .B2 (n_109));
INV_X4 sgo__c47 (.ZN (n_157), .A (sgo__sro_n187));
NOR3_X4 i_156 (.ZN (n_116), .A1 (Res_imm[32]), .A2 (Res_imm[38]), .A3 (Res_imm[39]));
AND4_X4 slo__xsl_c537 (.ZN (n_73), .A1 (n_74), .A2 (n_66), .A3 (n_56), .A4 (n_43));
INV_X1 slo__c602 (.ZN (slo__n437), .A (n_177));
AND2_X1 i_153 (.ZN (n_113), .A1 (n_107), .A2 (n_106));
NAND2_X4 i_152 (.ZN (n_112), .A1 (n_84), .A2 (n_113));
INV_X1 i_151 (.ZN (n_111), .A (n_112));
NOR2_X2 i_150 (.ZN (n_110), .A1 (slo__xsl_n335), .A2 (n_112));
INV_X1 i_149 (.ZN (n_109), .A (n_110));
AOI21_X1 i_148 (.ZN (p_0[39]), .A (n_110), .B1 (Res_imm[39]), .B2 (n_102));
INV_X1 i_147 (.ZN (n_108), .A (Res_imm[38]));
INV_X1 i_146 (.ZN (n_107), .A (Res_imm[37]));
INV_X4 i_145 (.ZN (n_106), .A (Res_imm[36]));
NAND3_X1 i_144 (.ZN (n_105), .A1 (n_84), .A2 (n_98), .A3 (n_106));
INV_X1 i_143 (.ZN (n_104), .A (n_105));
NOR2_X2 i_142 (.ZN (n_103), .A1 (Res_imm[37]), .A2 (n_105));
NAND2_X2 i_141 (.ZN (n_102), .A1 (n_108), .A2 (n_103));
OAI21_X2 i_140 (.ZN (n_101), .A (n_102), .B1 (n_108), .B2 (n_103));
INV_X1 i_139 (.ZN (p_0[38]), .A (n_101));
AND4_X2 slo__xsl_c411 (.ZN (n_192), .A1 (n_191), .A2 (n_181), .A3 (n_143), .A4 (n_84));
NOR3_X4 i_137 (.ZN (n_99), .A1 (Res_imm[35]), .A2 (Res_imm[33]), .A3 (Res_imm[34]));
AND2_X1 i_136 (.ZN (n_98), .A1 (n_90), .A2 (n_99));
NAND2_X1 i_135 (.ZN (n_97), .A1 (n_84), .A2 (n_98));
AOI22_X1 i_134 (.ZN (p_0[35]), .A1 (n_84), .A2 (n_98), .B1 (Res_imm[35]), .B2 (n_96));
INV_X1 i_133 (.ZN (n_96), .A (n_95));
AOI21_X1 i_132 (.ZN (p_0[34]), .A (n_95), .B1 (Res_imm[34]), .B2 (n_93));
NOR2_X1 i_131 (.ZN (n_95), .A1 (n_93), .A2 (Res_imm[34]));
INV_X1 i_130 (.ZN (n_94), .A (n_93));
NAND4_X1 i_129 (.ZN (n_93), .A1 (n_92), .A2 (n_73), .A3 (n_90), .A4 (n_86));
INV_X1 i_128 (.ZN (n_92), .A (Res_imm[33]));
AOI22_X2 CLOCK_slo__sro_c833 (.ZN (p_0[60]), .A1 (n_207), .A2 (n_209), .B1 (n_204), .B2 (Res_imm[60]));
INV_X1 i_126 (.ZN (n_90), .A (Res_imm[32]));
NAND2_X1 i_125 (.ZN (n_89), .A1 (n_84), .A2 (n_90));
AOI22_X1 i_124 (.ZN (p_0[32]), .A1 (n_84), .A2 (n_90), .B1 (sgo__sro_n238), .B2 (Res_imm[32]));
NAND4_X2 sgo__c113 (.ZN (CLOCK_slo__n781), .A1 (n_135), .A2 (n_138), .A3 (n_139), .A4 (n_87));
INV_X4 i_122 (.ZN (n_87), .A (Res_imm[31]));
AND3_X4 i_121 (.ZN (n_86), .A1 (n_82), .A2 (n_81), .A3 (n_87));
AND2_X4 slo__xsl_c499 (.ZN (n_115), .A1 (n_116), .A2 (n_99));
INV_X8 i_119 (.ZN (n_84), .A (sgo__sro_n238));
AOI21_X1 i_118 (.ZN (p_0[31]), .A (n_84), .B1 (Res_imm[31]), .B2 (n_78));
CLKBUF_X3 slo__c597 (.Z (slo__n432), .A (n_135));
INV_X1 i_116 (.ZN (n_82), .A (Res_imm[30]));
INV_X1 i_115 (.ZN (n_81), .A (Res_imm[29]));
NOR2_X1 i_114 (.ZN (n_80), .A1 (Res_imm[30]), .A2 (Res_imm[29]));
NOR2_X1 i_113 (.ZN (n_79), .A1 (slo__xsl_n363), .A2 (Res_imm[29]));
NAND2_X1 i_112 (.ZN (n_78), .A1 (n_82), .A2 (n_79));
OAI21_X1 i_111 (.ZN (n_77), .A (n_78), .B1 (n_82), .B2 (n_79));
INV_X1 i_110 (.ZN (p_0[30]), .A (n_77));
INV_X1 i_109 (.ZN (n_76), .A (CLOCK_slo_n763));
AND2_X2 sgo__sro_c302 (.ZN (sgo__sro_n188), .A1 (sgo__sro_n189), .A2 (n_64));
INV_X2 CLOCK_slo__c817 (.ZN (sgo__n70), .A (CLOCK_slo__n781));
AND2_X1 slo__sro_c616 (.ZN (slo__sro_n463), .A1 (n_195), .A2 (Res_imm[57]));
OAI21_X1 i_105 (.ZN (n_72), .A (slo__xsl_n363), .B1 (n_76), .B2 (n_68));
INV_X1 i_104 (.ZN (p_0[28]), .A (n_72));
INV_X4 sgo__c131 (.ZN (n_199), .A (sgo__n76));
NOR2_X1 i_102 (.ZN (n_70), .A1 (n_65), .A2 (Res_imm[26]));
INV_X1 i_101 (.ZN (n_69), .A (n_70));
NOR2_X1 i_100 (.ZN (n_68), .A1 (Res_imm[27]), .A2 (n_69));
AOI21_X1 i_99 (.ZN (p_0[27]), .A (n_68), .B1 (Res_imm[27]), .B2 (n_69));
NAND2_X4 sgo__sro_c303 (.ZN (sgo__sro_n187), .A1 (n_143), .A2 (sgo__sro_n188));
NOR3_X2 i_97 (.ZN (n_66), .A1 (Res_imm[25]), .A2 (Res_imm[24]), .A3 (Res_imm[23]));
NAND4_X1 i_96 (.ZN (n_65), .A1 (n_56), .A2 (n_58), .A3 (n_57), .A4 (n_66));
INV_X1 i_95 (.ZN (n_64), .A (n_65));
AOI21_X1 i_94 (.ZN (p_0[25]), .A (n_64), .B1 (Res_imm[25]), .B2 (n_61));
INV_X1 i_93 (.ZN (n_63), .A (Res_imm[24]));
NOR2_X1 i_92 (.ZN (n_62), .A1 (n_55), .A2 (Res_imm[23]));
NAND2_X1 i_91 (.ZN (n_61), .A1 (n_63), .A2 (n_62));
OAI21_X1 i_90 (.ZN (n_60), .A (n_61), .B1 (n_63), .B2 (n_62));
INV_X1 i_89 (.ZN (p_0[24]), .A (n_60));
INV_X1 i_88 (.ZN (n_59), .A (Res_imm[22]));
INV_X1 i_87 (.ZN (n_58), .A (n_44));
INV_X1 i_86 (.ZN (n_57), .A (n_45));
AND4_X1 i_85 (.ZN (n_56), .A1 (n_59), .A2 (n_53), .A3 (n_52), .A4 (n_48));
NAND3_X1 i_84 (.ZN (n_55), .A1 (n_58), .A2 (n_56), .A3 (n_57));
INV_X1 i_83 (.ZN (n_54), .A (n_55));
AOI21_X1 i_82 (.ZN (p_0[22]), .A (n_54), .B1 (Res_imm[22]), .B2 (n_51));
INV_X1 i_81 (.ZN (n_53), .A (Res_imm[21]));
INV_X2 i_80 (.ZN (n_52), .A (Res_imm[20]));
NAND4_X1 i_79 (.ZN (n_51), .A1 (n_53), .A2 (n_48), .A3 (n_52), .A4 (n_43));
NOR2_X1 i_78 (.ZN (n_50), .A1 (Res_imm[20]), .A2 (n_47));
OAI21_X1 i_77 (.ZN (n_49), .A (n_51), .B1 (n_53), .B2 (n_50));
INV_X1 i_76 (.ZN (p_0[21]), .A (n_49));
INV_X1 i_75 (.ZN (n_48), .A (Res_imm[19]));
NAND2_X1 i_74 (.ZN (n_47), .A1 (n_48), .A2 (n_43));
AOI22_X1 i_73 (.ZN (p_0[19]), .A1 (n_48), .A2 (n_43), .B1 (Res_imm[19]), .B2 (n_42));
NOR2_X1 i_72 (.ZN (n_46), .A1 (n_24), .A2 (n_37));
NAND2_X1 i_71 (.ZN (n_45), .A1 (n_39), .A2 (n_46));
OR2_X1 i_70 (.ZN (n_44), .A1 (Res_imm[18]), .A2 (Res_imm[17]));
NOR2_X1 i_69 (.ZN (n_43), .A1 (n_45), .A2 (n_44));
INV_X1 i_68 (.ZN (n_42), .A (n_43));
NOR2_X1 i_67 (.ZN (n_41), .A1 (Res_imm[17]), .A2 (n_35));
INV_X1 i_66 (.ZN (n_40), .A (n_41));
AOI21_X1 i_65 (.ZN (p_0[18]), .A (n_43), .B1 (Res_imm[18]), .B2 (n_40));
INV_X1 i_64 (.ZN (n_39), .A (Res_imm[16]));
INV_X1 i_63 (.ZN (n_38), .A (Res_imm[15]));
NAND4_X1 i_62 (.ZN (n_37), .A1 (n_38), .A2 (n_33), .A3 (n_32), .A4 (n_31));
NOR2_X1 i_61 (.ZN (n_36), .A1 (n_24), .A2 (n_37));
NAND2_X1 i_60 (.ZN (n_35), .A1 (n_39), .A2 (n_36));
OAI21_X1 i_59 (.ZN (n_34), .A (n_35), .B1 (n_39), .B2 (n_36));
INV_X1 i_58 (.ZN (p_0[16]), .A (n_34));
INV_X1 i_57 (.ZN (n_33), .A (Res_imm[14]));
INV_X1 i_56 (.ZN (n_32), .A (Res_imm[13]));
INV_X1 i_55 (.ZN (n_31), .A (Res_imm[12]));
NOR2_X1 i_54 (.ZN (n_30), .A1 (Res_imm[12]), .A2 (n_24));
INV_X1 i_53 (.ZN (n_29), .A (n_30));
NOR2_X1 i_52 (.ZN (n_28), .A1 (Res_imm[13]), .A2 (n_29));
INV_X1 i_51 (.ZN (n_27), .A (n_28));
NOR2_X1 i_50 (.ZN (n_26), .A1 (Res_imm[14]), .A2 (n_27));
AOI21_X1 i_49 (.ZN (p_0[14]), .A (n_26), .B1 (Res_imm[14]), .B2 (n_27));
INV_X1 i_48 (.ZN (n_25), .A (Res_imm[11]));
NAND4_X1 i_47 (.ZN (n_24), .A1 (n_1), .A2 (n_21), .A3 (n_20), .A4 (n_25));
OAI21_X1 i_45 (.ZN (n_23), .A (n_24), .B1 (n_25), .B2 (n_15));
INV_X1 i_44 (.ZN (p_0[11]), .A (n_23));
INV_X1 i_42 (.ZN (n_22), .A (n_1));
INV_X1 i_41 (.ZN (n_21), .A (Res_imm[10]));
NOR2_X1 i_40 (.ZN (n_20), .A1 (Res_imm[9]), .A2 (Res_imm[8]));
NOR2_X1 i_39 (.ZN (n_19), .A1 (n_22), .A2 (Res_imm[8]));
INV_X1 i_38 (.ZN (n_18), .A (n_19));
NAND2_X1 i_36 (.ZN (n_17), .A1 (n_1), .A2 (n_20));
INV_X1 i_35 (.ZN (n_16), .A (n_17));
NOR2_X1 i_33 (.ZN (n_15), .A1 (Res_imm[10]), .A2 (n_17));
AOI21_X1 i_32 (.ZN (p_0[10]), .A (n_15), .B1 (Res_imm[10]), .B2 (n_17));
NOR2_X1 i_31 (.ZN (n_14), .A1 (Res_imm[1]), .A2 (Res_imm[0]));
INV_X1 i_30 (.ZN (n_13), .A (n_14));
NOR2_X1 i_29 (.ZN (n_11), .A1 (Res_imm[2]), .A2 (n_13));
INV_X1 i_28 (.ZN (n_10), .A (n_11));
NOR2_X1 i_27 (.ZN (n_9), .A1 (Res_imm[3]), .A2 (n_10));
INV_X1 i_26 (.ZN (n_8), .A (n_9));
NOR4_X1 i_25 (.ZN (n_7), .A1 (Res_imm[6]), .A2 (Res_imm[5]), .A3 (Res_imm[4]), .A4 (n_8));
INV_X1 i_22 (.ZN (n_6), .A (n_7));
NOR2_X1 i_21 (.ZN (n_1), .A1 (Res_imm[7]), .A2 (n_6));
AOI21_X1 i_20 (.ZN (p_0[7]), .A (n_1), .B1 (Res_imm[7]), .B2 (n_6));
INV_X1 i_19 (.ZN (n_0), .A (n_223));
NAND4_X2 CLOCK_slo__sro_c747 (.ZN (CLOCK_slo__sro_n716), .A1 (n_139), .A2 (n_138)
    , .A3 (n_136), .A4 (n_137));
AOI21_X1 i_17 (.ZN (p_0[37]), .A (n_103), .B1 (Res_imm[37]), .B2 (n_105));
AOI21_X1 i_16 (.ZN (p_0[36]), .A (n_104), .B1 (Res_imm[36]), .B2 (n_97));
AOI21_X1 i_15 (.ZN (p_0[33]), .A (n_94), .B1 (Res_imm[33]), .B2 (n_89));
AOI21_X1 i_46 (.ZN (p_0[29]), .A (n_79), .B1 (Res_imm[29]), .B2 (slo__xsl_n363));
AOI21_X1 i_43 (.ZN (p_0[26]), .A (n_70), .B1 (Res_imm[26]), .B2 (n_65));
AOI21_X1 i_14 (.ZN (p_0[23]), .A (n_62), .B1 (Res_imm[23]), .B2 (n_55));
AOI21_X1 i_37 (.ZN (p_0[20]), .A (n_50), .B1 (Res_imm[20]), .B2 (n_47));
AOI21_X1 i_34 (.ZN (p_0[17]), .A (n_41), .B1 (Res_imm[17]), .B2 (n_35));
INV_X1 i_13 (.ZN (n_12), .A (n_26));
AOI21_X1 i_12 (.ZN (p_0[15]), .A (n_36), .B1 (Res_imm[15]), .B2 (n_12));
AOI21_X1 i_24 (.ZN (p_0[13]), .A (n_28), .B1 (Res_imm[13]), .B2 (n_29));
AOI21_X1 i_23 (.ZN (p_0[12]), .A (n_30), .B1 (Res_imm[12]), .B2 (n_24));
AOI21_X1 i_11 (.ZN (p_0[9]), .A (n_16), .B1 (Res_imm[9]), .B2 (n_18));
AOI21_X1 i_10 (.ZN (p_0[8]), .A (n_19), .B1 (Res_imm[8]), .B2 (n_22));
NOR2_X1 i_9 (.ZN (n_5), .A1 (Res_imm[4]), .A2 (n_8));
INV_X1 i_8 (.ZN (n_4), .A (n_5));
NOR2_X1 i_7 (.ZN (n_3), .A1 (Res_imm[5]), .A2 (n_4));
INV_X1 i_6 (.ZN (n_2), .A (n_3));
AOI21_X1 i_5 (.ZN (p_0[6]), .A (n_7), .B1 (Res_imm[6]), .B2 (n_2));
AOI21_X1 i_4 (.ZN (p_0[5]), .A (n_3), .B1 (Res_imm[5]), .B2 (n_4));
AOI21_X1 i_3 (.ZN (p_0[4]), .A (n_5), .B1 (Res_imm[4]), .B2 (n_8));
AOI21_X1 i_2 (.ZN (p_0[3]), .A (n_9), .B1 (Res_imm[3]), .B2 (n_10));
AOI21_X1 i_1 (.ZN (p_0[2]), .A (n_11), .B1 (Res_imm[2]), .B2 (n_13));
AOI21_X1 i_0 (.ZN (p_0[1]), .A (n_14), .B1 (Res_imm[1]), .B2 (Res_imm[0]));
AND2_X1 sgo__sro_c370 (.ZN (sgo__sro_n239), .A1 (n_54), .A2 (n_66));
NAND3_X4 sgo__sro_c371 (.ZN (sgo__sro_n238), .A1 (n_86), .A2 (sgo__sro_n239), .A3 (n_74));
AOI22_X1 slo__sro_c607 (.ZN (p_0[58]), .A1 (n_186), .A2 (n_196), .B1 (slo__xsl_n263), .B2 (Res_imm[58]));
NAND2_X1 sgo__sro_c277 (.ZN (sgo__sro_n170), .A1 (n_153), .A2 (n_154));
INV_X1 sgo__sro_c278 (.ZN (sgo__sro_n169), .A (sgo__sro_n170));
NAND2_X1 sgo__sro_c279 (.ZN (sgo__sro_n168), .A1 (n_155), .A2 (sgo__sro_n169));
INV_X2 sgo__sro_c280 (.ZN (sgo__sro_n167), .A (sgo__sro_n168));
NAND2_X4 sgo__sro_c281 (.ZN (sgo__sro_n166), .A1 (n_147), .A2 (sgo__sro_n167));
AOI21_X1 CLOCK_slo__sro_c759 (.ZN (p_0[56]), .A (CLOCK_slo__sro_n729), .B1 (n_186), .B2 (n_188));
INV_X1 CLOCK_slo__sro_c790 (.ZN (CLOCK_slo__sro_n765), .A (Res_imm[26]));
NAND2_X1 CLOCK_slo__sro_c791 (.ZN (CLOCK_slo__sro_n764), .A1 (CLOCK_slo__sro_n765), .A2 (CLOCK_slo__sro_n766));
NOR2_X4 CLOCK_slo__sro_c792 (.ZN (n_74), .A1 (Res_imm[28]), .A2 (CLOCK_slo__sro_n764));
AND2_X1 CLOCK_slo__c902 (.ZN (CLOCK_slo__n877), .A1 (n_164), .A2 (n_163));
NAND3_X1 CLOCK_slo__sro_c807 (.ZN (n_214), .A1 (n_181), .A2 (n_143), .A3 (n_84));

endmodule //datapath__0_119

module datapath (carry_in, Res_in, Res_out);

output [63:0] Res_out;
input [63:0] Res_in;
input [63:0] carry_in;
wire slo__xsl_n495;
wire CLOCK_slo__sro_n1317;
wire CLOCK_slo__xsl_n1578;
wire CLOCK_slo__sro_n1363;
wire slo__n476;
wire CLOCK_slo__n1548;
wire n_1;
wire n_22;
wire n_20;
wire n_17;
wire n_2;
wire n_5;
wire n_25;
wire n_19;
wire n_3;
wire n_4;
wire n_24;
wire n_16;
wire n_6;
wire n_21;
wire n_23;
wire n_31;
wire n_8;
wire CLOCK_slo__sro_n1388;
wire n_30;
wire n_18;
wire n_10;
wire n_11;
wire n_28;
wire n_29;
wire n_27;
wire n_50;
wire n_49;
wire n_34;
wire n_41;
wire n_35;
wire n_104;
wire n_92;
wire n_36;
wire n_39;
wire n_95;
wire n_0;
wire n_42;
wire n_37;
wire n_38;
wire n_40;
wire n_91;
wire n_78;
wire n_88;
wire n_93;
wire n_43;
wire n_44;
wire n_115;
wire n_119;
wire n_122;
wire n_45;
wire n_124;
wire n_46;
wire n_152;
wire n_86;
wire n_254;
wire n_76;
wire CLOCK_slo__xsl_n1508;
wire n_255;
wire n_96;
wire n_97;
wire n_110;
wire n_373;
wire n_390;
wire n_98;
wire n_102;
wire slo__n536;
wire n_391;
wire n_101;
wire n_99;
wire n_379;
wire n_106;
wire n_100;
wire n_268;
wire n_111;
wire n_267;
wire n_103;
wire n_272;
wire n_270;
wire n_107;
wire n_274;
wire n_108;
wire n_109;
wire n_237;
wire n_399;
wire n_114;
wire n_275;
wire n_378;
wire n_384;
wire n_116;
wire sgo__n190;
wire n_120;
wire n_284;
wire n_278;
wire n_118;
wire n_131;
wire n_177;
wire n_279;
wire n_121;
wire n_125;
wire n_178;
wire n_276;
wire n_128;
wire n_126;
wire n_132;
wire n_127;
wire n_130;
wire n_331;
wire CLOCK_slo__n1598;
wire n_280;
wire n_281;
wire n_285;
wire n_282;
wire n_140;
wire CLOCK_slo__sro_n1387;
wire n_144;
wire n_319;
wire n_167;
wire n_142;
wire n_295;
wire n_180;
wire n_166;
wire n_145;
wire n_318;
wire n_181;
wire n_183;
wire n_147;
wire n_146;
wire n_151;
wire n_294;
wire n_289;
wire n_150;
wire n_288;
wire n_298;
wire n_172;
wire n_324;
wire n_320;
wire n_154;
wire n_290;
wire n_163;
wire n_332;
wire n_165;
wire n_296;
wire n_313;
wire n_312;
wire n_173;
wire n_184;
wire sgo__sro_n74;
wire n_193;
wire n_190;
wire n_302;
wire n_195;
wire n_341;
wire n_345;
wire n_207;
wire n_208;
wire sgo__sro_n75;
wire n_212;
wire n_335;
wire n_210;
wire n_342;
wire n_211;
wire n_334;
wire n_213;
wire n_344;
wire n_233;
wire n_238;
wire n_219;
wire n_216;
wire n_221;
wire n_218;
wire n_217;
wire n_355;
wire n_339;
wire n_227;
wire n_220;
wire n_340;
wire n_224;
wire n_222;
wire n_228;
wire n_223;
wire n_226;
wire n_356;
wire n_388;
wire n_225;
wire n_354;
wire n_346;
wire n_337;
wire n_338;
wire n_410;
wire n_400;
wire n_416;
wire n_263;
wire n_432;
wire n_436;
wire n_434;
wire n_433;
wire n_7;
wire n_252;
wire n_371;
wire n_283;
wire n_386;
wire n_277;
wire n_202;
wire n_196;
wire n_194;
wire n_293;
wire sgo__sro_n144;
wire n_198;
wire n_292;
wire n_352;
wire n_326;
wire n_203;
wire n_206;
wire n_300;
wire n_205;
wire n_236;
wire sgo__sro_n48;
wire n_240;
wire n_303;
wire n_242;
wire n_305;
wire n_304;
wire n_257;
wire n_311;
wire slo__sro_n375;
wire n_261;
wire n_308;
wire n_307;
wire slo__n516;
wire n_358;
wire n_301;
wire n_262;
wire n_306;
wire n_269;
wire n_309;
wire n_271;
wire n_314;
wire n_350;
wire n_357;
wire n_362;
wire n_347;
wire n_374;
wire n_418;
wire n_385;
wire n_395;
wire n_409;
wire n_408;
wire n_13;
wire n_12;
wire n_14;
wire n_15;
wire n_26;
wire n_33;
wire n_32;
wire n_48;
wire n_51;
wire sgo__sro_n26;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_62;
wire n_59;
wire n_61;
wire n_60;
wire n_65;
wire n_64;
wire n_63;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_72;
wire n_71;
wire n_75;
wire n_74;
wire n_73;
wire n_77;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire sgo__sro_n145;
wire n_84;
wire n_85;
wire n_87;
wire n_89;
wire n_90;
wire n_94;
wire n_105;
wire n_112;
wire n_113;
wire n_123;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_139;
wire n_138;
wire n_148;
wire n_143;
wire n_149;
wire n_153;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire CLOCK_sgo__n1177;
wire n_168;
wire n_169;
wire n_171;
wire n_170;
wire n_175;
wire n_174;
wire n_179;
wire n_188;
wire n_182;
wire CLOCK_slo__n1604;
wire n_185;
wire n_187;
wire n_189;
wire n_191;
wire CLOCK_slo__n1537;
wire n_199;
wire n_200;
wire sgo__sro_n49;
wire n_204;
wire n_214;
wire n_215;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_235;
wire n_239;
wire n_241;
wire n_243;
wire n_244;
wire n_248;
wire n_245;
wire n_247;
wire n_246;
wire n_249;
wire n_250;
wire n_251;
wire n_253;
wire n_259;
wire sgo__sro_n25;
wire slo__mro_n397;
wire n_265;
wire n_287;
wire n_286;
wire n_291;
wire n_299;
wire n_297;
wire n_310;
wire n_316;
wire n_322;
wire n_315;
wire n_325;
wire n_323;
wire n_317;
wire n_321;
wire n_329;
wire n_327;
wire n_333;
wire n_330;
wire n_328;
wire n_336;
wire n_343;
wire n_351;
wire n_349;
wire n_359;
wire n_360;
wire n_361;
wire n_363;
wire n_364;
wire n_365;
wire n_367;
wire n_368;
wire sgo__sro_n76;
wire n_370;
wire n_372;
wire n_375;
wire n_376;
wire sgo__sro_n108;
wire sgo__sro_n11;
wire n_381;
wire n_382;
wire n_383;
wire slo__sro_n469;
wire n_389;
wire n_392;
wire n_393;
wire n_394;
wire n_396;
wire n_397;
wire n_398;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_406;
wire n_407;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_417;
wire n_421;
wire n_419;
wire n_420;
wire n_423;
wire n_422;
wire n_426;
wire n_429;
wire n_425;
wire n_424;
wire n_427;
wire n_428;
wire n_431;
wire n_430;
wire n_435;
wire slo__xsl_n594;
wire sgo__sro_n109;
wire sgo__sro_n110;
wire sgo__sro_n146;
wire sgo__sro_n210;
wire sgo__sro_n211;
wire sgo__sro_n174;
wire CLOCK_slo__sro_n1333;
wire sgo__sro_n176;
wire sgo__sro_n177;
wire sgo__sro_n178;
wire CLOCK_slo__mro_n1456;
wire sgo__sro_n301;
wire sgo__sro_n302;
wire sgo__sro_n303;
wire sgo__n290;
wire slo__mro_n380;
wire slo__mro_n414;
wire slo__mro_n415;
wire slo__mro_n416;
wire slo__n543;
wire slo__n626;
wire slo__xsl_n558;
wire opt_ipo_n883;
wire CLOCK_slo__sro_n1310;
wire CLOCK_opt_ipo_n1035;
wire CLOCK_slo__sro_n1364;
wire opt_ipo_n987;
wire CLOCK_slo__sro_n1389;
wire CLOCK_slo__mro_n1454;
wire CLOCK_slo__mro_n1455;
wire opt_ipo_n1006;
wire opt_ipo_n1007;
wire CLOCK_slo__mro_n1453;
wire opt_ipo_n737;
wire CLOCK_opt_ipo_n1068;
wire CLOCK_slo__mro_n1442;


INV_X1 i_491 (.ZN (n_436), .A (carry_in[62]));
INV_X1 i_490 (.ZN (n_435), .A (n_424));
AOI21_X2 slo__mro_c666 (.ZN (slo__mro_n380), .A (n_259), .B1 (n_254), .B2 (opt_ipo_n737));
AOI21_X1 i_488 (.ZN (n_433), .A (n_435), .B1 (n_425), .B2 (n_426));
AND3_X4 i_487 (.ZN (n_432), .A1 (n_434), .A2 (n_433), .A3 (n_436));
NAND2_X1 i_486 (.ZN (n_431), .A1 (n_400), .A2 (n_415));
NAND2_X1 i_485 (.ZN (n_430), .A1 (n_396), .A2 (n_420));
NOR2_X1 i_484 (.ZN (n_429), .A1 (n_431), .A2 (n_430));
AOI21_X1 i_483 (.ZN (n_428), .A (n_431), .B1 (n_397), .B2 (n_401));
AOI21_X1 i_482 (.ZN (n_427), .A (n_428), .B1 (carry_in[59]), .B2 (Res_in[59]));
OAI21_X1 i_481 (.ZN (n_426), .A (n_419), .B1 (n_421), .B2 (n_427));
OR2_X1 i_480 (.ZN (n_425), .A1 (carry_in[61]), .A2 (Res_in[61]));
NAND2_X1 i_479 (.ZN (n_424), .A1 (carry_in[61]), .A2 (Res_in[61]));
NAND2_X1 i_478 (.ZN (n_423), .A1 (n_425), .A2 (n_424));
AOI21_X2 i_477 (.ZN (n_422), .A (n_426), .B1 (n_395), .B2 (n_429));
XOR2_X2 i_476 (.Z (Res_out[61]), .A (n_422), .B (n_423));
NOR2_X1 i_475 (.ZN (n_421), .A1 (carry_in[60]), .A2 (Res_in[60]));
INV_X1 i_474 (.ZN (n_420), .A (n_421));
NAND2_X1 i_473 (.ZN (n_419), .A1 (carry_in[60]), .A2 (Res_in[60]));
AOI21_X1 i_472 (.ZN (n_418), .A (n_421), .B1 (carry_in[60]), .B2 (Res_in[60]));
XOR2_X2 i_471 (.Z (Res_out[59]), .A (n_414), .B (n_417));
NAND2_X1 i_470 (.ZN (n_417), .A1 (n_415), .A2 (n_416));
NAND2_X1 i_469 (.ZN (n_416), .A1 (carry_in[59]), .A2 (Res_in[59]));
INV_X1 i_468 (.ZN (n_415), .A (n_409));
NAND2_X2 i_467 (.ZN (n_414), .A1 (n_412), .A2 (n_413));
INV_X1 i_466 (.ZN (n_413), .A (n_408));
NAND3_X2 i_465 (.ZN (n_412), .A1 (n_411), .A2 (sgo__sro_n174), .A3 (n_410));
INV_X2 i_464 (.ZN (n_411), .A (n_403));
AND3_X1 i_463 (.ZN (n_410), .A1 (n_396), .A2 (n_397), .A3 (n_401));
NOR2_X1 i_462 (.ZN (n_409), .A1 (carry_in[59]), .A2 (Res_in[59]));
AOI21_X1 i_461 (.ZN (n_408), .A (n_407), .B1 (n_400), .B2 (n_396));
INV_X1 i_460 (.ZN (n_407), .A (n_401));
XNOR2_X2 i_459 (.ZN (Res_out[58]), .A (slo__mro_n397), .B (n_406));
NAND2_X1 i_458 (.ZN (n_406), .A1 (n_400), .A2 (n_401));
XNOR2_X2 slo__sro_c773 (.ZN (Res_out[32]), .A (n_200), .B (slo__sro_n469));
OR2_X1 slo__mro_c750 (.ZN (n_56), .A1 (Res_in[17]), .A2 (carry_in[17]));
NAND2_X4 i_455 (.ZN (n_403), .A1 (n_364), .A2 (n_394));
INV_X4 i_454 (.ZN (n_402), .A (sgo__sro_n174));
NAND2_X1 i_453 (.ZN (n_401), .A1 (carry_in[58]), .A2 (Res_in[58]));
OR2_X1 i_452 (.ZN (n_400), .A1 (carry_in[58]), .A2 (Res_in[58]));
INV_X2 i_451 (.ZN (n_399), .A (sgo__sro_n74));
XNOR2_X2 i_450 (.ZN (Res_out[57]), .A (n_395), .B (n_398));
NAND2_X1 i_449 (.ZN (n_398), .A1 (n_396), .A2 (n_397));
NAND2_X1 i_448 (.ZN (n_397), .A1 (carry_in[57]), .A2 (Res_in[57]));
OR2_X1 i_447 (.ZN (n_396), .A1 (carry_in[57]), .A2 (Res_in[57]));
NAND3_X4 i_446 (.ZN (n_395), .A1 (sgo__sro_n174), .A2 (n_364), .A3 (n_394));
OAI21_X2 i_445 (.ZN (n_394), .A (n_356), .B1 (n_392), .B2 (n_393));
NAND2_X1 i_444 (.ZN (n_393), .A1 (n_388), .A2 (n_339));
INV_X1 CLOCK_slo__mro_c1948 (.ZN (CLOCK_slo__mro_n1455), .A (n_331));
INV_X1 i_442 (.ZN (n_389), .A (n_337));
NAND2_X1 i_441 (.ZN (n_388), .A1 (carry_in[56]), .A2 (Res_in[56]));
AOI21_X2 slo__c840 (.ZN (slo__n536), .A (n_103), .B1 (n_110), .B2 (n_373));
NAND2_X4 i_439 (.ZN (n_386), .A1 (n_378), .A2 (n_384));
INV_X4 i_438 (.ZN (n_384), .A (n_383));
OAI21_X2 i_437 (.ZN (n_383), .A (n_270), .B1 (n_381), .B2 (n_382));
INV_X1 i_436 (.ZN (n_382), .A (n_272));
AOI21_X2 i_435 (.ZN (n_381), .A (n_111), .B1 (n_372), .B2 (n_7));
AND2_X1 sgo__sro_c11 (.ZN (sgo__sro_n11), .A1 (Res_in[32]), .A2 (carry_in[32]));
NAND2_X1 i_433 (.ZN (n_379), .A1 (carry_in[39]), .A2 (Res_in[39]));
OAI21_X2 i_432 (.ZN (n_378), .A (n_375), .B1 (n_371), .B2 (sgo__sro_n74));
NAND2_X4 sgo__sro_c174 (.ZN (sgo__sro_n110), .A1 (n_66), .A2 (n_61));
INV_X4 i_430 (.ZN (n_376), .A (n_115));
AND3_X2 i_429 (.ZN (n_375), .A1 (n_372), .A2 (n_373), .A3 (n_272));
OR2_X1 i_428 (.ZN (n_373), .A1 (carry_in[37]), .A2 (Res_in[37]));
AND2_X4 i_427 (.ZN (n_372), .A1 (n_274), .A2 (n_267));
OAI21_X2 i_426 (.ZN (n_371), .A (n_368), .B1 (n_230), .B2 (slo__xsl_n558));
OR2_X2 slo__xsl_c914 (.ZN (n_329), .A1 (Res_in[44]), .A2 (carry_in[44]));
NOR2_X4 sgo__sro_c113 (.ZN (sgo__sro_n74), .A1 (n_376), .A2 (sgo__sro_n75));
AOI22_X2 i_423 (.ZN (n_368), .A1 (n_367), .A2 (n_251), .B1 (carry_in[36]), .B2 (Res_in[36]));
OAI21_X2 i_422 (.ZN (n_367), .A (n_255), .B1 (n_365), .B2 (CLOCK_slo__sro_n1317));
INV_X1 CLOCK_slo__sro_c1807 (.ZN (CLOCK_slo__sro_n1333), .A (n_245));
AOI22_X2 i_420 (.ZN (n_365), .A1 (Res_in[33]), .A2 (carry_in[33]), .B1 (carry_in[34]), .B2 (Res_in[34]));
OAI21_X4 i_419 (.ZN (n_364), .A (n_363), .B1 (n_357), .B2 (n_362));
AND4_X2 i_418 (.ZN (n_363), .A1 (n_355), .A2 (n_356), .A3 (n_341), .A4 (n_337));
NAND2_X4 i_417 (.ZN (n_362), .A1 (n_361), .A2 (n_307));
OAI21_X4 i_416 (.ZN (n_361), .A (n_308), .B1 (n_360), .B2 (n_358));
AOI21_X2 i_415 (.ZN (n_360), .A (n_359), .B1 (n_301), .B2 (n_312));
NAND2_X4 i_414 (.ZN (n_359), .A1 (n_302), .A2 (n_305));
INV_X1 i_413 (.ZN (n_358), .A (n_304));
AOI21_X4 i_412 (.ZN (n_357), .A (n_349), .B1 (n_321), .B2 (n_315));
OR2_X1 i_411 (.ZN (n_356), .A1 (carry_in[56]), .A2 (Res_in[56]));
INV_X1 i_410 (.ZN (n_355), .A (n_354));
NOR2_X1 i_409 (.ZN (n_354), .A1 (carry_in[55]), .A2 (Res_in[55]));
NAND2_X2 slo__sro_c966 (.ZN (n_290), .A1 (Res_in[47]), .A2 (carry_in[47]));
AND3_X4 i_407 (.ZN (n_352), .A1 (n_330), .A2 (n_277), .A3 (n_329));
NAND2_X4 i_406 (.ZN (n_351), .A1 (n_322), .A2 (n_352));
INV_X4 i_405 (.ZN (n_350), .A (n_351));
NAND4_X4 i_404 (.ZN (n_349), .A1 (n_313), .A2 (n_302), .A3 (n_305), .A4 (CLOCK_slo__n1604));
NAND2_X4 CLOCK_slo__mro_c1951 (.ZN (n_128), .A1 (CLOCK_slo__mro_n1454), .A2 (CLOCK_slo__mro_n1453));
NOR2_X2 i_402 (.ZN (n_347), .A1 (n_351), .A2 (n_349));
INV_X1 i_401 (.ZN (n_346), .A (n_336));
NAND2_X1 i_400 (.ZN (n_345), .A1 (carry_in[53]), .A2 (Res_in[53]));
INV_X1 i_399 (.ZN (n_344), .A (n_345));
NOR2_X1 i_398 (.ZN (n_343), .A1 (n_346), .A2 (n_344));
NOR2_X2 i_397 (.ZN (n_342), .A1 (carry_in[53]), .A2 (Res_in[53]));
INV_X2 i_396 (.ZN (n_341), .A (n_342));
NOR3_X1 i_395 (.ZN (n_340), .A1 (n_346), .A2 (n_344), .A3 (n_342));
NAND2_X1 i_394 (.ZN (n_339), .A1 (carry_in[55]), .A2 (Res_in[55]));
AND3_X1 i_393 (.ZN (n_338), .A1 (n_337), .A2 (n_340), .A3 (n_339));
OR2_X1 i_392 (.ZN (n_337), .A1 (carry_in[54]), .A2 (Res_in[54]));
NAND2_X1 i_391 (.ZN (n_336), .A1 (carry_in[54]), .A2 (Res_in[54]));
NAND2_X1 i_390 (.ZN (n_335), .A1 (n_337), .A2 (n_336));
INV_X1 i_389 (.ZN (n_334), .A (n_335));
INV_X1 i_388 (.ZN (n_333), .A (n_280));
INV_X1 i_387 (.ZN (n_332), .A (n_295));
NAND2_X1 i_386 (.ZN (n_331), .A1 (Res_in[44]), .A2 (carry_in[44]));
AOI21_X4 i_385 (.ZN (n_330), .A (n_281), .B1 (n_287), .B2 (n_286));
NOR2_X2 CLOCK_sgo__c1560 (.ZN (CLOCK_sgo__n1177), .A1 (Res_in[51]), .A2 (carry_in[51]));
NAND2_X2 i_383 (.ZN (n_328), .A1 (n_276), .A2 (CLOCK_slo__n1548));
AOI21_X2 i_382 (.ZN (n_327), .A (n_333), .B1 (n_330), .B2 (n_328));
OAI21_X1 i_381 (.ZN (n_326), .A (n_331), .B1 (n_327), .B2 (slo__xsl_n594));
NOR2_X2 i_380 (.ZN (n_325), .A1 (Res_in[48]), .A2 (carry_in[48]));
INV_X2 i_379 (.ZN (n_324), .A (n_325));
NAND3_X4 i_378 (.ZN (n_323), .A1 (n_296), .A2 (n_291), .A3 (n_324));
NOR2_X4 i_377 (.ZN (n_322), .A1 (n_323), .A2 (n_295));
NAND2_X2 i_376 (.ZN (n_321), .A1 (slo__n543), .A2 (n_322));
NAND2_X1 i_375 (.ZN (n_320), .A1 (Res_in[48]), .A2 (carry_in[48]));
NAND2_X2 i_374 (.ZN (n_319), .A1 (Res_in[45]), .A2 (carry_in[45]));
INV_X2 i_373 (.ZN (n_318), .A (n_319));
AOI21_X2 i_372 (.ZN (n_317), .A (n_318), .B1 (Res_in[46]), .B2 (carry_in[46]));
INV_X1 sgo__sro_c515 (.ZN (sgo__sro_n303), .A (n_308));
INV_X2 i_370 (.ZN (n_315), .A (n_316));
AOI21_X1 i_369 (.ZN (n_314), .A (n_316), .B1 (n_326), .B2 (n_322));
OR2_X2 i_368 (.ZN (n_313), .A1 (carry_in[49]), .A2 (Res_in[49]));
NAND2_X1 i_367 (.ZN (n_312), .A1 (carry_in[49]), .A2 (Res_in[49]));
NAND3_X1 i_366 (.ZN (n_311), .A1 (n_301), .A2 (n_312), .A3 (n_313));
NAND2_X1 i_365 (.ZN (n_310), .A1 (n_302), .A2 (n_304));
NOR2_X1 i_364 (.ZN (n_309), .A1 (n_311), .A2 (n_310));
OR2_X1 i_363 (.ZN (n_308), .A1 (carry_in[52]), .A2 (Res_in[52]));
NAND2_X1 i_362 (.ZN (n_307), .A1 (carry_in[52]), .A2 (Res_in[52]));
NAND2_X1 i_361 (.ZN (n_306), .A1 (n_308), .A2 (n_307));
XNOR2_X2 CLOCK_slo__sro_c1808 (.ZN (Res_out[34]), .A (n_248), .B (CLOCK_slo__sro_n1333));
NAND2_X1 i_359 (.ZN (n_304), .A1 (Res_in[51]), .A2 (carry_in[51]));
AND2_X1 i_358 (.ZN (n_303), .A1 (n_305), .A2 (n_304));
OR2_X4 i_357 (.ZN (n_302), .A1 (Res_in[50]), .A2 (carry_in[50]));
NAND2_X1 i_356 (.ZN (n_301), .A1 (Res_in[50]), .A2 (carry_in[50]));
AND2_X1 i_355 (.ZN (n_300), .A1 (n_302), .A2 (n_301));
INV_X1 i_354 (.ZN (n_299), .A (n_290));
NAND2_X1 i_353 (.ZN (n_298), .A1 (Res_in[46]), .A2 (carry_in[46]));
NOR2_X2 i_352 (.ZN (n_297), .A1 (Res_in[46]), .A2 (carry_in[46]));
INV_X2 i_351 (.ZN (n_296), .A (n_297));
NOR2_X2 i_350 (.ZN (n_295), .A1 (Res_in[45]), .A2 (carry_in[45]));
OAI21_X1 i_349 (.ZN (n_294), .A (n_298), .B1 (n_297), .B2 (n_295));
OAI21_X1 i_348 (.ZN (n_293), .A (n_291), .B1 (n_299), .B2 (n_294));
INV_X1 i_347 (.ZN (n_292), .A (n_293));
OR2_X2 i_346 (.ZN (n_291), .A1 (Res_in[47]), .A2 (carry_in[47]));
OR2_X2 CLOCK_slo__sro_c1797 (.ZN (CLOCK_slo__sro_n1310), .A1 (n_242), .A2 (n_303));
NAND2_X1 i_344 (.ZN (n_289), .A1 (n_291), .A2 (n_290));
INV_X1 i_343 (.ZN (n_288), .A (n_289));
INV_X1 i_342 (.ZN (n_287), .A (carry_in[42]));
INV_X1 i_341 (.ZN (n_286), .A (Res_in[42]));
NAND2_X1 i_340 (.ZN (n_285), .A1 (n_287), .A2 (n_286));
NAND2_X1 i_339 (.ZN (n_284), .A1 (carry_in[42]), .A2 (Res_in[42]));
NAND2_X1 i_338 (.ZN (n_283), .A1 (n_285), .A2 (n_284));
AND3_X1 i_337 (.ZN (n_282), .A1 (n_285), .A2 (n_284), .A3 (n_280));
NOR2_X2 i_336 (.ZN (n_281), .A1 (Res_in[43]), .A2 (carry_in[43]));
NAND2_X1 i_335 (.ZN (n_280), .A1 (carry_in[43]), .A2 (Res_in[43]));
AOI21_X1 i_334 (.ZN (n_279), .A (n_281), .B1 (carry_in[43]), .B2 (Res_in[43]));
INV_X1 i_333 (.ZN (n_278), .A (n_279));
OR2_X2 i_332 (.ZN (n_277), .A1 (Res_in[41]), .A2 (carry_in[41]));
NOR2_X4 slo__sro_c944 (.ZN (n_250), .A1 (Res_in[36]), .A2 (carry_in[36]));
NAND2_X1 i_330 (.ZN (n_275), .A1 (n_277), .A2 (CLOCK_opt_ipo_n1068));
NAND2_X1 CLOCK_slo__c2060 (.ZN (CLOCK_slo__n1548), .A1 (carry_in[42]), .A2 (Res_in[42]));
OR2_X2 i_327 (.ZN (n_272), .A1 (Res_in[40]), .A2 (carry_in[40]));
NAND2_X1 i_326 (.ZN (n_270), .A1 (Res_in[40]), .A2 (carry_in[40]));
NAND2_X1 i_325 (.ZN (n_268), .A1 (n_272), .A2 (n_270));
INV_X1 slo__xsl_c911 (.ZN (slo__xsl_n594), .A (n_329));
OAI21_X2 slo__c847 (.ZN (slo__n543), .A (n_331), .B1 (n_327), .B2 (slo__xsl_n594));
NAND2_X2 slo__mro_c683 (.ZN (slo__mro_n397), .A1 (n_404), .A2 (n_397));
AOI21_X1 i_321 (.ZN (n_265), .A (n_250), .B1 (Res_in[36]), .B2 (carry_in[36]));
OAI21_X2 slo__mro_c682 (.ZN (n_404), .A (n_396), .B1 (n_403), .B2 (n_402));
NOR2_X4 sgo__sro_c111 (.ZN (sgo__sro_n76), .A1 (n_231), .A2 (n_159));
INV_X1 i_318 (.ZN (n_259), .A (n_255));
NAND2_X1 i_317 (.ZN (n_255), .A1 (Res_in[35]), .A2 (carry_in[35]));
OAI21_X4 i_316 (.ZN (n_254), .A (n_246), .B1 (n_248), .B2 (n_253));
INV_X1 i_315 (.ZN (n_253), .A (n_247));
NOR2_X4 i_314 (.ZN (n_252), .A1 (Res_in[35]), .A2 (carry_in[35]));
INV_X1 i_313 (.ZN (n_251), .A (n_250));
NAND2_X1 slo__c958 (.ZN (slo__n626), .A1 (Res_in[38]), .A2 (carry_in[38]));
INV_X1 i_311 (.ZN (n_249), .A (n_243));
AOI21_X2 i_310 (.ZN (n_248), .A (n_249), .B1 (n_235), .B2 (n_241));
OR2_X1 i_309 (.ZN (n_247), .A1 (carry_in[34]), .A2 (Res_in[34]));
NAND2_X1 i_308 (.ZN (n_246), .A1 (carry_in[34]), .A2 (Res_in[34]));
NAND2_X1 i_307 (.ZN (n_245), .A1 (n_247), .A2 (n_246));
AND2_X1 CLOCK_slo__sro_c1830 (.ZN (CLOCK_slo__sro_n1364), .A1 (n_167), .A2 (n_319));
XNOR2_X1 i_305 (.ZN (Res_out[33]), .A (n_235), .B (n_244));
NAND2_X1 i_304 (.ZN (n_244), .A1 (n_241), .A2 (n_243));
NAND2_X1 i_303 (.ZN (n_243), .A1 (Res_in[33]), .A2 (carry_in[33]));
INV_X1 i_302 (.ZN (n_241), .A (n_239));
NOR2_X2 i_301 (.ZN (n_239), .A1 (Res_in[33]), .A2 (carry_in[33]));
OAI21_X2 i_300 (.ZN (n_235), .A (n_230), .B1 (n_232), .B2 (n_231));
NAND2_X1 i_299 (.ZN (n_232), .A1 (n_115), .A2 (n_168));
NAND3_X4 i_298 (.ZN (n_231), .A1 (CLOCK_slo__n1598), .A2 (n_160), .A3 (n_175));
NAND2_X1 sgo__sro_c240 (.ZN (sgo__sro_n146), .A1 (n_278), .A2 (n_284));
AND2_X2 i_296 (.ZN (n_229), .A1 (n_187), .A2 (n_191));
INV_X2 sgo__sro_c175 (.ZN (sgo__sro_n109), .A (sgo__sro_n110));
NAND3_X2 i_294 (.ZN (n_214), .A1 (Res_in[29]), .A2 (carry_in[29]), .A3 (n_175));
NAND3_X2 i_293 (.ZN (n_204), .A1 (opt_ipo_n883), .A2 (n_160), .A3 (n_175));
OAI21_X2 sgo__sro_c80 (.ZN (sgo__sro_n48), .A (sgo__sro_n49), .B1 (n_210), .B2 (n_342));
OAI21_X4 slo__c778 (.ZN (slo__n476), .A (n_49), .B1 (n_53), .B2 (n_54));
OAI21_X2 i_290 (.ZN (n_200), .A (n_185), .B1 (n_188), .B2 (CLOCK_slo__xsl_n1578));
AOI21_X1 i_289 (.ZN (n_199), .A (CLOCK_slo__xsl_n1508), .B1 (Res_in[32]), .B2 (carry_in[32]));
NAND2_X2 CLOCK_slo__c2049 (.ZN (CLOCK_slo__n1537), .A1 (n_271), .A2 (n_314));
AND2_X4 CLOCK_slo__c2120 (.ZN (CLOCK_slo__n1598), .A1 (n_187), .A2 (n_191));
INV_X1 i_286 (.ZN (n_189), .A (n_174));
AOI21_X4 i_285 (.ZN (n_188), .A (n_189), .B1 (n_171), .B2 (n_175));
OR2_X2 CLOCK_slo__c2129 (.ZN (CLOCK_slo__n1604), .A1 (carry_in[52]), .A2 (Res_in[52]));
NAND2_X1 i_282 (.ZN (n_185), .A1 (Res_in[31]), .A2 (carry_in[31]));
NAND2_X1 i_281 (.ZN (n_182), .A1 (n_187), .A2 (n_185));
OR2_X4 CLOCK_slo__c2001 (.ZN (n_274), .A1 (Res_in[39]), .A2 (carry_in[39]));
INV_X1 i_279 (.ZN (n_179), .A (n_160));
INV_X1 slo__xsl_c795 (.ZN (slo__xsl_n495), .A (n_267));
NAND2_X1 i_277 (.ZN (n_174), .A1 (Res_in[30]), .A2 (carry_in[30]));
OAI21_X2 i_276 (.ZN (n_171), .A (n_161), .B1 (n_169), .B2 (n_179));
NAND2_X1 i_275 (.ZN (n_170), .A1 (n_175), .A2 (n_174));
XNOR2_X1 i_274 (.ZN (Res_out[30]), .A (n_171), .B (n_170));
XOR2_X1 i_273 (.Z (Res_out[29]), .A (n_162), .B (n_169));
AOI21_X1 i_272 (.ZN (n_169), .A (opt_ipo_n883), .B1 (n_115), .B2 (n_168));
INV_X1 i_271 (.ZN (n_168), .A (n_159));
NAND2_X4 CLOCK_slo__sro_c1798 (.ZN (Res_out[51]), .A1 (n_240), .A2 (CLOCK_slo__sro_n1310));
NAND2_X1 i_269 (.ZN (n_162), .A1 (n_160), .A2 (n_161));
NAND2_X1 i_268 (.ZN (n_161), .A1 (Res_in[29]), .A2 (carry_in[29]));
OR2_X4 i_267 (.ZN (n_160), .A1 (Res_in[29]), .A2 (carry_in[29]));
NAND4_X2 i_266 (.ZN (n_159), .A1 (n_152), .A2 (n_135), .A3 (n_148), .A4 (n_119));
AOI21_X4 i_265 (.ZN (n_158), .A (n_153), .B1 (n_157), .B2 (n_148));
OAI21_X2 i_264 (.ZN (n_157), .A (n_136), .B1 (n_156), .B2 (n_155));
NAND2_X4 i_263 (.ZN (n_156), .A1 (n_135), .A2 (n_152));
AOI22_X2 i_262 (.ZN (n_155), .A1 (Res_in[25]), .A2 (carry_in[25]), .B1 (Res_in[26]), .B2 (carry_in[26]));
INV_X1 i_261 (.ZN (n_153), .A (n_143));
INV_X4 i_260 (.ZN (n_152), .A (n_133));
INV_X1 i_259 (.ZN (n_149), .A (n_136));
OR2_X2 i_258 (.ZN (n_148), .A1 (carry_in[28]), .A2 (Res_in[28]));
NAND2_X1 i_257 (.ZN (n_143), .A1 (carry_in[28]), .A2 (Res_in[28]));
AOI21_X1 i_256 (.ZN (n_139), .A (n_149), .B1 (n_134), .B2 (n_135));
NAND2_X1 i_255 (.ZN (n_138), .A1 (n_148), .A2 (n_143));
XOR2_X2 i_254 (.Z (Res_out[28]), .A (n_139), .B (n_138));
XNOR2_X1 i_253 (.ZN (Res_out[27]), .A (n_134), .B (n_137));
NAND2_X1 i_252 (.ZN (n_137), .A1 (n_135), .A2 (n_136));
NAND2_X1 i_251 (.ZN (n_136), .A1 (Res_in[27]), .A2 (carry_in[27]));
OR2_X4 i_250 (.ZN (n_135), .A1 (Res_in[27]), .A2 (carry_in[27]));
OAI21_X2 i_249 (.ZN (n_134), .A (n_86), .B1 (n_124), .B2 (n_133));
NOR2_X4 i_248 (.ZN (n_133), .A1 (Res_in[26]), .A2 (carry_in[26]));
AOI21_X1 i_247 (.ZN (n_124), .A (n_123), .B1 (n_115), .B2 (n_119));
INV_X1 i_246 (.ZN (n_123), .A (n_122));
NAND2_X1 i_245 (.ZN (n_122), .A1 (Res_in[25]), .A2 (carry_in[25]));
OR2_X2 i_244 (.ZN (n_119), .A1 (Res_in[25]), .A2 (carry_in[25]));
AOI21_X4 i_243 (.ZN (n_115), .A (n_87), .B1 (n_105), .B2 (n_113));
AOI21_X2 i_242 (.ZN (n_113), .A (n_112), .B1 (Res_in[23]), .B2 (carry_in[23]));
INV_X1 i_241 (.ZN (n_112), .A (n_93));
NAND3_X2 i_240 (.ZN (n_105), .A1 (n_94), .A2 (n_95), .A3 (n_104));
OR2_X2 i_239 (.ZN (n_104), .A1 (Res_in[22]), .A2 (carry_in[22]));
OR2_X2 i_238 (.ZN (n_95), .A1 (Res_in[23]), .A2 (carry_in[23]));
NAND3_X2 i_237 (.ZN (n_94), .A1 (n_91), .A2 (n_78), .A3 (n_92));
NAND2_X1 i_236 (.ZN (n_93), .A1 (Res_in[24]), .A2 (carry_in[24]));
NAND2_X2 i_235 (.ZN (n_92), .A1 (Res_in[22]), .A2 (carry_in[22]));
OAI21_X2 i_234 (.ZN (n_91), .A (n_77), .B1 (n_89), .B2 (n_90));
INV_X1 i_233 (.ZN (n_90), .A (n_73));
NAND2_X2 i_232 (.ZN (n_89), .A1 (slo__n516), .A2 (n_81));
INV_X1 i_231 (.ZN (n_88), .A (n_87));
NOR2_X1 i_230 (.ZN (n_87), .A1 (Res_in[24]), .A2 (carry_in[24]));
NAND2_X1 i_229 (.ZN (n_86), .A1 (Res_in[26]), .A2 (carry_in[26]));
XNOR2_X1 i_228 (.ZN (Res_out[21]), .A (n_84), .B (n_85));
NAND2_X1 i_227 (.ZN (n_85), .A1 (n_77), .A2 (n_78));
NAND3_X1 i_226 (.ZN (n_84), .A1 (n_81), .A2 (n_73), .A3 (sgo__sro_n108));
OAI21_X2 sgo__sro_c242 (.ZN (sgo__sro_n144), .A (sgo__sro_n145), .B1 (n_118), .B2 (n_131));
INV_X4 i_224 (.ZN (n_82), .A (n_63));
OAI211_X2 i_223 (.ZN (n_81), .A (n_66), .B (n_74), .C1 (n_79), .C2 (n_80));
NAND2_X1 i_222 (.ZN (n_80), .A1 (n_60), .A2 (n_67));
AOI21_X2 i_221 (.ZN (n_79), .A (n_57), .B1 (n_65), .B2 (n_64));
NAND2_X2 i_220 (.ZN (n_78), .A1 (Res_in[21]), .A2 (carry_in[21]));
OR2_X2 i_219 (.ZN (n_77), .A1 (Res_in[21]), .A2 (carry_in[21]));
INV_X1 i_218 (.ZN (n_75), .A (n_67));
OR2_X4 i_217 (.ZN (n_74), .A1 (Res_in[20]), .A2 (carry_in[20]));
NAND2_X1 i_216 (.ZN (n_73), .A1 (Res_in[20]), .A2 (carry_in[20]));
NAND2_X1 i_215 (.ZN (n_72), .A1 (n_74), .A2 (n_73));
AOI21_X1 i_214 (.ZN (n_71), .A (n_75), .B1 (n_70), .B2 (n_66));
XOR2_X2 i_213 (.Z (Res_out[20]), .A (n_72), .B (n_71));
XNOR2_X1 i_212 (.ZN (Res_out[19]), .A (n_68), .B (n_70));
NAND2_X1 i_211 (.ZN (n_70), .A1 (n_69), .A2 (n_60));
NAND2_X1 i_210 (.ZN (n_69), .A1 (n_62), .A2 (n_61));
NAND2_X1 i_209 (.ZN (n_68), .A1 (n_66), .A2 (n_67));
NAND2_X2 i_208 (.ZN (n_67), .A1 (Res_in[19]), .A2 (carry_in[19]));
OAI21_X1 sgo__sro_c342 (.ZN (sgo__sro_n211), .A (n_320), .B1 (n_290), .B2 (n_325));
INV_X2 i_206 (.ZN (n_65), .A (Res_in[18]));
INV_X1 i_205 (.ZN (n_64), .A (carry_in[18]));
NAND2_X4 i_204 (.ZN (n_63), .A1 (slo__n476), .A2 (n_56));
NAND2_X1 i_203 (.ZN (n_62), .A1 (n_57), .A2 (n_63));
NAND2_X2 i_202 (.ZN (n_61), .A1 (n_65), .A2 (n_64));
NAND2_X2 i_201 (.ZN (n_60), .A1 (Res_in[18]), .A2 (carry_in[18]));
NAND2_X1 i_200 (.ZN (n_59), .A1 (n_61), .A2 (n_60));
XNOR2_X1 i_199 (.ZN (Res_out[18]), .A (n_62), .B (n_59));
XNOR2_X1 i_198 (.ZN (Res_out[17]), .A (n_55), .B (n_58));
NAND2_X1 i_197 (.ZN (n_58), .A1 (n_56), .A2 (n_57));
NAND2_X2 i_196 (.ZN (n_57), .A1 (Res_in[17]), .A2 (carry_in[17]));
OAI21_X2 slo__sro_c768 (.ZN (n_316), .A (sgo__sro_n210), .B1 (n_317), .B2 (n_323));
OAI21_X1 i_194 (.ZN (n_55), .A (n_49), .B1 (n_53), .B2 (n_54));
OAI21_X4 i_193 (.ZN (n_54), .A (n_50), .B1 (Res_in[15]), .B2 (carry_in[15]));
AOI22_X4 i_192 (.ZN (n_53), .A1 (n_51), .A2 (opt_ipo_n987), .B1 (Res_in[15]), .B2 (carry_in[15]));
AND2_X1 sgo__sro_c79 (.ZN (sgo__sro_n49), .A1 (n_335), .A2 (n_345));
NAND3_X2 i_190 (.ZN (n_51), .A1 (n_33), .A2 (n_32), .A3 (n_30));
OR2_X4 i_189 (.ZN (n_50), .A1 (Res_in[16]), .A2 (carry_in[16]));
NAND2_X1 i_188 (.ZN (n_49), .A1 (Res_in[16]), .A2 (carry_in[16]));
NOR2_X1 i_187 (.ZN (n_48), .A1 (Res_in[14]), .A2 (carry_in[14]));
INV_X1 CLOCK_slo__sro_c1859 (.ZN (CLOCK_slo__sro_n1388), .A (n_389));
OAI21_X2 i_185 (.ZN (n_33), .A (n_13), .B1 (Res_in[13]), .B2 (carry_in[13]));
NAND2_X1 i_184 (.ZN (n_32), .A1 (Res_in[13]), .A2 (carry_in[13]));
NAND2_X1 i_183 (.ZN (n_31), .A1 (n_33), .A2 (n_32));
NAND2_X1 i_182 (.ZN (n_30), .A1 (Res_in[14]), .A2 (carry_in[14]));
AOI22_X1 i_181 (.ZN (n_29), .A1 (Res_in[14]), .A2 (carry_in[14]), .B1 (opt_ipo_n987), .B2 (n_31));
OR2_X1 i_180 (.ZN (n_28), .A1 (Res_in[15]), .A2 (carry_in[15]));
NAND2_X1 i_179 (.ZN (n_27), .A1 (Res_in[15]), .A2 (carry_in[15]));
NAND2_X1 i_178 (.ZN (n_26), .A1 (n_28), .A2 (n_27));
XOR2_X1 i_177 (.Z (Res_out[15]), .A (n_29), .B (n_26));
OR2_X2 i_176 (.ZN (n_25), .A1 (Res_in[11]), .A2 (carry_in[11]));
OR2_X1 i_175 (.ZN (n_24), .A1 (Res_in[12]), .A2 (carry_in[12]));
NAND2_X2 i_174 (.ZN (n_23), .A1 (Res_in[9]), .A2 (carry_in[9]));
INV_X1 i_173 (.ZN (n_22), .A (n_23));
NOR2_X2 i_172 (.ZN (n_21), .A1 (Res_in[10]), .A2 (carry_in[10]));
INV_X1 i_171 (.ZN (n_20), .A (n_21));
NAND2_X2 i_170 (.ZN (n_19), .A1 (Res_in[11]), .A2 (carry_in[11]));
NAND2_X2 i_169 (.ZN (n_17), .A1 (Res_in[10]), .A2 (carry_in[10]));
NAND2_X1 i_168 (.ZN (n_16), .A1 (Res_in[12]), .A2 (carry_in[12]));
OAI211_X2 i_167 (.ZN (n_15), .A (n_19), .B (n_17), .C1 (n_23), .C2 (n_21));
NAND3_X1 i_166 (.ZN (n_14), .A1 (n_15), .A2 (n_24), .A3 (n_25));
NAND2_X2 i_165 (.ZN (n_13), .A1 (n_14), .A2 (n_16));
XOR2_X1 i_164 (.Z (n_12), .A (Res_in[13]), .B (carry_in[13]));
XOR2_X1 i_163 (.Z (Res_out[13]), .A (n_13), .B (n_12));
XOR2_X1 i_162 (.Z (Res_out[9]), .A (Res_in[9]), .B (carry_in[9]));
AOI21_X1 i_161 (.ZN (n_385), .A (n_409), .B1 (n_408), .B2 (n_416));
OAI21_X2 i_160 (.ZN (n_374), .A (n_385), .B1 (n_395), .B2 (n_263));
XNOR2_X2 i_159 (.ZN (Res_out[60]), .A (n_374), .B (n_418));
NAND2_X2 i_158 (.ZN (n_233), .A1 (n_386), .A2 (n_347));
NOR2_X2 i_157 (.ZN (n_238), .A1 (n_357), .A2 (n_362));
NAND2_X2 i_156 (.ZN (n_211), .A1 (n_233), .A2 (n_238));
XNOR2_X2 i_155 (.ZN (Res_out[53]), .A (n_211), .B (n_207));
NAND2_X2 i_154 (.ZN (n_271), .A1 (n_386), .A2 (n_350));
NAND2_X2 i_153 (.ZN (n_184), .A1 (n_271), .A2 (n_314));
INV_X1 i_152 (.ZN (n_269), .A (n_184));
NAND2_X2 i_151 (.ZN (n_262), .A1 (n_269), .A2 (n_309));
NAND3_X2 i_150 (.ZN (n_261), .A1 (n_262), .A2 (n_306), .A3 (n_190));
NAND3_X4 slo__c825 (.ZN (slo__n516), .A1 (n_82), .A2 (sgo__sro_n109), .A3 (n_74));
NAND2_X1 i_148 (.ZN (n_257), .A1 (n_195), .A2 (n_301));
OAI21_X1 i_147 (.ZN (n_193), .A (n_305), .B1 (n_257), .B2 (n_358));
AND2_X1 slo__sro_c659 (.ZN (slo__sro_n375), .A1 (n_429), .A2 (n_425));
NAND2_X2 slo__sro_c850 (.ZN (n_276), .A1 (carry_in[41]), .A2 (Res_in[41]));
OAI21_X2 i_144 (.ZN (n_242), .A (n_257), .B1 (CLOCK_slo__n1537), .B2 (n_311));
NAND3_X1 i_143 (.ZN (n_240), .A1 (n_242), .A2 (n_305), .A3 (n_304));
OAI21_X4 CLOCK_slo__sro_c1803 (.ZN (CLOCK_slo__sro_n1317), .A (opt_ipo_n737), .B1 (Res_in[34]), .B2 (carry_in[34]));
INV_X1 i_141 (.ZN (n_236), .A (n_312));
INV_X4 opt_ipo_c1196 (.ZN (opt_ipo_n883), .A (n_158));
AOI21_X2 i_139 (.ZN (n_206), .A (n_236), .B1 (CLOCK_slo__n1537), .B2 (n_313));
NAND2_X1 i_138 (.ZN (n_205), .A1 (n_184), .A2 (n_313));
NAND3_X2 i_137 (.ZN (n_203), .A1 (n_205), .A2 (n_312), .A3 (n_300));
OAI21_X4 i_136 (.ZN (Res_out[50]), .A (n_203), .B1 (n_206), .B2 (n_300));
XNOR2_X2 i_135 (.ZN (Res_out[49]), .A (CLOCK_slo__n1537), .B (n_173));
INV_X1 i_134 (.ZN (n_183), .A (n_326));
NAND2_X2 i_133 (.ZN (n_181), .A1 (n_386), .A2 (n_352));
NAND2_X4 i_132 (.ZN (n_180), .A1 (n_181), .A2 (n_183));
OAI211_X1 i_131 (.ZN (n_202), .A (n_154), .B (n_292), .C1 (n_180), .C2 (n_163));
INV_X1 i_130 (.ZN (n_198), .A (n_163));
AOI21_X4 sgo__sro_c12 (.ZN (n_230), .A (sgo__sro_n11), .B1 (n_215), .B2 (n_229));
AOI21_X1 i_128 (.ZN (n_196), .A (n_293), .B1 (n_142), .B2 (n_198));
NAND2_X1 i_127 (.ZN (n_194), .A1 (n_324), .A2 (n_320));
OAI21_X2 i_126 (.ZN (Res_out[48]), .A (n_202), .B1 (n_196), .B2 (n_194));
XNOR2_X2 i_125 (.ZN (Res_out[45]), .A (n_180), .B (n_165));
NAND2_X4 i_124 (.ZN (n_178), .A1 (n_386), .A2 (n_277));
NAND2_X2 i_123 (.ZN (n_177), .A1 (n_178), .A2 (CLOCK_opt_ipo_n1068));
XNOR2_X2 i_122 (.ZN (Res_out[42]), .A (n_177), .B (n_283));
NAND2_X1 i_121 (.ZN (n_0), .A1 (Res_in[23]), .A2 (carry_in[23]));
INV_X1 i_120 (.ZN (n_237), .A (n_371));
INV_X1 i_119 (.ZN (n_172), .A (n_165));
INV_X1 CLOCK_slo__xsl_c2016 (.ZN (CLOCK_slo__xsl_n1508), .A (n_191));
NAND2_X1 i_117 (.ZN (n_391), .A1 (Res_in[38]), .A2 (carry_in[38]));
NAND2_X1 i_116 (.ZN (n_390), .A1 (Res_in[37]), .A2 (carry_in[37]));
NAND2_X1 i_115 (.ZN (n_7), .A1 (n_390), .A2 (slo__n626));
AOI21_X4 i_114 (.ZN (Res_out[63]), .A (n_436), .B1 (n_434), .B2 (n_433));
NOR2_X2 i_113 (.ZN (Res_out[62]), .A1 (n_432), .A2 (Res_out[63]));
NAND3_X1 i_112 (.ZN (n_263), .A1 (n_410), .A2 (n_400), .A3 (n_416));
NAND3_X1 i_111 (.ZN (n_228), .A1 (n_233), .A2 (n_238), .A3 (n_338));
AOI21_X1 i_110 (.ZN (n_227), .A (n_346), .B1 (n_341), .B2 (n_337));
AOI21_X1 i_109 (.ZN (n_226), .A (n_354), .B1 (n_227), .B2 (n_339));
NAND2_X1 i_108 (.ZN (n_225), .A1 (n_228), .A2 (n_226));
NAND3_X1 i_107 (.ZN (n_224), .A1 (n_225), .A2 (n_356), .A3 (n_388));
NAND2_X1 i_106 (.ZN (n_223), .A1 (n_356), .A2 (n_388));
NAND3_X1 i_105 (.ZN (n_222), .A1 (n_228), .A2 (n_223), .A3 (n_226));
NAND2_X2 i_104 (.ZN (Res_out[56]), .A1 (n_224), .A2 (n_222));
NAND3_X1 i_103 (.ZN (n_221), .A1 (n_233), .A2 (n_238), .A3 (n_340));
INV_X1 i_102 (.ZN (n_220), .A (n_221));
OAI211_X2 i_101 (.ZN (n_219), .A (n_355), .B (n_339), .C1 (n_220), .C2 (n_227));
INV_X1 i_100 (.ZN (n_218), .A (n_227));
NAND2_X1 i_99 (.ZN (n_217), .A1 (n_355), .A2 (n_339));
NAND3_X1 i_98 (.ZN (n_216), .A1 (n_221), .A2 (n_218), .A3 (n_217));
NAND2_X4 i_97 (.ZN (Res_out[55]), .A1 (n_219), .A2 (n_216));
AOI21_X2 i_96 (.ZN (n_213), .A (n_342), .B1 (n_233), .B2 (n_238));
OAI21_X1 i_95 (.ZN (n_212), .A (n_334), .B1 (n_213), .B2 (n_344));
INV_X1 i_94 (.ZN (n_210), .A (n_211));
NAND2_X2 sgo__sro_c112 (.ZN (sgo__sro_n75), .A1 (sgo__sro_n76), .A2 (n_370));
NAND2_X2 i_92 (.ZN (n_208), .A1 (sgo__sro_n48), .A2 (n_212));
INV_X4 i_91 (.ZN (Res_out[54]), .A (n_208));
NAND2_X1 i_90 (.ZN (n_207), .A1 (n_341), .A2 (n_345));
NAND2_X1 i_89 (.ZN (n_195), .A1 (n_313), .A2 (n_302));
INV_X1 i_88 (.ZN (n_190), .A (n_193));
INV_X1 sgo__sro_c241 (.ZN (sgo__sro_n145), .A (sgo__sro_n146));
NAND2_X1 i_86 (.ZN (n_173), .A1 (n_313), .A2 (n_312));
NAND2_X1 i_85 (.ZN (n_167), .A1 (n_296), .A2 (n_298));
INV_X1 i_84 (.ZN (n_166), .A (n_167));
NAND2_X1 i_83 (.ZN (n_165), .A1 (n_332), .A2 (n_319));
NAND3_X1 i_82 (.ZN (n_163), .A1 (n_166), .A2 (n_290), .A3 (n_172));
NAND2_X1 i_81 (.ZN (n_154), .A1 (n_324), .A2 (n_320));
NAND4_X1 i_80 (.ZN (n_151), .A1 (n_181), .A2 (n_183), .A3 (n_298), .A4 (n_172));
NAND2_X1 i_79 (.ZN (n_150), .A1 (n_151), .A2 (n_294));
NAND2_X1 i_78 (.ZN (n_147), .A1 (n_150), .A2 (n_288));
NAND3_X2 i_77 (.ZN (n_146), .A1 (n_151), .A2 (n_294), .A3 (n_289));
NAND2_X4 i_76 (.ZN (Res_out[47]), .A1 (n_147), .A2 (n_146));
AOI21_X1 i_75 (.ZN (n_145), .A (n_295), .B1 (n_181), .B2 (n_183));
OAI21_X1 i_74 (.ZN (n_144), .A (n_166), .B1 (n_145), .B2 (n_318));
INV_X2 i_73 (.ZN (n_142), .A (n_180));
INV_X1 CLOCK_slo__sro_c1858 (.ZN (CLOCK_slo__sro_n1389), .A (n_354));
NAND2_X1 i_71 (.ZN (n_140), .A1 (CLOCK_slo__sro_n1363), .A2 (n_144));
INV_X4 i_70 (.ZN (Res_out[46]), .A (n_140));
NAND3_X2 i_69 (.ZN (n_132), .A1 (n_178), .A2 (CLOCK_opt_ipo_n1068), .A3 (n_282));
INV_X1 i_68 (.ZN (n_131), .A (n_285));
OAI21_X1 i_67 (.ZN (n_130), .A (n_280), .B1 (n_131), .B2 (n_281));
INV_X1 CLOCK_slo__xsl_c2091 (.ZN (CLOCK_slo__xsl_n1578), .A (n_187));
NAND2_X1 i_64 (.ZN (n_127), .A1 (n_329), .A2 (n_331));
NAND3_X1 i_63 (.ZN (n_126), .A1 (n_132), .A2 (n_127), .A3 (n_130));
OR2_X4 CLOCK_slo__xsl_c2094 (.ZN (n_187), .A1 (carry_in[31]), .A2 (Res_in[31]));
INV_X1 i_61 (.ZN (n_125), .A (n_284));
AOI21_X1 i_60 (.ZN (n_121), .A (n_131), .B1 (n_178), .B2 (CLOCK_opt_ipo_n1068));
OAI21_X1 i_59 (.ZN (n_120), .A (n_279), .B1 (n_121), .B2 (n_125));
INV_X1 i_58 (.ZN (n_118), .A (n_177));
NOR2_X2 sgo__c303 (.ZN (sgo__n190), .A1 (Res_in[19]), .A2 (carry_in[19]));
NAND2_X2 i_56 (.ZN (n_116), .A1 (sgo__sro_n144), .A2 (n_120));
INV_X4 i_55 (.ZN (Res_out[43]), .A (n_116));
NAND2_X1 i_54 (.ZN (n_114), .A1 (n_378), .A2 (n_384));
XNOR2_X1 i_53 (.ZN (Res_out[41]), .A (n_114), .B (n_275));
INV_X1 i_52 (.ZN (n_111), .A (n_379));
NAND2_X2 i_51 (.ZN (n_110), .A1 (n_237), .A2 (n_399));
NAND2_X1 i_50 (.ZN (n_109), .A1 (n_110), .A2 (n_373));
NAND3_X1 i_49 (.ZN (n_108), .A1 (n_109), .A2 (n_391), .A3 (n_390));
AOI21_X1 i_48 (.ZN (n_107), .A (n_111), .B1 (n_108), .B2 (n_267));
OAI211_X2 i_47 (.ZN (n_106), .A (n_272), .B (n_270), .C1 (n_107), .C2 (opt_ipo_n1007));
INV_X1 i_46 (.ZN (n_103), .A (n_390));
AOI21_X1 i_45 (.ZN (n_102), .A (n_103), .B1 (n_110), .B2 (n_373));
AOI21_X2 i_44 (.ZN (n_101), .A (slo__xsl_n495), .B1 (slo__n536), .B2 (n_391));
OAI211_X1 i_43 (.ZN (n_100), .A (opt_ipo_n1006), .B (n_268), .C1 (n_101), .C2 (n_111));
NAND2_X4 i_42 (.ZN (Res_out[40]), .A1 (n_106), .A2 (n_100));
NAND2_X1 i_41 (.ZN (n_99), .A1 (opt_ipo_n1006), .A2 (n_379));
XNOR2_X2 i_40 (.ZN (Res_out[39]), .A (n_101), .B (n_99));
NAND2_X1 i_39 (.ZN (n_98), .A1 (n_267), .A2 (n_391));
XOR2_X2 i_38 (.Z (Res_out[38]), .A (n_102), .B (n_98));
NAND2_X1 i_37 (.ZN (n_97), .A1 (n_373), .A2 (n_390));
XOR2_X1 i_36 (.Z (n_96), .A (n_97), .B (n_110));
INV_X1 i_35 (.ZN (Res_out[37]), .A (n_96));
NAND2_X1 i_34 (.ZN (n_76), .A1 (opt_ipo_n737), .A2 (n_255));
XNOR2_X2 i_33 (.ZN (Res_out[35]), .A (n_254), .B (n_76));
NAND2_X1 i_32 (.ZN (n_46), .A1 (n_152), .A2 (n_86));
XNOR2_X1 i_31 (.ZN (n_45), .A (n_124), .B (n_46));
INV_X1 i_30 (.ZN (Res_out[26]), .A (n_45));
NAND2_X1 i_29 (.ZN (n_44), .A1 (n_119), .A2 (n_122));
XOR2_X1 i_28 (.Z (n_43), .A (n_44), .B (n_115));
INV_X1 i_27 (.ZN (Res_out[25]), .A (n_43));
NAND2_X1 i_26 (.ZN (n_42), .A1 (n_88), .A2 (n_93));
AND2_X1 i_25 (.ZN (n_41), .A1 (n_91), .A2 (n_78));
NAND2_X1 i_24 (.ZN (n_40), .A1 (n_41), .A2 (n_92));
NAND2_X1 i_23 (.ZN (n_39), .A1 (n_40), .A2 (n_104));
NAND2_X1 i_22 (.ZN (n_38), .A1 (n_39), .A2 (n_0));
NAND2_X1 i_21 (.ZN (n_37), .A1 (n_38), .A2 (n_95));
XOR2_X1 i_20 (.Z (Res_out[24]), .A (n_42), .B (n_37));
NAND2_X1 i_19 (.ZN (n_36), .A1 (n_95), .A2 (n_0));
XOR2_X1 i_18 (.Z (Res_out[23]), .A (n_36), .B (n_39));
NAND2_X1 i_17 (.ZN (n_35), .A1 (n_104), .A2 (n_92));
XNOR2_X1 i_16 (.ZN (n_34), .A (n_41), .B (n_35));
INV_X1 i_15 (.ZN (Res_out[22]), .A (n_34));
NAND2_X1 i_14 (.ZN (n_18), .A1 (n_50), .A2 (n_49));
NAND2_X1 i_13 (.ZN (n_11), .A1 (n_29), .A2 (n_27));
NAND2_X1 i_12 (.ZN (n_10), .A1 (n_11), .A2 (n_28));
XOR2_X1 i_11 (.Z (Res_out[16]), .A (n_18), .B (n_10));
NAND2_X1 i_10 (.ZN (n_8), .A1 (opt_ipo_n987), .A2 (n_30));
XNOR2_X1 i_9 (.ZN (Res_out[14]), .A (n_31), .B (n_8));
INV_X1 i_8 (.ZN (n_6), .A (n_19));
AOI21_X1 i_7 (.ZN (n_5), .A (n_21), .B1 (n_17), .B2 (n_23));
OAI21_X1 i_6 (.ZN (n_4), .A (n_25), .B1 (n_5), .B2 (n_6));
NAND2_X1 i_5 (.ZN (n_3), .A1 (n_24), .A2 (n_16));
XOR2_X1 i_4 (.Z (Res_out[12]), .A (n_3), .B (n_4));
NAND2_X1 i_3 (.ZN (n_2), .A1 (n_25), .A2 (n_19));
XNOR2_X1 i_2 (.ZN (Res_out[11]), .A (n_2), .B (n_5));
NAND2_X1 i_1 (.ZN (n_1), .A1 (n_20), .A2 (n_17));
XNOR2_X1 i_0 (.ZN (Res_out[10]), .A (n_1), .B (n_22));
NAND2_X1 sgo__sro_c34 (.ZN (sgo__sro_n26), .A1 (n_174), .A2 (n_185));
INV_X1 sgo__sro_c35 (.ZN (sgo__sro_n25), .A (sgo__sro_n26));
NAND3_X2 sgo__sro_c36 (.ZN (n_215), .A1 (n_204), .A2 (n_214), .A3 (sgo__sro_n25));
NAND3_X1 sgo__sro_c176 (.ZN (sgo__sro_n108), .A1 (n_82), .A2 (sgo__sro_n109), .A3 (n_74));
INV_X4 sgo__c305 (.ZN (n_66), .A (sgo__n190));
INV_X1 sgo__sro_c343 (.ZN (sgo__sro_n210), .A (sgo__sro_n211));
INV_X1 slo__sro_c772 (.ZN (slo__sro_n469), .A (n_199));
INV_X1 sgo__sro_c516 (.ZN (sgo__sro_n302), .A (n_307));
NOR2_X1 sgo__sro_c517 (.ZN (sgo__sro_n301), .A1 (sgo__sro_n303), .A2 (sgo__sro_n302));
NOR2_X2 CLOCK_slo__mro_c1950 (.ZN (CLOCK_slo__mro_n1453), .A1 (CLOCK_slo__mro_n1455), .A2 (CLOCK_slo__mro_n1456));
INV_X1 sgo__sro_c285 (.ZN (sgo__sro_n178), .A (n_363));
NOR2_X4 sgo__sro_c286 (.ZN (sgo__sro_n177), .A1 (sgo__sro_n178), .A2 (n_349));
NAND2_X4 sgo__sro_c287 (.ZN (sgo__sro_n176), .A1 (n_350), .A2 (sgo__sro_n177));
INV_X4 CLOCK_sgo__c1562 (.ZN (n_305), .A (CLOCK_sgo__n1177));
NAND2_X4 sgo__sro_c289 (.ZN (sgo__sro_n174), .A1 (n_386), .A2 (CLOCK_opt_ipo_n1035));
OAI21_X4 slo__sro_c660 (.ZN (n_434), .A (slo__sro_n375), .B1 (n_403), .B2 (n_402));
XNOR2_X2 slo__mro_c667 (.ZN (Res_out[36]), .A (slo__mro_n380), .B (n_265));
INV_X1 slo__mro_c705 (.ZN (slo__mro_n416), .A (sgo__sro_n301));
INV_X1 slo__mro_c706 (.ZN (slo__mro_n415), .A (n_193));
AND2_X2 slo__mro_c707 (.ZN (slo__mro_n414), .A1 (n_262), .A2 (slo__mro_n415));
OAI21_X4 slo__mro_c708 (.ZN (Res_out[52]), .A (n_261), .B1 (slo__mro_n414), .B2 (slo__mro_n416));
NOR2_X2 sgo__c502 (.ZN (sgo__n290), .A1 (Res_in[30]), .A2 (carry_in[30]));
INV_X4 sgo__c504 (.ZN (n_175), .A (sgo__n290));
OR2_X4 slo__xsl_c798 (.ZN (n_267), .A1 (carry_in[38]), .A2 (Res_in[38]));
INV_X1 slo__xsl_c867 (.ZN (slo__xsl_n558), .A (n_370));
NOR3_X4 slo__xsl_c870 (.ZN (n_370), .A1 (CLOCK_slo__sro_n1317), .A2 (n_250), .A3 (n_239));
INV_X4 CLOCK_opt_ipo_c1336 (.ZN (CLOCK_opt_ipo_n1035), .A (sgo__sro_n176));
OAI21_X2 CLOCK_slo__sro_c1831 (.ZN (CLOCK_slo__sro_n1363), .A (CLOCK_slo__sro_n1364)
    , .B1 (n_142), .B2 (n_295));
OR2_X2 CLOCK_slo__xsl_c2019 (.ZN (n_191), .A1 (carry_in[32]), .A2 (Res_in[32]));
INV_X1 opt_ipo_c1292 (.ZN (opt_ipo_n987), .A (n_48));
NAND2_X1 CLOCK_slo__sro_c1860 (.ZN (CLOCK_slo__sro_n1387), .A1 (CLOCK_slo__sro_n1388), .A2 (CLOCK_slo__sro_n1389));
NOR2_X1 CLOCK_slo__sro_c1861 (.ZN (n_392), .A1 (CLOCK_slo__sro_n1387), .A2 (n_343));
NAND2_X2 CLOCK_slo__mro_c1949 (.ZN (CLOCK_slo__mro_n1454), .A1 (n_132), .A2 (n_130));
INV_X2 CLOCK_slo__mro_c1936 (.ZN (CLOCK_slo__mro_n1442), .A (n_182));
NAND2_X4 CLOCK_slo__mro_c1952 (.ZN (Res_out[44]), .A1 (n_126), .A2 (n_128));
INV_X1 opt_ipo_c1311 (.ZN (opt_ipo_n1006), .A (opt_ipo_n1007));
INV_X1 opt_ipo_c1312 (.ZN (opt_ipo_n1007), .A (n_274));
INV_X2 CLOCK_slo__mro_c1947 (.ZN (CLOCK_slo__mro_n1456), .A (n_329));
INV_X4 opt_ipo_c1084 (.ZN (opt_ipo_n737), .A (n_252));
BUF_X1 CLOCK_opt_ipo_c1367 (.Z (CLOCK_opt_ipo_n1068), .A (n_276));
XNOR2_X2 CLOCK_slo__mro_c1937 (.ZN (Res_out[31]), .A (n_188), .B (CLOCK_slo__mro_n1442));

endmodule //datapath

module addResWithCarry (Res_out, Res_in, carry_in);

output [63:0] Res_out;
input [63:0] Res_in;
input [63:0] carry_in;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire uc_28;
wire uc_29;


datapath i_0 (.Res_out ({Res_out[63], Res_out[62], Res_out[61], Res_out[60], Res_out[59], 
    Res_out[58], Res_out[57], Res_out[56], Res_out[55], Res_out[54], Res_out[53], 
    Res_out[52], Res_out[51], Res_out[50], Res_out[49], Res_out[48], Res_out[47], 
    Res_out[46], Res_out[45], Res_out[44], Res_out[43], Res_out[42], Res_out[41], 
    Res_out[40], Res_out[39], Res_out[38], Res_out[37], Res_out[36], Res_out[35], 
    Res_out[34], Res_out[33], Res_out[32], Res_out[31], Res_out[30], Res_out[29], 
    Res_out[28], Res_out[27], Res_out[26], Res_out[25], Res_out[24], Res_out[23], 
    Res_out[22], Res_out[21], Res_out[20], Res_out[19], Res_out[18], Res_out[17], 
    Res_out[16], Res_out[15], Res_out[14], Res_out[13], Res_out[12], Res_out[11], 
    Res_out[10], Res_out[9], uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, 
    uc_29}), .Res_in ({uc_10, uc_11, Res_in[61], Res_in[60], Res_in[59], Res_in[58], 
    Res_in[57], Res_in[56], Res_in[55], Res_in[54], Res_in[53], Res_in[52], Res_in[51], 
    Res_in[50], Res_in[49], Res_in[48], Res_in[47], Res_in[46], Res_in[45], Res_in[44], 
    Res_in[43], Res_in[42], Res_in[41], Res_in[40], Res_in[39], Res_in[38], Res_in[37], 
    Res_in[36], Res_in[35], Res_in[34], Res_in[33], Res_in[32], Res_in[31], Res_in[30], 
    Res_in[29], Res_in[28], Res_in[27], Res_in[26], Res_in[25], Res_in[24], Res_in[23], 
    Res_in[22], Res_in[21], Res_in[20], Res_in[19], Res_in[18], Res_in[17], Res_in[16], 
    Res_in[15], Res_in[14], Res_in[13], Res_in[12], Res_in[11], Res_in[10], Res_in[9], 
    uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, uc_20}), .carry_in ({
    uc_0, carry_in[62], carry_in[61], carry_in[60], carry_in[59], carry_in[58], carry_in[57], 
    carry_in[56], carry_in[55], carry_in[54], carry_in[53], carry_in[52], carry_in[51], 
    carry_in[50], carry_in[49], carry_in[48], carry_in[47], carry_in[46], carry_in[45], 
    carry_in[44], carry_in[43], carry_in[42], carry_in[41], carry_in[40], carry_in[39], 
    carry_in[38], carry_in[37], carry_in[36], carry_in[35], carry_in[34], carry_in[33], 
    carry_in[32], carry_in[31], carry_in[30], carry_in[29], carry_in[28], carry_in[27], 
    carry_in[26], carry_in[25], carry_in[24], carry_in[23], carry_in[22], carry_in[21], 
    carry_in[20], carry_in[19], carry_in[18], carry_in[17], carry_in[16], carry_in[15], 
    carry_in[14], carry_in[13], carry_in[12], carry_in[11], carry_in[10], carry_in[9], 
    uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, uc_9}));

endmodule //addResWithCarry

module multiplyAllBits (B_7_PP_0, B_24_PP_0, B_4_PP_0, normalizedWires, A, B);

output [2047:0] normalizedWires;
input [31:0] A;
input [31:0] B;
input B_7_PP_0;
input B_24_PP_0;
input B_4_PP_0;
wire slo__n1036;
wire CLOCK_slo__n2403;
wire CLOCK_slo__n3235;
wire slo___n867;
wire opt_ipo_n1525;
wire opt_ipo_n1677;
wire slo___n1215;
wire CLOCK_slo__n2927;
wire slo__n298;
wire spw__n3533;
wire CLOCK_slo__n2250;
wire CLOCK_slo___n2514;
wire slo__n1191;
wire CLOCK_sgo__n1891;
wire CLOCK_slo___n3081;
wire slo_n1330;
wire slo_n705;
wire CLOCK_slo_n2535;
wire n_0_20;
wire CLOCK_slo__n3242;
wire n_0_25;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_36;
wire n_0_39;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_48;
wire n_0_51;
wire n_0_54;
wire n_0_57;
wire n_0_58;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_56;
wire n_0_5;
wire n_0_3;
wire n_0_2;
wire n_0_73;
wire sgo__n27;
wire opt_ipo_n1649;
wire sgo__n32;
wire n_0_15;
wire n_0_68;
wire n_0_67;
wire n_0_11;
wire n_0_19;
wire n_0_14;
wire n_0_13;
wire n_0_12;
wire n_0_10;
wire sgo__n175;
wire n_0_65;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_74;
wire opt_ipo_n1532;
wire sgo__n110;
wire n_0_76;
wire n_0_55;
wire n_0_53;
wire n_0_52;
wire n_0_50;
wire n_0_49;
wire n_0_47;
wire n_0_46;
wire n_0_40;
wire n_0_38;
wire n_0_35;
wire n_0_34;
wire sgo__n131;
wire n_0_33;
wire n_0_16;
wire n_0_32;
wire n_0_28;
wire n_0_27;
wire n_0_26;
wire n_0_23;
wire n_0_22;
wire n_0_21;
wire n_0_18;
wire n_0_17;
wire n_0_9;
wire CLOCK_slo___n2515;
wire n_0_4;
wire n_0_0;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_81;
wire n_0_82;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire sgo__n168;
wire n_0_106;
wire opt_ipo_n1647;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire opt_ipo_n1658;
wire sgo__n85;
wire CLOCK_slo__n2299;
wire slo__n302;
wire slo__n332;
wire slo__n317;
wire slo__n381;
wire slo___n436;
wire slo__n791;
wire CLOCK_slo__n3319;
wire slo__n616;
wire slo__n494;
wire slo__n785;
wire slo__n907;
wire slo__n1004;
wire CLOCK_slo__n2695;
wire slo__n1013;
wire slo__n1127;
wire slo__n1158;
wire CLOCK_sgo__n1896;
wire slo__n1306;
wire slo__n1353;
wire CLOCK_slo__n2241;
wire opt_ipo_n1648;
wire opt_ipo_n1675;
wire opt_ipo_n1550;
wire opt_ipo_n1556;
wire spw__n3534;
wire spw__n3569;
wire spw__n3498;
wire CLOCK_slo__n2545;
wire spw__n3570;
wire spw__n3571;
wire CLOCK_slo___n3082;
wire opt_ipo_n1710;
wire spw__n3572;
wire spw__n3573;
wire CLOCK_slo__n3096;
wire spw__n3574;
wire spw__n3575;


AND2_X4 i_0_534 (.ZN (normalizedWires[22]), .A1 (A[22]), .A2 (B[0]));
BUF_X8 opt_ipo_c1514 (.Z (opt_ipo_n1658), .A (n_0_20));
AND2_X1 i_0_1122 (.ZN (normalizedWires[1647]), .A1 (A[22]), .A2 (B[25]));
INV_X1 opt_ipo_c1503 (.ZN (opt_ipo_n1647), .A (opt_ipo_n1648));
AND2_X2 i_0_1120 (.ZN (normalizedWires[1582]), .A1 (A[22]), .A2 (slo_n1330));
INV_X1 slo__c1091 (.ZN (slo__n1191), .A (A[9]));
AND2_X4 i_0_1118 (.ZN (normalizedWires[79]), .A1 (A[14]), .A2 (B[1]));
AND2_X1 i_0_1117 (.ZN (normalizedWires[73]), .A1 (A[8]), .A2 (B[1]));
AND2_X1 i_0_1116 (.ZN (normalizedWires[71]), .A1 (A[6]), .A2 (B[1]));
AND2_X2 i_0_1115 (.ZN (normalizedWires[15]), .A1 (A[15]), .A2 (B[0]));
AND2_X1 i_0_1114 (.ZN (normalizedWires[13]), .A1 (A[13]), .A2 (B[0]));
AND2_X1 i_0_1113 (.ZN (normalizedWires[12]), .A1 (A[12]), .A2 (B[0]));
AND2_X1 i_0_1112 (.ZN (normalizedWires[11]), .A1 (A[11]), .A2 (B[0]));
AND2_X1 i_0_1111 (.ZN (normalizedWires[10]), .A1 (A[10]), .A2 (B[0]));
AND2_X1 i_0_1110 (.ZN (normalizedWires[6]), .A1 (A[6]), .A2 (B[0]));
NAND2_X1 i_0_1109 (.ZN (n_0_129), .A1 (sgo__n32), .A2 (B[25]));
INV_X1 i_0_1108 (.ZN (normalizedWires[1646]), .A (n_0_129));
NAND2_X1 i_0_1107 (.ZN (n_0_128), .A1 (sgo__n32), .A2 (slo_n1330));
INV_X1 i_0_1106 (.ZN (normalizedWires[1581]), .A (n_0_128));
NAND2_X1 i_0_1105 (.ZN (n_0_127), .A1 (A[25]), .A2 (B[22]));
INV_X1 i_0_1104 (.ZN (normalizedWires[1455]), .A (n_0_127));
NAND2_X1 i_0_1103 (.ZN (n_0_126), .A1 (A[22]), .A2 (B[22]));
INV_X1 i_0_1102 (.ZN (normalizedWires[1452]), .A (n_0_126));
NAND2_X1 i_0_1101 (.ZN (n_0_125), .A1 (sgo__n32), .A2 (B[22]));
INV_X1 i_0_1100 (.ZN (normalizedWires[1451]), .A (n_0_125));
NAND2_X1 i_0_1099 (.ZN (n_0_124), .A1 (A[26]), .A2 (B[21]));
INV_X1 i_0_1098 (.ZN (normalizedWires[1391]), .A (n_0_124));
NAND2_X1 i_0_1097 (.ZN (n_0_123), .A1 (A[22]), .A2 (B[21]));
INV_X1 i_0_1096 (.ZN (normalizedWires[1387]), .A (n_0_123));
NAND2_X1 i_0_1095 (.ZN (n_0_122), .A1 (sgo__n32), .A2 (B[21]));
INV_X1 i_0_1094 (.ZN (normalizedWires[1386]), .A (n_0_122));
NAND2_X1 i_0_1093 (.ZN (n_0_121), .A1 (A[26]), .A2 (B[19]));
INV_X1 i_0_1092 (.ZN (normalizedWires[1261]), .A (n_0_121));
NAND2_X1 i_0_1091 (.ZN (n_0_120), .A1 (A[25]), .A2 (slo__n494));
INV_X1 i_0_1090 (.ZN (normalizedWires[1260]), .A (n_0_120));
NAND2_X1 i_0_1089 (.ZN (n_0_119), .A1 (A[22]), .A2 (B[19]));
INV_X1 i_0_1088 (.ZN (normalizedWires[1257]), .A (n_0_119));
NAND2_X1 i_0_1087 (.ZN (n_0_118), .A1 (sgo__n32), .A2 (slo__n494));
INV_X1 i_0_1086 (.ZN (normalizedWires[1256]), .A (n_0_118));
NAND2_X1 i_0_1085 (.ZN (n_0_117), .A1 (A[26]), .A2 (B[18]));
INV_X1 i_0_1084 (.ZN (normalizedWires[1196]), .A (n_0_117));
NAND2_X1 i_0_1083 (.ZN (n_0_116), .A1 (A[25]), .A2 (B[18]));
INV_X1 i_0_1082 (.ZN (normalizedWires[1195]), .A (n_0_116));
NAND2_X1 i_0_1081 (.ZN (n_0_115), .A1 (A[22]), .A2 (B[18]));
INV_X1 i_0_1080 (.ZN (normalizedWires[1192]), .A (n_0_115));
NAND2_X2 i_0_1079 (.ZN (n_0_114), .A1 (A[27]), .A2 (B[16]));
INV_X2 i_0_1078 (.ZN (normalizedWires[1067]), .A (n_0_114));
NAND2_X1 i_0_1077 (.ZN (n_0_113), .A1 (A[26]), .A2 (B[16]));
INV_X2 i_0_1076 (.ZN (normalizedWires[1066]), .A (n_0_113));
NAND2_X1 i_0_1075 (.ZN (n_0_112), .A1 (A[25]), .A2 (B[16]));
INV_X1 i_0_1074 (.ZN (normalizedWires[1065]), .A (n_0_112));
NAND2_X1 i_0_1073 (.ZN (n_0_111), .A1 (A[22]), .A2 (B[16]));
INV_X2 i_0_1072 (.ZN (normalizedWires[1062]), .A (n_0_111));
NAND2_X2 i_0_1071 (.ZN (n_0_110), .A1 (A[27]), .A2 (B[15]));
INV_X2 i_0_1070 (.ZN (normalizedWires[1002]), .A (n_0_110));
NAND2_X1 i_0_1069 (.ZN (n_0_109), .A1 (A[26]), .A2 (B[15]));
INV_X2 i_0_1068 (.ZN (normalizedWires[1001]), .A (n_0_109));
NAND2_X1 i_0_1067 (.ZN (n_0_108), .A1 (A[22]), .A2 (B[15]));
INV_X1 i_0_1066 (.ZN (normalizedWires[997]), .A (n_0_108));
BUF_X4 sgo__c206 (.Z (sgo__n168), .A (n_0_27));
NAND2_X1 i_0_1064 (.ZN (n_0_106), .A1 (opt_ipo_n1648), .A2 (A[2]));
INV_X1 i_0_1063 (.ZN (normalizedWires[652]), .A (n_0_106));
INV_X8 opt_ipo_c1392 (.ZN (opt_ipo_n1532), .A (A[23]));
NAND2_X1 i_0_1061 (.ZN (n_0_104), .A1 (B[9]), .A2 (A[4]));
INV_X1 i_0_1060 (.ZN (normalizedWires[589]), .A (n_0_104));
NAND2_X1 i_0_1059 (.ZN (n_0_103), .A1 (B[9]), .A2 (A[3]));
INV_X1 i_0_1058 (.ZN (normalizedWires[588]), .A (n_0_103));
NAND2_X1 i_0_1057 (.ZN (n_0_102), .A1 (slo_n705), .A2 (A[3]));
INV_X2 i_0_1055 (.ZN (normalizedWires[458]), .A (n_0_102));
NAND2_X1 i_0_962 (.ZN (n_0_101), .A1 (B[6]), .A2 (A[5]));
INV_X1 i_0_961 (.ZN (normalizedWires[395]), .A (n_0_101));
NAND2_X1 i_0_960 (.ZN (n_0_100), .A1 (B[6]), .A2 (A[4]));
INV_X1 i_0_959 (.ZN (normalizedWires[394]), .A (n_0_100));
NAND2_X1 i_0_932 (.ZN (n_0_99), .A1 (B[6]), .A2 (A[3]));
INV_X1 i_0_931 (.ZN (normalizedWires[393]), .A (n_0_99));
NAND2_X1 i_0_930 (.ZN (n_0_98), .A1 (CLOCK_slo_n2535), .A2 (A[7]));
INV_X1 i_0_929 (.ZN (normalizedWires[267]), .A (n_0_98));
NAND2_X1 i_0_854 (.ZN (n_0_97), .A1 (sgo__n32), .A2 (B[3]));
INV_X1 i_0_853 (.ZN (normalizedWires[216]), .A (n_0_97));
NAND2_X1 i_0_822 (.ZN (n_0_96), .A1 (A[7]), .A2 (B[3]));
INV_X1 i_0_821 (.ZN (normalizedWires[202]), .A (n_0_96));
NAND2_X1 i_0_799 (.ZN (n_0_95), .A1 (A[8]), .A2 (B[2]));
INV_X1 i_0_761 (.ZN (normalizedWires[138]), .A (n_0_95));
NAND2_X1 i_0_758 (.ZN (n_0_94), .A1 (A[7]), .A2 (B[2]));
INV_X1 i_0_757 (.ZN (normalizedWires[137]), .A (n_0_94));
NAND2_X1 i_0_735 (.ZN (n_0_93), .A1 (A[21]), .A2 (B[1]));
INV_X1 i_0_730 (.ZN (normalizedWires[86]), .A (n_0_93));
NAND2_X1 i_0_726 (.ZN (n_0_92), .A1 (A[17]), .A2 (B[1]));
INV_X1 i_0_725 (.ZN (normalizedWires[82]), .A (n_0_92));
NAND2_X4 i_0_703 (.ZN (n_0_91), .A1 (A[15]), .A2 (B[1]));
INV_X4 i_0_666 (.ZN (normalizedWires[80]), .A (n_0_91));
NAND2_X2 i_0_665 (.ZN (n_0_90), .A1 (A[13]), .A2 (B[1]));
INV_X4 i_0_662 (.ZN (normalizedWires[78]), .A (n_0_90));
NAND2_X1 i_0_661 (.ZN (n_0_89), .A1 (A[12]), .A2 (B[1]));
INV_X1 i_0_639 (.ZN (normalizedWires[77]), .A (n_0_89));
NAND2_X1 i_0_634 (.ZN (n_0_88), .A1 (A[11]), .A2 (B[1]));
INV_X1 i_0_633 (.ZN (normalizedWires[76]), .A (n_0_88));
NAND2_X1 i_0_630 (.ZN (n_0_87), .A1 (A[10]), .A2 (B[1]));
INV_X1 i_0_607 (.ZN (normalizedWires[75]), .A (n_0_87));
NAND2_X1 i_0_571 (.ZN (n_0_86), .A1 (A[9]), .A2 (B[1]));
INV_X1 i_0_570 (.ZN (normalizedWires[74]), .A (n_0_86));
NAND2_X1 i_0_569 (.ZN (n_0_85), .A1 (A[7]), .A2 (B[1]));
INV_X2 i_0_566 (.ZN (normalizedWires[72]), .A (n_0_85));
NAND2_X1 i_0_543 (.ZN (n_0_84), .A1 (A[5]), .A2 (B[1]));
INV_X1 i_0_539 (.ZN (normalizedWires[70]), .A (n_0_84));
NAND2_X1 i_0_511 (.ZN (n_0_82), .A1 (A[20]), .A2 (B[0]));
INV_X1 i_0_355 (.ZN (normalizedWires[20]), .A (n_0_82));
NAND2_X4 i_0_354 (.ZN (n_0_81), .A1 (A[16]), .A2 (B[0]));
INV_X4 i_0_353 (.ZN (normalizedWires[16]), .A (n_0_81));
NAND2_X2 i_0_351 (.ZN (normalizedWires[14]), .A1 (A[14]), .A2 (B[0]));
CLKBUF_X3 CLOCK_sgo__c1758 (.Z (CLOCK_sgo__n1891), .A (n_0_15));
NAND2_X1 i_0_323 (.ZN (n_0_79), .A1 (A[9]), .A2 (B[0]));
INV_X1 i_0_319 (.ZN (normalizedWires[9]), .A (n_0_79));
NAND2_X1 i_0_259 (.ZN (n_0_78), .A1 (A[8]), .A2 (B[0]));
INV_X1 i_0_255 (.ZN (normalizedWires[8]), .A (n_0_78));
NAND2_X1 i_0_229 (.ZN (n_0_77), .A1 (A[7]), .A2 (B[0]));
INV_X1 i_0_228 (.ZN (normalizedWires[7]), .A (n_0_77));
INV_X2 i_0_227 (.ZN (n_0_0), .A (B[0]));
INV_X4 i_0_223 (.ZN (n_0_4), .A (A[3]));
NOR2_X4 CLOCK_slo__sro_c2694 (.ZN (normalizedWires[673]), .A1 (opt_ipo_n1532), .A2 (opt_ipo_n1649));
INV_X4 i_0_166 (.ZN (n_0_9), .A (A[8]));
INV_X4 i_0_159 (.ZN (n_0_17), .A (A[16]));
INV_X1 i_0_149 (.ZN (n_0_18), .A (A[17]));
INV_X16 i_0_135 (.ZN (n_0_21), .A (A[20]));
INV_X8 i_0_134 (.ZN (n_0_22), .A (A[21]));
INV_X8 i_0_127 (.ZN (n_0_23), .A (A[22]));
INV_X8 i_0_104 (.ZN (n_0_26), .A (A[25]));
INV_X8 i_0_103 (.ZN (n_0_27), .A (A[26]));
INV_X8 i_0_95 (.ZN (n_0_28), .A (A[27]));
INV_X8 i_0_86 (.ZN (n_0_32), .A (B[1]));
INV_X4 i_0_85 (.ZN (n_0_16), .A (A[15]));
INV_X4 i_0_81 (.ZN (n_0_33), .A (B[2]));
BUF_X4 sgo__c138 (.Z (sgo__n110), .A (n_0_23));
INV_X4 i_0_76 (.ZN (n_0_34), .A (B[3]));
INV_X4 i_0_75 (.ZN (n_0_35), .A (B[4]));
INV_X4 i_0_74 (.ZN (spw__n3498), .A (B[6]));
INV_X16 i_0_72 (.ZN (n_0_38), .A (B[7]));
INV_X8 i_0_71 (.ZN (n_0_40), .A (B[9]));
INV_X8 i_0_70 (.ZN (n_0_46), .A (B[15]));
INV_X8 i_0_69 (.ZN (n_0_47), .A (B[16]));
INV_X8 i_0_55 (.ZN (n_0_49), .A (B[18]));
INV_X8 i_0_53 (.ZN (n_0_50), .A (B[19]));
INV_X4 i_0_51 (.ZN (n_0_52), .A (B[21]));
INV_X16 i_0_46 (.ZN (n_0_53), .A (B[22]));
INV_X4 i_0_45 (.ZN (n_0_55), .A (B[24]));
INV_X8 i_0_43 (.ZN (n_0_76), .A (A[7]));
CLKBUF_X3 sgo__c112 (.Z (sgo__n85), .A (n_0_50));
INV_X1 CLOCK_slo__c2137 (.ZN (CLOCK_slo__n2299), .A (B[16]));
NAND2_X1 i_0_38 (.ZN (n_0_74), .A1 (B[10]), .A2 (A[3]));
INV_X1 i_0_37 (.ZN (normalizedWires[653]), .A (n_0_74));
NOR2_X1 slo__mro_c283 (.ZN (normalizedWires[1369]), .A1 (n_0_52), .A2 (opt_ipo_n1710));
NAND2_X1 i_0_34 (.ZN (n_0_71), .A1 (opt_ipo_n1648), .A2 (A[1]));
INV_X1 i_0_33 (.ZN (normalizedWires[651]), .A (n_0_71));
NAND2_X1 i_0_32 (.ZN (n_0_70), .A1 (A[6]), .A2 (CLOCK_slo___n2514));
INV_X1 i_0_31 (.ZN (normalizedWires[266]), .A (n_0_70));
NAND2_X1 i_0_28 (.ZN (n_0_69), .A1 (A[6]), .A2 (B[3]));
INV_X1 i_0_26 (.ZN (normalizedWires[201]), .A (n_0_69));
NAND2_X1 i_0_25 (.ZN (n_0_65), .A1 (A[18]), .A2 (B[0]));
INV_X1 i_0_24 (.ZN (normalizedWires[18]), .A (n_0_65));
BUF_X4 sgo__c168 (.Z (sgo__n131), .A (n_0_29));
INV_X4 i_0_20 (.ZN (n_0_10), .A (A[9]));
INV_X8 i_0_18 (.ZN (n_0_12), .A (A[11]));
INV_X4 i_0_17 (.ZN (n_0_13), .A (A[12]));
INV_X8 i_0_16 (.ZN (n_0_14), .A (A[13]));
INV_X16 i_0_14 (.ZN (n_0_19), .A (A[18]));
INV_X4 i_0_13 (.ZN (n_0_11), .A (A[10]));
NOR2_X2 CLOCK_slo__mro_c1872 (.ZN (normalizedWires[1777]), .A1 (sgo__n110), .A2 (n_0_58));
INV_X8 i_0_7 (.ZN (n_0_67), .A (A[6]));
INV_X8 i_0_5 (.ZN (n_0_68), .A (A[5]));
INV_X8 i_0_1056 (.ZN (n_0_15), .A (A[14]));
BUF_X4 sgo__c38 (.Z (sgo__n32), .A (A[21]));
BUF_X4 sgo__c33 (.Z (sgo__n27), .A (n_0_26));
INV_X8 opt_ipo_c1505 (.ZN (opt_ipo_n1649), .A (B[10]));
NOR2_X1 i_0_838 (.ZN (normalizedWires[1888]), .A1 (n_0_63), .A2 (CLOCK_slo___n3082));
NOR2_X1 i_0_837 (.ZN (normalizedWires[1887]), .A1 (n_0_63), .A2 (n_0_3));
NOR2_X1 i_0_836 (.ZN (normalizedWires[1886]), .A1 (n_0_63), .A2 (n_0_2));
NOR2_X1 i_0_835 (.ZN (normalizedWires[1885]), .A1 (n_0_63), .A2 (n_0_73));
NOR2_X1 i_0_834 (.ZN (normalizedWires[1824]), .A1 (n_0_64), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_833 (.ZN (normalizedWires[1823]), .A1 (n_0_64), .A2 (CLOCK_slo___n3082));
NOR2_X1 i_0_831 (.ZN (normalizedWires[1822]), .A1 (n_0_64), .A2 (n_0_3));
NOR2_X1 i_0_78 (.ZN (normalizedWires[1821]), .A1 (n_0_64), .A2 (n_0_2));
NOR2_X2 i_0_77 (.ZN (normalizedWires[1632]), .A1 (n_0_56), .A2 (n_0_76));
NOR2_X2 i_0_73 (.ZN (normalizedWires[1631]), .A1 (n_0_56), .A2 (n_0_67));
NOR2_X2 i_0_63 (.ZN (normalizedWires[1630]), .A1 (n_0_56), .A2 (sgo__n175));
NOR2_X1 i_0_30 (.ZN (normalizedWires[1629]), .A1 (n_0_56), .A2 (opt_ipo_n1710));
NOR2_X2 CLOCK_slo__sro_c2674 (.ZN (normalizedWires[282]), .A1 (n_0_23), .A2 (n_0_35));
NOR2_X1 i_0_27 (.ZN (normalizedWires[1627]), .A1 (n_0_56), .A2 (n_0_3));
NOR2_X1 i_0_22 (.ZN (normalizedWires[1626]), .A1 (n_0_56), .A2 (n_0_2));
INV_X2 i_0_21 (.ZN (n_0_73), .A (A[0]));
INV_X4 i_0_19 (.ZN (n_0_2), .A (A[1]));
INV_X4 i_0_15 (.ZN (n_0_3), .A (A[2]));
INV_X8 i_0_11 (.ZN (n_0_5), .A (A[4]));
INV_X8 i_0_3 (.ZN (n_0_56), .A (B[25]));
INV_X16 i_0_1 (.ZN (n_0_64), .A (B[28]));
INV_X2 i_0_0 (.ZN (n_0_63), .A (B[29]));
NOR2_X1 i_0_1054 (.ZN (normalizedWires[2045]), .A1 (slo__n785), .A2 (n_0_62));
NOR2_X1 i_0_1053 (.ZN (normalizedWires[2044]), .A1 (slo__n332), .A2 (n_0_62));
NOR2_X1 i_0_1052 (.ZN (normalizedWires[2043]), .A1 (sgo__n131), .A2 (n_0_62));
NOR2_X1 i_0_1051 (.ZN (normalizedWires[2042]), .A1 (spw__n3534), .A2 (n_0_62));
NOR2_X1 i_0_1050 (.ZN (normalizedWires[2041]), .A1 (sgo__n168), .A2 (n_0_62));
NOR2_X1 i_0_1049 (.ZN (normalizedWires[2040]), .A1 (sgo__n27), .A2 (n_0_62));
NOR2_X1 i_0_1048 (.ZN (normalizedWires[2039]), .A1 (opt_ipo_n1677), .A2 (n_0_62));
NOR2_X1 i_0_1047 (.ZN (normalizedWires[2038]), .A1 (slo___n1215), .A2 (n_0_62));
NOR2_X1 i_0_1046 (.ZN (normalizedWires[2037]), .A1 (sgo__n110), .A2 (n_0_62));
NOR2_X1 i_0_1045 (.ZN (normalizedWires[2036]), .A1 (slo__n302), .A2 (n_0_62));
NOR2_X1 i_0_1044 (.ZN (normalizedWires[2035]), .A1 (n_0_21), .A2 (n_0_62));
NOR2_X1 i_0_1043 (.ZN (normalizedWires[2034]), .A1 (opt_ipo_n1658), .A2 (n_0_62));
NOR2_X1 i_0_1042 (.ZN (normalizedWires[2033]), .A1 (n_0_19), .A2 (n_0_62));
NOR2_X1 i_0_1041 (.ZN (normalizedWires[2032]), .A1 (slo__n298), .A2 (n_0_62));
NOR2_X1 i_0_1040 (.ZN (normalizedWires[2031]), .A1 (opt_ipo_n1550), .A2 (n_0_62));
NOR2_X1 i_0_1039 (.ZN (normalizedWires[2030]), .A1 (n_0_16), .A2 (n_0_62));
NOR2_X1 i_0_1038 (.ZN (normalizedWires[2029]), .A1 (CLOCK_sgo__n1891), .A2 (n_0_62));
NOR2_X1 i_0_1037 (.ZN (normalizedWires[2028]), .A1 (n_0_14), .A2 (n_0_62));
NOR2_X1 i_0_1036 (.ZN (normalizedWires[2027]), .A1 (CLOCK_sgo__n1896), .A2 (n_0_62));
NOR2_X1 i_0_1035 (.ZN (normalizedWires[2026]), .A1 (opt_ipo_n1525), .A2 (n_0_62));
NOR2_X1 i_0_1034 (.ZN (normalizedWires[2025]), .A1 (n_0_11), .A2 (n_0_62));
NOR2_X1 i_0_1033 (.ZN (normalizedWires[2024]), .A1 (opt_ipo_n1556), .A2 (n_0_62));
NOR2_X1 i_0_1032 (.ZN (normalizedWires[2023]), .A1 (n_0_9), .A2 (n_0_62));
NOR2_X1 i_0_1031 (.ZN (normalizedWires[2022]), .A1 (slo__n1013), .A2 (n_0_62));
NOR2_X1 i_0_1030 (.ZN (normalizedWires[2021]), .A1 (n_0_67), .A2 (n_0_62));
NOR2_X1 i_0_1029 (.ZN (normalizedWires[2020]), .A1 (sgo__n175), .A2 (n_0_62));
NOR2_X1 i_0_1028 (.ZN (normalizedWires[2019]), .A1 (opt_ipo_n1710), .A2 (n_0_62));
NOR2_X1 i_0_1027 (.ZN (normalizedWires[2018]), .A1 (CLOCK_slo___n3082), .A2 (n_0_62));
NOR2_X1 i_0_1026 (.ZN (normalizedWires[2017]), .A1 (n_0_3), .A2 (n_0_62));
NOR2_X1 i_0_1025 (.ZN (normalizedWires[2016]), .A1 (n_0_2), .A2 (n_0_62));
NOR2_X1 i_0_1024 (.ZN (normalizedWires[2015]), .A1 (n_0_73), .A2 (n_0_62));
INV_X2 i_0_1023 (.ZN (n_0_62), .A (B[31]));
NOR2_X1 i_0_1022 (.ZN (normalizedWires[1980]), .A1 (n_0_61), .A2 (slo__n785));
NOR2_X1 i_0_1021 (.ZN (normalizedWires[1979]), .A1 (n_0_61), .A2 (slo__n332));
NOR2_X1 i_0_1020 (.ZN (normalizedWires[1978]), .A1 (n_0_61), .A2 (sgo__n131));
NOR2_X1 i_0_1019 (.ZN (normalizedWires[1977]), .A1 (n_0_61), .A2 (spw__n3534));
NOR2_X1 i_0_1018 (.ZN (normalizedWires[1976]), .A1 (n_0_61), .A2 (sgo__n168));
NOR2_X1 i_0_1017 (.ZN (normalizedWires[1975]), .A1 (n_0_61), .A2 (sgo__n27));
NOR2_X1 i_0_1016 (.ZN (normalizedWires[1974]), .A1 (n_0_61), .A2 (opt_ipo_n1677));
NOR2_X1 i_0_1015 (.ZN (normalizedWires[1973]), .A1 (n_0_61), .A2 (slo___n1215));
NOR2_X1 i_0_1014 (.ZN (normalizedWires[1972]), .A1 (n_0_61), .A2 (sgo__n110));
NOR2_X1 i_0_1013 (.ZN (normalizedWires[1971]), .A1 (n_0_61), .A2 (slo__n302));
NOR2_X1 i_0_1012 (.ZN (normalizedWires[1970]), .A1 (n_0_61), .A2 (n_0_21));
NOR2_X1 i_0_1011 (.ZN (normalizedWires[1969]), .A1 (n_0_61), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_1010 (.ZN (normalizedWires[1968]), .A1 (n_0_61), .A2 (n_0_19));
NOR2_X1 i_0_1009 (.ZN (normalizedWires[1967]), .A1 (n_0_61), .A2 (slo__n298));
NOR2_X1 i_0_1008 (.ZN (normalizedWires[1966]), .A1 (n_0_61), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_1007 (.ZN (normalizedWires[1965]), .A1 (n_0_61), .A2 (n_0_16));
NOR2_X1 i_0_1006 (.ZN (normalizedWires[1964]), .A1 (n_0_61), .A2 (CLOCK_sgo__n1891));
NOR2_X1 i_0_1005 (.ZN (normalizedWires[1963]), .A1 (n_0_61), .A2 (n_0_14));
NOR2_X1 i_0_1004 (.ZN (normalizedWires[1962]), .A1 (n_0_61), .A2 (CLOCK_sgo__n1896));
NOR2_X1 i_0_1003 (.ZN (normalizedWires[1961]), .A1 (n_0_61), .A2 (opt_ipo_n1525));
NOR2_X1 i_0_1002 (.ZN (normalizedWires[1960]), .A1 (n_0_61), .A2 (n_0_11));
NOR2_X1 i_0_1001 (.ZN (normalizedWires[1959]), .A1 (n_0_61), .A2 (opt_ipo_n1556));
NOR2_X1 i_0_1000 (.ZN (normalizedWires[1958]), .A1 (n_0_61), .A2 (n_0_9));
NOR2_X1 i_0_999 (.ZN (normalizedWires[1957]), .A1 (n_0_61), .A2 (slo__n1013));
NOR2_X1 i_0_998 (.ZN (normalizedWires[1956]), .A1 (n_0_61), .A2 (n_0_67));
NOR2_X1 i_0_997 (.ZN (normalizedWires[1955]), .A1 (n_0_61), .A2 (sgo__n175));
NOR2_X1 i_0_996 (.ZN (normalizedWires[1954]), .A1 (n_0_61), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_995 (.ZN (normalizedWires[1953]), .A1 (n_0_61), .A2 (CLOCK_slo___n3082));
NOR2_X1 i_0_994 (.ZN (normalizedWires[1952]), .A1 (n_0_61), .A2 (n_0_3));
NOR2_X1 i_0_993 (.ZN (normalizedWires[1951]), .A1 (n_0_61), .A2 (n_0_2));
NOR2_X1 i_0_992 (.ZN (normalizedWires[1950]), .A1 (n_0_61), .A2 (n_0_73));
INV_X2 i_0_991 (.ZN (n_0_61), .A (B[30]));
NOR2_X1 i_0_990 (.ZN (normalizedWires[1915]), .A1 (n_0_63), .A2 (slo__n785));
NOR2_X1 i_0_989 (.ZN (normalizedWires[1914]), .A1 (n_0_63), .A2 (slo__n332));
NOR2_X1 i_0_988 (.ZN (normalizedWires[1913]), .A1 (n_0_63), .A2 (sgo__n131));
NOR2_X1 i_0_987 (.ZN (normalizedWires[1912]), .A1 (n_0_63), .A2 (spw__n3534));
NOR2_X1 i_0_986 (.ZN (normalizedWires[1911]), .A1 (n_0_63), .A2 (sgo__n168));
NOR2_X1 i_0_985 (.ZN (normalizedWires[1910]), .A1 (n_0_63), .A2 (sgo__n27));
NOR2_X1 i_0_984 (.ZN (normalizedWires[1909]), .A1 (n_0_63), .A2 (opt_ipo_n1677));
NOR2_X1 i_0_983 (.ZN (normalizedWires[1908]), .A1 (n_0_63), .A2 (slo___n1215));
NOR2_X1 i_0_982 (.ZN (normalizedWires[1907]), .A1 (n_0_63), .A2 (sgo__n110));
NOR2_X1 i_0_981 (.ZN (normalizedWires[1906]), .A1 (n_0_63), .A2 (slo__n302));
NOR2_X1 i_0_980 (.ZN (normalizedWires[1905]), .A1 (n_0_63), .A2 (n_0_21));
NOR2_X1 i_0_979 (.ZN (normalizedWires[1904]), .A1 (n_0_63), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_978 (.ZN (normalizedWires[1903]), .A1 (n_0_63), .A2 (n_0_19));
NOR2_X1 i_0_977 (.ZN (normalizedWires[1902]), .A1 (n_0_63), .A2 (slo__n298));
NOR2_X1 i_0_976 (.ZN (normalizedWires[1901]), .A1 (n_0_63), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_975 (.ZN (normalizedWires[1900]), .A1 (n_0_63), .A2 (n_0_16));
NOR2_X1 i_0_974 (.ZN (normalizedWires[1899]), .A1 (n_0_63), .A2 (CLOCK_sgo__n1891));
NOR2_X1 i_0_973 (.ZN (normalizedWires[1898]), .A1 (n_0_63), .A2 (n_0_14));
NOR2_X1 i_0_972 (.ZN (normalizedWires[1897]), .A1 (n_0_63), .A2 (CLOCK_sgo__n1896));
NOR2_X1 i_0_971 (.ZN (normalizedWires[1896]), .A1 (n_0_63), .A2 (opt_ipo_n1525));
NOR2_X1 i_0_970 (.ZN (normalizedWires[1895]), .A1 (n_0_63), .A2 (n_0_11));
NOR2_X1 i_0_969 (.ZN (normalizedWires[1894]), .A1 (n_0_63), .A2 (opt_ipo_n1556));
NOR2_X1 i_0_968 (.ZN (normalizedWires[1893]), .A1 (n_0_63), .A2 (n_0_9));
NOR2_X1 i_0_967 (.ZN (normalizedWires[1892]), .A1 (n_0_63), .A2 (slo__n1013));
NOR2_X1 i_0_966 (.ZN (normalizedWires[1891]), .A1 (n_0_63), .A2 (n_0_67));
NOR2_X1 i_0_965 (.ZN (normalizedWires[1890]), .A1 (n_0_63), .A2 (sgo__n175));
NOR2_X1 i_0_964 (.ZN (normalizedWires[1889]), .A1 (n_0_63), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_958 (.ZN (normalizedWires[1850]), .A1 (n_0_64), .A2 (slo__n785));
NOR2_X1 i_0_957 (.ZN (normalizedWires[1849]), .A1 (n_0_64), .A2 (slo__n332));
NOR2_X1 i_0_956 (.ZN (normalizedWires[1848]), .A1 (n_0_64), .A2 (sgo__n131));
NOR2_X1 i_0_955 (.ZN (normalizedWires[1847]), .A1 (n_0_64), .A2 (spw__n3533));
NOR2_X1 i_0_954 (.ZN (normalizedWires[1846]), .A1 (n_0_64), .A2 (sgo__n168));
NOR2_X1 i_0_953 (.ZN (normalizedWires[1845]), .A1 (n_0_64), .A2 (sgo__n27));
NOR2_X1 i_0_952 (.ZN (normalizedWires[1844]), .A1 (n_0_64), .A2 (opt_ipo_n1677));
NOR2_X1 i_0_951 (.ZN (normalizedWires[1843]), .A1 (n_0_64), .A2 (slo___n1215));
NOR2_X1 i_0_950 (.ZN (normalizedWires[1842]), .A1 (sgo__n110), .A2 (n_0_64));
NOR2_X1 i_0_949 (.ZN (normalizedWires[1841]), .A1 (n_0_64), .A2 (slo__n302));
NOR2_X1 i_0_948 (.ZN (normalizedWires[1840]), .A1 (n_0_64), .A2 (n_0_21));
NOR2_X1 i_0_947 (.ZN (normalizedWires[1839]), .A1 (opt_ipo_n1658), .A2 (n_0_64));
NOR2_X1 i_0_946 (.ZN (normalizedWires[1838]), .A1 (n_0_64), .A2 (n_0_19));
NOR2_X1 i_0_945 (.ZN (normalizedWires[1837]), .A1 (n_0_64), .A2 (slo__n317));
NOR2_X1 i_0_944 (.ZN (normalizedWires[1836]), .A1 (n_0_64), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_943 (.ZN (normalizedWires[1835]), .A1 (n_0_64), .A2 (n_0_16));
NOR2_X2 slo__sro_c659 (.ZN (normalizedWires[1183]), .A1 (n_0_49), .A2 (n_0_14));
NOR2_X1 i_0_941 (.ZN (normalizedWires[1833]), .A1 (n_0_64), .A2 (n_0_14));
NOR2_X1 i_0_940 (.ZN (normalizedWires[1832]), .A1 (n_0_64), .A2 (n_0_13));
NOR2_X1 i_0_939 (.ZN (normalizedWires[1831]), .A1 (n_0_64), .A2 (opt_ipo_n1525));
NOR2_X1 i_0_938 (.ZN (normalizedWires[1830]), .A1 (n_0_64), .A2 (n_0_11));
NOR2_X1 i_0_937 (.ZN (normalizedWires[1829]), .A1 (n_0_64), .A2 (opt_ipo_n1556));
NOR2_X1 i_0_936 (.ZN (normalizedWires[1828]), .A1 (n_0_64), .A2 (n_0_9));
NOR2_X1 i_0_935 (.ZN (normalizedWires[1827]), .A1 (n_0_64), .A2 (slo__n1013));
NOR2_X1 i_0_934 (.ZN (normalizedWires[1826]), .A1 (n_0_64), .A2 (n_0_67));
NOR2_X1 i_0_933 (.ZN (normalizedWires[1825]), .A1 (n_0_64), .A2 (sgo__n175));
NOR2_X1 i_0_928 (.ZN (normalizedWires[1820]), .A1 (n_0_64), .A2 (n_0_73));
NOR2_X1 i_0_926 (.ZN (normalizedWires[1785]), .A1 (n_0_58), .A2 (slo__n785));
NOR2_X1 i_0_925 (.ZN (normalizedWires[1784]), .A1 (n_0_58), .A2 (slo__n332));
NOR2_X1 i_0_924 (.ZN (normalizedWires[1783]), .A1 (n_0_58), .A2 (sgo__n131));
NOR2_X1 i_0_923 (.ZN (normalizedWires[1782]), .A1 (n_0_58), .A2 (spw__n3533));
NOR2_X1 i_0_922 (.ZN (normalizedWires[1781]), .A1 (n_0_58), .A2 (sgo__n168));
NOR2_X1 i_0_921 (.ZN (normalizedWires[1780]), .A1 (n_0_58), .A2 (sgo__n27));
NOR2_X1 i_0_920 (.ZN (normalizedWires[1779]), .A1 (n_0_58), .A2 (opt_ipo_n1677));
NOR2_X1 i_0_919 (.ZN (normalizedWires[1778]), .A1 (n_0_58), .A2 (slo___n1215));
NOR2_X1 CLOCK_slo__mro_c1893 (.ZN (normalizedWires[209]), .A1 (n_0_15), .A2 (n_0_34));
NOR2_X1 i_0_917 (.ZN (normalizedWires[1776]), .A1 (n_0_58), .A2 (slo__n302));
NOR2_X1 i_0_916 (.ZN (normalizedWires[1775]), .A1 (n_0_58), .A2 (n_0_21));
NOR2_X1 i_0_915 (.ZN (normalizedWires[1774]), .A1 (n_0_58), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_914 (.ZN (normalizedWires[1773]), .A1 (n_0_58), .A2 (n_0_19));
NOR2_X1 i_0_913 (.ZN (normalizedWires[1772]), .A1 (slo__n298), .A2 (n_0_58));
NOR2_X1 i_0_912 (.ZN (normalizedWires[1771]), .A1 (n_0_58), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_911 (.ZN (normalizedWires[1770]), .A1 (n_0_58), .A2 (n_0_16));
NOR2_X1 i_0_910 (.ZN (normalizedWires[1769]), .A1 (n_0_58), .A2 (n_0_15));
NOR2_X1 i_0_909 (.ZN (normalizedWires[1768]), .A1 (n_0_58), .A2 (n_0_14));
NOR2_X1 i_0_908 (.ZN (normalizedWires[1767]), .A1 (n_0_58), .A2 (n_0_13));
NOR2_X1 i_0_907 (.ZN (normalizedWires[1766]), .A1 (n_0_58), .A2 (opt_ipo_n1525));
NOR2_X1 i_0_906 (.ZN (normalizedWires[1765]), .A1 (n_0_58), .A2 (n_0_11));
NOR2_X1 i_0_905 (.ZN (normalizedWires[1764]), .A1 (n_0_58), .A2 (opt_ipo_n1556));
NOR2_X1 i_0_904 (.ZN (normalizedWires[1763]), .A1 (n_0_58), .A2 (n_0_9));
NOR2_X1 i_0_903 (.ZN (normalizedWires[1762]), .A1 (n_0_58), .A2 (slo__n1013));
NOR2_X1 i_0_902 (.ZN (normalizedWires[1761]), .A1 (n_0_58), .A2 (n_0_67));
NOR2_X1 i_0_901 (.ZN (normalizedWires[1760]), .A1 (n_0_58), .A2 (sgo__n175));
NOR2_X1 i_0_900 (.ZN (normalizedWires[1759]), .A1 (n_0_58), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_899 (.ZN (normalizedWires[1758]), .A1 (n_0_58), .A2 (CLOCK_slo___n3082));
NOR2_X1 i_0_898 (.ZN (normalizedWires[1757]), .A1 (n_0_58), .A2 (n_0_3));
NOR2_X1 i_0_897 (.ZN (normalizedWires[1756]), .A1 (n_0_58), .A2 (n_0_2));
NOR2_X1 i_0_896 (.ZN (normalizedWires[1755]), .A1 (n_0_58), .A2 (n_0_73));
INV_X8 i_0_895 (.ZN (n_0_58), .A (B[27]));
NOR2_X1 i_0_894 (.ZN (normalizedWires[1720]), .A1 (n_0_57), .A2 (slo__n785));
NOR2_X1 i_0_893 (.ZN (normalizedWires[1719]), .A1 (n_0_57), .A2 (slo__n332));
NOR2_X1 i_0_892 (.ZN (normalizedWires[1718]), .A1 (n_0_57), .A2 (sgo__n131));
NOR2_X1 i_0_891 (.ZN (normalizedWires[1717]), .A1 (n_0_57), .A2 (spw__n3533));
NOR2_X1 i_0_890 (.ZN (normalizedWires[1716]), .A1 (n_0_57), .A2 (sgo__n168));
NOR2_X1 i_0_889 (.ZN (normalizedWires[1715]), .A1 (n_0_57), .A2 (sgo__n27));
NOR2_X1 i_0_888 (.ZN (normalizedWires[1714]), .A1 (n_0_57), .A2 (opt_ipo_n1677));
NOR2_X1 i_0_887 (.ZN (normalizedWires[1713]), .A1 (n_0_57), .A2 (slo___n1215));
NOR2_X1 i_0_886 (.ZN (normalizedWires[1712]), .A1 (n_0_57), .A2 (sgo__n110));
NOR2_X1 i_0_885 (.ZN (normalizedWires[1711]), .A1 (n_0_57), .A2 (slo__n302));
NOR2_X1 i_0_884 (.ZN (normalizedWires[1710]), .A1 (n_0_57), .A2 (n_0_21));
NOR2_X1 i_0_883 (.ZN (normalizedWires[1709]), .A1 (n_0_57), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_882 (.ZN (normalizedWires[1708]), .A1 (n_0_57), .A2 (n_0_19));
NOR2_X1 i_0_881 (.ZN (normalizedWires[1707]), .A1 (n_0_57), .A2 (slo__n298));
NOR2_X1 i_0_880 (.ZN (normalizedWires[1706]), .A1 (n_0_57), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_879 (.ZN (normalizedWires[1705]), .A1 (n_0_57), .A2 (n_0_16));
NOR2_X1 i_0_878 (.ZN (normalizedWires[1704]), .A1 (n_0_57), .A2 (n_0_15));
NOR2_X1 i_0_877 (.ZN (normalizedWires[1703]), .A1 (n_0_57), .A2 (n_0_14));
NOR2_X1 i_0_876 (.ZN (normalizedWires[1702]), .A1 (n_0_57), .A2 (n_0_13));
NOR2_X1 i_0_875 (.ZN (normalizedWires[1701]), .A1 (n_0_57), .A2 (opt_ipo_n1525));
NOR2_X1 i_0_874 (.ZN (normalizedWires[1700]), .A1 (n_0_57), .A2 (n_0_11));
NOR2_X1 i_0_873 (.ZN (normalizedWires[1699]), .A1 (n_0_57), .A2 (opt_ipo_n1556));
NOR2_X1 i_0_872 (.ZN (normalizedWires[1698]), .A1 (n_0_57), .A2 (n_0_9));
NOR2_X1 i_0_871 (.ZN (normalizedWires[1697]), .A1 (n_0_57), .A2 (n_0_76));
NOR2_X1 i_0_870 (.ZN (normalizedWires[1696]), .A1 (n_0_57), .A2 (n_0_67));
NOR2_X1 i_0_869 (.ZN (normalizedWires[1695]), .A1 (n_0_57), .A2 (sgo__n175));
NOR2_X1 i_0_868 (.ZN (normalizedWires[1694]), .A1 (n_0_57), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_867 (.ZN (normalizedWires[1693]), .A1 (n_0_57), .A2 (CLOCK_slo___n3082));
NOR2_X1 i_0_866 (.ZN (normalizedWires[1692]), .A1 (n_0_57), .A2 (n_0_3));
NOR2_X1 i_0_865 (.ZN (normalizedWires[1691]), .A1 (n_0_57), .A2 (n_0_2));
NOR2_X1 i_0_864 (.ZN (normalizedWires[1690]), .A1 (n_0_57), .A2 (n_0_73));
INV_X4 i_0_863 (.ZN (n_0_57), .A (B[26]));
NOR2_X1 i_0_862 (.ZN (normalizedWires[1655]), .A1 (n_0_56), .A2 (slo__n785));
NOR2_X1 i_0_861 (.ZN (normalizedWires[1654]), .A1 (n_0_56), .A2 (slo__n332));
NOR2_X1 i_0_860 (.ZN (normalizedWires[1653]), .A1 (n_0_56), .A2 (sgo__n131));
NOR2_X1 i_0_859 (.ZN (normalizedWires[1652]), .A1 (n_0_56), .A2 (opt_ipo_n1675));
NOR2_X1 i_0_858 (.ZN (normalizedWires[1651]), .A1 (n_0_27), .A2 (n_0_56));
NOR2_X1 i_0_857 (.ZN (normalizedWires[1650]), .A1 (n_0_56), .A2 (CLOCK_slo__n3096));
NOR2_X1 i_0_856 (.ZN (normalizedWires[1649]), .A1 (n_0_56), .A2 (n_0_25));
NOR2_X1 i_0_855 (.ZN (normalizedWires[1648]), .A1 (n_0_56), .A2 (opt_ipo_n1532));
NOR2_X2 CLOCK_slo__mro_c2640 (.ZN (normalizedWires[1628]), .A1 (n_0_56), .A2 (CLOCK_slo___n3082));
NOR2_X2 slo__mro_c340 (.ZN (normalizedWires[271]), .A1 (n_0_12), .A2 (n_0_35));
NOR2_X2 i_0_850 (.ZN (normalizedWires[1643]), .A1 (n_0_56), .A2 (n_0_19));
NOR2_X2 i_0_849 (.ZN (normalizedWires[1642]), .A1 (n_0_56), .A2 (slo___n436));
NOR2_X1 i_0_848 (.ZN (normalizedWires[1641]), .A1 (n_0_56), .A2 (opt_ipo_n1550));
NOR2_X2 i_0_847 (.ZN (normalizedWires[1640]), .A1 (n_0_56), .A2 (n_0_16));
NOR2_X1 i_0_846 (.ZN (normalizedWires[1639]), .A1 (n_0_56), .A2 (n_0_15));
NOR2_X1 i_0_845 (.ZN (normalizedWires[1638]), .A1 (n_0_56), .A2 (n_0_14));
NOR2_X1 i_0_844 (.ZN (normalizedWires[1637]), .A1 (n_0_56), .A2 (n_0_13));
NOR2_X1 i_0_843 (.ZN (normalizedWires[1636]), .A1 (n_0_56), .A2 (n_0_12));
NOR2_X1 i_0_842 (.ZN (normalizedWires[1635]), .A1 (n_0_56), .A2 (n_0_11));
NOR2_X1 i_0_841 (.ZN (normalizedWires[1634]), .A1 (n_0_56), .A2 (n_0_10));
NOR2_X1 i_0_840 (.ZN (normalizedWires[1633]), .A1 (n_0_56), .A2 (n_0_9));
NOR2_X1 i_0_832 (.ZN (normalizedWires[1625]), .A1 (n_0_56), .A2 (n_0_73));
NOR2_X1 i_0_830 (.ZN (normalizedWires[1590]), .A1 (slo__n1306), .A2 (slo__n785));
NOR2_X4 i_0_829 (.ZN (normalizedWires[1589]), .A1 (slo__n1306), .A2 (slo__n332));
NOR2_X1 i_0_828 (.ZN (normalizedWires[1588]), .A1 (slo__n1306), .A2 (sgo__n131));
NOR2_X2 i_0_827 (.ZN (normalizedWires[1587]), .A1 (n_0_55), .A2 (n_0_28));
NOR2_X2 i_0_826 (.ZN (normalizedWires[1586]), .A1 (n_0_55), .A2 (n_0_27));
NOR2_X1 i_0_825 (.ZN (normalizedWires[1585]), .A1 (n_0_55), .A2 (n_0_26));
NOR2_X1 i_0_824 (.ZN (normalizedWires[1584]), .A1 (n_0_55), .A2 (n_0_25));
NOR2_X2 i_0_823 (.ZN (normalizedWires[1583]), .A1 (n_0_55), .A2 (opt_ipo_n1532));
NOR2_X2 i_0_820 (.ZN (normalizedWires[1580]), .A1 (n_0_55), .A2 (n_0_21));
NOR2_X1 i_0_819 (.ZN (normalizedWires[1579]), .A1 (n_0_55), .A2 (n_0_20));
NOR2_X1 i_0_818 (.ZN (normalizedWires[1578]), .A1 (n_0_55), .A2 (n_0_19));
NOR2_X1 i_0_817 (.ZN (normalizedWires[1577]), .A1 (n_0_55), .A2 (slo__n381));
NOR2_X2 i_0_816 (.ZN (normalizedWires[1576]), .A1 (opt_ipo_n1550), .A2 (n_0_55));
NOR2_X2 i_0_815 (.ZN (normalizedWires[1575]), .A1 (n_0_55), .A2 (n_0_16));
NOR2_X1 i_0_814 (.ZN (normalizedWires[1574]), .A1 (n_0_55), .A2 (n_0_15));
NOR2_X2 i_0_813 (.ZN (normalizedWires[1573]), .A1 (n_0_55), .A2 (n_0_14));
NOR2_X1 i_0_812 (.ZN (normalizedWires[1572]), .A1 (n_0_55), .A2 (n_0_13));
NOR2_X1 i_0_811 (.ZN (normalizedWires[1571]), .A1 (n_0_55), .A2 (n_0_12));
NOR2_X2 i_0_810 (.ZN (normalizedWires[1570]), .A1 (n_0_55), .A2 (n_0_11));
NOR2_X1 i_0_809 (.ZN (normalizedWires[1569]), .A1 (n_0_55), .A2 (n_0_10));
NOR2_X2 i_0_808 (.ZN (normalizedWires[1568]), .A1 (n_0_55), .A2 (n_0_9));
NOR2_X2 i_0_807 (.ZN (normalizedWires[1567]), .A1 (n_0_55), .A2 (n_0_76));
NOR2_X1 i_0_806 (.ZN (normalizedWires[1566]), .A1 (n_0_55), .A2 (n_0_67));
NOR2_X1 i_0_805 (.ZN (normalizedWires[1565]), .A1 (n_0_55), .A2 (sgo__n175));
NOR2_X1 i_0_804 (.ZN (normalizedWires[1564]), .A1 (n_0_55), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_803 (.ZN (normalizedWires[1563]), .A1 (n_0_55), .A2 (CLOCK_slo___n3082));
NOR2_X1 i_0_802 (.ZN (normalizedWires[1562]), .A1 (n_0_55), .A2 (n_0_3));
NOR2_X1 i_0_801 (.ZN (normalizedWires[1561]), .A1 (slo__n1306), .A2 (n_0_2));
NOR2_X1 i_0_800 (.ZN (normalizedWires[1560]), .A1 (slo__n1306), .A2 (n_0_73));
NOR2_X1 i_0_798 (.ZN (normalizedWires[1525]), .A1 (n_0_54), .A2 (slo__n785));
NOR2_X1 i_0_797 (.ZN (normalizedWires[1524]), .A1 (n_0_54), .A2 (slo__n332));
NOR2_X1 i_0_796 (.ZN (normalizedWires[1523]), .A1 (n_0_54), .A2 (sgo__n131));
NOR2_X1 i_0_795 (.ZN (normalizedWires[1522]), .A1 (n_0_54), .A2 (opt_ipo_n1675));
NOR2_X1 i_0_794 (.ZN (normalizedWires[1521]), .A1 (n_0_54), .A2 (sgo__n168));
NOR2_X1 i_0_793 (.ZN (normalizedWires[1520]), .A1 (n_0_54), .A2 (sgo__n27));
NOR2_X1 i_0_792 (.ZN (normalizedWires[1519]), .A1 (n_0_54), .A2 (opt_ipo_n1677));
NOR2_X1 i_0_791 (.ZN (normalizedWires[1518]), .A1 (n_0_54), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_790 (.ZN (normalizedWires[1517]), .A1 (n_0_54), .A2 (n_0_23));
NOR2_X1 i_0_789 (.ZN (normalizedWires[1516]), .A1 (n_0_54), .A2 (slo__n302));
NOR2_X1 i_0_788 (.ZN (normalizedWires[1515]), .A1 (n_0_54), .A2 (n_0_21));
NOR2_X1 i_0_787 (.ZN (normalizedWires[1514]), .A1 (n_0_54), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_786 (.ZN (normalizedWires[1513]), .A1 (n_0_54), .A2 (n_0_19));
NOR2_X1 i_0_785 (.ZN (normalizedWires[1512]), .A1 (n_0_54), .A2 (slo__n298));
NOR2_X1 i_0_784 (.ZN (normalizedWires[1511]), .A1 (n_0_54), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_783 (.ZN (normalizedWires[1510]), .A1 (n_0_54), .A2 (n_0_16));
NOR2_X1 i_0_782 (.ZN (normalizedWires[1509]), .A1 (n_0_54), .A2 (CLOCK_sgo__n1891));
NOR2_X1 i_0_781 (.ZN (normalizedWires[1508]), .A1 (n_0_54), .A2 (n_0_14));
NOR2_X1 i_0_780 (.ZN (normalizedWires[1507]), .A1 (n_0_54), .A2 (CLOCK_sgo__n1896));
NOR2_X1 i_0_779 (.ZN (normalizedWires[1506]), .A1 (n_0_54), .A2 (opt_ipo_n1525));
NOR2_X1 i_0_778 (.ZN (normalizedWires[1505]), .A1 (n_0_54), .A2 (n_0_11));
NOR2_X1 i_0_777 (.ZN (normalizedWires[1504]), .A1 (n_0_54), .A2 (opt_ipo_n1556));
NOR2_X1 i_0_776 (.ZN (normalizedWires[1503]), .A1 (n_0_54), .A2 (n_0_9));
NOR2_X1 i_0_775 (.ZN (normalizedWires[1502]), .A1 (n_0_54), .A2 (slo__n1013));
NOR2_X1 i_0_774 (.ZN (normalizedWires[1501]), .A1 (n_0_54), .A2 (n_0_67));
NOR2_X1 i_0_773 (.ZN (normalizedWires[1500]), .A1 (n_0_54), .A2 (sgo__n175));
NOR2_X1 i_0_772 (.ZN (normalizedWires[1499]), .A1 (n_0_54), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_771 (.ZN (normalizedWires[1498]), .A1 (n_0_54), .A2 (CLOCK_slo___n3082));
NOR2_X1 i_0_770 (.ZN (normalizedWires[1497]), .A1 (n_0_54), .A2 (n_0_3));
NOR2_X1 i_0_769 (.ZN (normalizedWires[1496]), .A1 (n_0_54), .A2 (n_0_2));
NOR2_X1 i_0_768 (.ZN (normalizedWires[1495]), .A1 (n_0_54), .A2 (n_0_73));
INV_X4 i_0_767 (.ZN (n_0_54), .A (B[23]));
NOR2_X1 i_0_766 (.ZN (normalizedWires[1460]), .A1 (n_0_53), .A2 (slo__n785));
NOR2_X1 i_0_765 (.ZN (normalizedWires[1459]), .A1 (n_0_53), .A2 (slo__n332));
NOR2_X1 i_0_764 (.ZN (normalizedWires[1458]), .A1 (n_0_53), .A2 (n_0_29));
NOR2_X1 i_0_763 (.ZN (normalizedWires[1457]), .A1 (n_0_53), .A2 (n_0_28));
NOR2_X1 i_0_762 (.ZN (normalizedWires[1456]), .A1 (n_0_53), .A2 (n_0_27));
NOR2_X1 i_0_760 (.ZN (normalizedWires[1454]), .A1 (n_0_53), .A2 (n_0_25));
NOR2_X1 i_0_759 (.ZN (normalizedWires[1453]), .A1 (n_0_53), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_756 (.ZN (normalizedWires[1450]), .A1 (n_0_53), .A2 (n_0_21));
NOR2_X1 i_0_755 (.ZN (normalizedWires[1449]), .A1 (n_0_53), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_754 (.ZN (normalizedWires[1448]), .A1 (n_0_53), .A2 (n_0_19));
NOR2_X1 i_0_753 (.ZN (normalizedWires[1447]), .A1 (slo___n436), .A2 (n_0_53));
NOR2_X1 i_0_752 (.ZN (normalizedWires[1446]), .A1 (n_0_53), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_751 (.ZN (normalizedWires[1445]), .A1 (n_0_53), .A2 (n_0_16));
NOR2_X1 i_0_750 (.ZN (normalizedWires[1444]), .A1 (n_0_53), .A2 (n_0_15));
NOR2_X1 i_0_749 (.ZN (normalizedWires[1443]), .A1 (n_0_53), .A2 (n_0_14));
NOR2_X1 i_0_748 (.ZN (normalizedWires[1442]), .A1 (n_0_53), .A2 (n_0_13));
NOR2_X1 i_0_747 (.ZN (normalizedWires[1441]), .A1 (n_0_53), .A2 (n_0_12));
NOR2_X1 i_0_746 (.ZN (normalizedWires[1440]), .A1 (n_0_53), .A2 (n_0_11));
NOR2_X1 i_0_745 (.ZN (normalizedWires[1439]), .A1 (n_0_53), .A2 (n_0_10));
NOR2_X4 i_0_744 (.ZN (normalizedWires[1438]), .A1 (n_0_53), .A2 (n_0_9));
NOR2_X1 i_0_743 (.ZN (normalizedWires[1437]), .A1 (n_0_53), .A2 (n_0_76));
NOR2_X1 i_0_742 (.ZN (normalizedWires[1436]), .A1 (n_0_53), .A2 (n_0_67));
NOR2_X1 i_0_741 (.ZN (normalizedWires[1435]), .A1 (n_0_53), .A2 (sgo__n175));
NOR2_X1 i_0_740 (.ZN (normalizedWires[1434]), .A1 (n_0_53), .A2 (n_0_5));
NOR2_X1 i_0_739 (.ZN (normalizedWires[1433]), .A1 (n_0_53), .A2 (CLOCK_slo___n3082));
NOR2_X1 i_0_738 (.ZN (normalizedWires[1432]), .A1 (n_0_53), .A2 (n_0_3));
NOR2_X1 i_0_737 (.ZN (normalizedWires[1431]), .A1 (n_0_53), .A2 (n_0_2));
NOR2_X1 i_0_736 (.ZN (normalizedWires[1430]), .A1 (n_0_53), .A2 (n_0_73));
NOR2_X1 i_0_734 (.ZN (normalizedWires[1395]), .A1 (n_0_52), .A2 (slo__n785));
NOR2_X1 i_0_733 (.ZN (normalizedWires[1394]), .A1 (n_0_52), .A2 (n_0_30));
NOR2_X1 i_0_732 (.ZN (normalizedWires[1393]), .A1 (n_0_52), .A2 (n_0_29));
NOR2_X1 i_0_731 (.ZN (normalizedWires[1392]), .A1 (n_0_52), .A2 (n_0_28));
NOR2_X1 i_0_729 (.ZN (normalizedWires[1390]), .A1 (n_0_52), .A2 (n_0_26));
NOR2_X1 i_0_728 (.ZN (normalizedWires[1389]), .A1 (n_0_52), .A2 (n_0_25));
NOR2_X1 i_0_727 (.ZN (normalizedWires[1388]), .A1 (n_0_52), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_724 (.ZN (normalizedWires[1385]), .A1 (n_0_52), .A2 (n_0_21));
NOR2_X2 i_0_723 (.ZN (normalizedWires[1384]), .A1 (n_0_52), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_722 (.ZN (normalizedWires[1383]), .A1 (n_0_52), .A2 (n_0_19));
NOR2_X1 i_0_721 (.ZN (normalizedWires[1382]), .A1 (n_0_52), .A2 (slo___n436));
NOR2_X1 i_0_720 (.ZN (normalizedWires[1381]), .A1 (n_0_52), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_719 (.ZN (normalizedWires[1380]), .A1 (n_0_52), .A2 (n_0_16));
NOR2_X1 i_0_718 (.ZN (normalizedWires[1379]), .A1 (n_0_52), .A2 (n_0_15));
NOR2_X1 i_0_717 (.ZN (normalizedWires[1378]), .A1 (n_0_52), .A2 (n_0_14));
NOR2_X1 i_0_716 (.ZN (normalizedWires[1377]), .A1 (n_0_52), .A2 (n_0_13));
NOR2_X1 i_0_715 (.ZN (normalizedWires[1376]), .A1 (n_0_52), .A2 (n_0_12));
NOR2_X1 i_0_714 (.ZN (normalizedWires[1375]), .A1 (n_0_52), .A2 (n_0_11));
NOR2_X1 slo__sro_c677 (.ZN (normalizedWires[661]), .A1 (n_0_12), .A2 (opt_ipo_n1649));
NOR2_X1 i_0_712 (.ZN (normalizedWires[1373]), .A1 (n_0_52), .A2 (n_0_9));
NOR2_X1 i_0_711 (.ZN (normalizedWires[1372]), .A1 (n_0_52), .A2 (n_0_76));
NOR2_X1 i_0_710 (.ZN (normalizedWires[1371]), .A1 (n_0_52), .A2 (n_0_67));
NOR2_X1 i_0_709 (.ZN (normalizedWires[1370]), .A1 (n_0_52), .A2 (sgo__n175));
CLKBUF_X2 CLOCK_slo__c2494 (.Z (CLOCK_slo__n2695), .A (n_0_12));
NOR2_X1 i_0_707 (.ZN (normalizedWires[1368]), .A1 (n_0_52), .A2 (CLOCK_slo___n3082));
NOR2_X1 i_0_706 (.ZN (normalizedWires[1367]), .A1 (n_0_52), .A2 (n_0_3));
NOR2_X1 i_0_705 (.ZN (normalizedWires[1366]), .A1 (n_0_52), .A2 (n_0_2));
NOR2_X1 i_0_704 (.ZN (normalizedWires[1365]), .A1 (n_0_52), .A2 (n_0_73));
NOR2_X1 i_0_702 (.ZN (normalizedWires[1330]), .A1 (n_0_51), .A2 (slo__n785));
NOR2_X1 i_0_701 (.ZN (normalizedWires[1329]), .A1 (n_0_51), .A2 (slo__n332));
NOR2_X1 i_0_700 (.ZN (normalizedWires[1328]), .A1 (n_0_51), .A2 (sgo__n131));
NOR2_X1 i_0_699 (.ZN (normalizedWires[1327]), .A1 (n_0_51), .A2 (opt_ipo_n1675));
NOR2_X1 i_0_698 (.ZN (normalizedWires[1326]), .A1 (n_0_51), .A2 (sgo__n168));
NOR2_X1 i_0_697 (.ZN (normalizedWires[1325]), .A1 (n_0_51), .A2 (sgo__n27));
NOR2_X1 i_0_696 (.ZN (normalizedWires[1324]), .A1 (n_0_51), .A2 (opt_ipo_n1677));
NOR2_X1 i_0_695 (.ZN (normalizedWires[1323]), .A1 (n_0_51), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_694 (.ZN (normalizedWires[1322]), .A1 (n_0_51), .A2 (n_0_23));
NOR2_X1 i_0_693 (.ZN (normalizedWires[1321]), .A1 (n_0_51), .A2 (slo__n302));
NOR2_X1 i_0_692 (.ZN (normalizedWires[1320]), .A1 (n_0_51), .A2 (n_0_21));
NOR2_X1 i_0_691 (.ZN (normalizedWires[1319]), .A1 (n_0_51), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_690 (.ZN (normalizedWires[1318]), .A1 (n_0_51), .A2 (n_0_19));
NOR2_X1 i_0_689 (.ZN (normalizedWires[1317]), .A1 (n_0_51), .A2 (slo__n298));
NOR2_X1 i_0_688 (.ZN (normalizedWires[1316]), .A1 (n_0_51), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_687 (.ZN (normalizedWires[1315]), .A1 (n_0_51), .A2 (n_0_16));
NOR2_X1 i_0_686 (.ZN (normalizedWires[1314]), .A1 (n_0_51), .A2 (CLOCK_sgo__n1891));
NOR2_X1 i_0_685 (.ZN (normalizedWires[1313]), .A1 (n_0_51), .A2 (n_0_14));
NOR2_X1 i_0_684 (.ZN (normalizedWires[1312]), .A1 (n_0_51), .A2 (n_0_13));
NOR2_X1 i_0_683 (.ZN (normalizedWires[1311]), .A1 (n_0_51), .A2 (opt_ipo_n1525));
NOR2_X1 i_0_682 (.ZN (normalizedWires[1310]), .A1 (n_0_51), .A2 (n_0_11));
NOR2_X1 i_0_681 (.ZN (normalizedWires[1309]), .A1 (n_0_51), .A2 (opt_ipo_n1556));
NOR2_X1 i_0_680 (.ZN (normalizedWires[1308]), .A1 (n_0_51), .A2 (n_0_9));
NOR2_X1 i_0_679 (.ZN (normalizedWires[1307]), .A1 (n_0_51), .A2 (n_0_76));
NOR2_X1 i_0_678 (.ZN (normalizedWires[1306]), .A1 (n_0_51), .A2 (n_0_67));
NOR2_X1 i_0_677 (.ZN (normalizedWires[1305]), .A1 (n_0_51), .A2 (sgo__n175));
NOR2_X1 i_0_676 (.ZN (normalizedWires[1304]), .A1 (n_0_51), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_675 (.ZN (normalizedWires[1303]), .A1 (n_0_51), .A2 (CLOCK_slo___n3082));
NOR2_X1 i_0_674 (.ZN (normalizedWires[1302]), .A1 (n_0_51), .A2 (n_0_3));
NOR2_X1 i_0_673 (.ZN (normalizedWires[1301]), .A1 (n_0_51), .A2 (n_0_2));
NOR2_X1 i_0_672 (.ZN (normalizedWires[1300]), .A1 (n_0_51), .A2 (n_0_73));
INV_X4 i_0_671 (.ZN (n_0_51), .A (B[20]));
NOR2_X1 i_0_670 (.ZN (normalizedWires[1265]), .A1 (sgo__n85), .A2 (n_0_31));
NOR2_X1 i_0_669 (.ZN (normalizedWires[1264]), .A1 (n_0_50), .A2 (n_0_30));
NOR2_X1 i_0_668 (.ZN (normalizedWires[1263]), .A1 (n_0_50), .A2 (n_0_29));
NOR2_X1 i_0_667 (.ZN (normalizedWires[1262]), .A1 (n_0_50), .A2 (n_0_28));
NOR2_X2 i_0_664 (.ZN (normalizedWires[1259]), .A1 (n_0_50), .A2 (slo__n1158));
NOR2_X2 CLOCK_slo__sro_c2759 (.ZN (normalizedWires[207]), .A1 (slo__n1127), .A2 (n_0_34));
NOR2_X4 i_0_660 (.ZN (normalizedWires[1255]), .A1 (n_0_21), .A2 (n_0_50));
NOR2_X1 i_0_659 (.ZN (normalizedWires[1254]), .A1 (n_0_50), .A2 (n_0_20));
NOR2_X1 i_0_658 (.ZN (normalizedWires[1253]), .A1 (n_0_50), .A2 (n_0_19));
NOR2_X1 i_0_657 (.ZN (normalizedWires[1252]), .A1 (n_0_50), .A2 (slo__n381));
NOR2_X1 i_0_656 (.ZN (normalizedWires[1251]), .A1 (n_0_50), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_655 (.ZN (normalizedWires[1250]), .A1 (n_0_50), .A2 (n_0_16));
NOR2_X1 i_0_654 (.ZN (normalizedWires[1249]), .A1 (n_0_50), .A2 (n_0_15));
NOR2_X2 i_0_653 (.ZN (normalizedWires[1248]), .A1 (n_0_50), .A2 (n_0_14));
NOR2_X4 CLOCK_slo__mro_c2585 (.ZN (normalizedWires[610]), .A1 (n_0_26), .A2 (n_0_40));
NOR2_X2 i_0_651 (.ZN (normalizedWires[1246]), .A1 (n_0_50), .A2 (n_0_12));
NOR2_X4 i_0_650 (.ZN (normalizedWires[1245]), .A1 (n_0_50), .A2 (n_0_11));
NOR2_X1 i_0_649 (.ZN (normalizedWires[1244]), .A1 (n_0_50), .A2 (n_0_10));
INV_X2 slo__c954 (.ZN (slo__n1036), .A (B[10]));
NOR2_X1 i_0_647 (.ZN (normalizedWires[1242]), .A1 (n_0_50), .A2 (n_0_76));
NOR2_X1 i_0_646 (.ZN (normalizedWires[1241]), .A1 (n_0_50), .A2 (n_0_67));
NOR2_X1 i_0_645 (.ZN (normalizedWires[1240]), .A1 (n_0_50), .A2 (n_0_68));
NOR2_X1 i_0_644 (.ZN (normalizedWires[1239]), .A1 (n_0_50), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_643 (.ZN (normalizedWires[1238]), .A1 (sgo__n85), .A2 (CLOCK_slo___n3082));
NOR2_X1 i_0_642 (.ZN (normalizedWires[1237]), .A1 (sgo__n85), .A2 (n_0_3));
NOR2_X1 i_0_641 (.ZN (normalizedWires[1236]), .A1 (sgo__n85), .A2 (n_0_2));
NOR2_X1 i_0_640 (.ZN (normalizedWires[1235]), .A1 (sgo__n85), .A2 (n_0_73));
NOR2_X1 i_0_638 (.ZN (normalizedWires[1200]), .A1 (n_0_49), .A2 (n_0_31));
NOR2_X1 i_0_637 (.ZN (normalizedWires[1199]), .A1 (n_0_49), .A2 (n_0_30));
NOR2_X1 i_0_636 (.ZN (normalizedWires[1198]), .A1 (n_0_49), .A2 (n_0_29));
NOR2_X2 CLOCK_slo__sro_c2075 (.ZN (normalizedWires[200]), .A1 (n_0_68), .A2 (n_0_34));
INV_X4 CLOCK_slo__c2226 (.ZN (CLOCK_slo__n2403), .A (A[17]));
NOR2_X1 i_0_631 (.ZN (normalizedWires[1193]), .A1 (n_0_49), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_629 (.ZN (normalizedWires[1191]), .A1 (n_0_49), .A2 (n_0_22));
NOR2_X2 i_0_628 (.ZN (normalizedWires[1190]), .A1 (n_0_49), .A2 (n_0_21));
NOR2_X2 i_0_627 (.ZN (normalizedWires[1189]), .A1 (n_0_49), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_626 (.ZN (normalizedWires[1188]), .A1 (n_0_49), .A2 (n_0_19));
NOR2_X1 i_0_625 (.ZN (normalizedWires[1187]), .A1 (n_0_49), .A2 (slo___n436));
NOR2_X1 i_0_624 (.ZN (normalizedWires[1186]), .A1 (n_0_49), .A2 (opt_ipo_n1550));
NOR2_X2 i_0_623 (.ZN (normalizedWires[1185]), .A1 (n_0_49), .A2 (n_0_16));
NOR2_X2 CLOCK_slo__sro_c2044 (.ZN (normalizedWires[1179]), .A1 (n_0_49), .A2 (n_0_10));
CLKBUF_X1 slo___L1_c1_c665 (.Z (slo_n705), .A (B_7_PP_0));
BUF_X1 CLOCK_slo__c2920 (.Z (CLOCK_slo__n3235), .A (n_0_29));
CLKBUF_X1 slo___L1_c1_c1203 (.Z (slo_n1330), .A (B_24_PP_0));
NOR2_X1 CLOCK_slo__mro_c2530 (.ZN (normalizedWires[24]), .A1 (n_0_25), .A2 (n_0_0));
NOR2_X2 CLOCK_slo__sro_c2066 (.ZN (normalizedWires[1197]), .A1 (n_0_49), .A2 (n_0_28));
NOR2_X2 CLOCK_slo__sro_c2038 (.ZN (normalizedWires[1184]), .A1 (n_0_49), .A2 (n_0_15));
NOR2_X1 i_0_615 (.ZN (normalizedWires[1177]), .A1 (n_0_49), .A2 (n_0_76));
NOR2_X1 i_0_614 (.ZN (normalizedWires[1176]), .A1 (n_0_49), .A2 (n_0_67));
NOR2_X1 i_0_613 (.ZN (normalizedWires[1175]), .A1 (n_0_49), .A2 (sgo__n175));
NOR2_X1 i_0_612 (.ZN (normalizedWires[1174]), .A1 (slo___n867), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_611 (.ZN (normalizedWires[1173]), .A1 (slo___n867), .A2 (CLOCK_slo___n3082));
NOR2_X1 i_0_610 (.ZN (normalizedWires[1172]), .A1 (slo___n867), .A2 (n_0_3));
NOR2_X1 i_0_609 (.ZN (normalizedWires[1171]), .A1 (slo___n867), .A2 (n_0_2));
NOR2_X1 i_0_608 (.ZN (normalizedWires[1170]), .A1 (slo___n867), .A2 (n_0_73));
NOR2_X1 i_0_606 (.ZN (normalizedWires[1135]), .A1 (n_0_48), .A2 (slo__n785));
NOR2_X1 i_0_605 (.ZN (normalizedWires[1134]), .A1 (n_0_48), .A2 (slo__n332));
NOR2_X1 i_0_604 (.ZN (normalizedWires[1133]), .A1 (n_0_48), .A2 (sgo__n131));
NOR2_X1 i_0_603 (.ZN (normalizedWires[1132]), .A1 (n_0_48), .A2 (opt_ipo_n1675));
NOR2_X1 i_0_602 (.ZN (normalizedWires[1131]), .A1 (n_0_48), .A2 (n_0_27));
NOR2_X1 i_0_601 (.ZN (normalizedWires[1130]), .A1 (n_0_48), .A2 (n_0_26));
NOR2_X1 i_0_600 (.ZN (normalizedWires[1129]), .A1 (n_0_48), .A2 (n_0_25));
NOR2_X1 i_0_599 (.ZN (normalizedWires[1128]), .A1 (n_0_48), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_598 (.ZN (normalizedWires[1127]), .A1 (n_0_48), .A2 (n_0_23));
NOR2_X1 i_0_597 (.ZN (normalizedWires[1126]), .A1 (n_0_48), .A2 (n_0_22));
NOR2_X1 i_0_596 (.ZN (normalizedWires[1125]), .A1 (n_0_48), .A2 (n_0_21));
NOR2_X1 i_0_595 (.ZN (normalizedWires[1124]), .A1 (n_0_48), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_594 (.ZN (normalizedWires[1123]), .A1 (n_0_48), .A2 (n_0_19));
NOR2_X1 i_0_593 (.ZN (normalizedWires[1122]), .A1 (n_0_48), .A2 (slo__n298));
NOR2_X1 i_0_592 (.ZN (normalizedWires[1121]), .A1 (n_0_48), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_591 (.ZN (normalizedWires[1120]), .A1 (n_0_48), .A2 (n_0_16));
NOR2_X2 i_0_590 (.ZN (normalizedWires[1119]), .A1 (n_0_48), .A2 (CLOCK_sgo__n1891));
NOR2_X1 i_0_589 (.ZN (normalizedWires[1118]), .A1 (n_0_48), .A2 (n_0_14));
NOR2_X1 i_0_588 (.ZN (normalizedWires[1117]), .A1 (n_0_48), .A2 (CLOCK_sgo__n1896));
NOR2_X1 i_0_587 (.ZN (normalizedWires[1116]), .A1 (n_0_48), .A2 (opt_ipo_n1525));
NOR2_X1 i_0_586 (.ZN (normalizedWires[1115]), .A1 (n_0_48), .A2 (n_0_11));
NOR2_X1 i_0_585 (.ZN (normalizedWires[1114]), .A1 (n_0_48), .A2 (opt_ipo_n1556));
NOR2_X1 i_0_584 (.ZN (normalizedWires[1113]), .A1 (n_0_48), .A2 (n_0_9));
NOR2_X1 i_0_583 (.ZN (normalizedWires[1112]), .A1 (n_0_48), .A2 (slo__n1013));
NOR2_X1 i_0_582 (.ZN (normalizedWires[1111]), .A1 (n_0_48), .A2 (n_0_67));
NOR2_X1 i_0_581 (.ZN (normalizedWires[1110]), .A1 (n_0_48), .A2 (sgo__n175));
NOR2_X1 i_0_580 (.ZN (normalizedWires[1109]), .A1 (n_0_48), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_579 (.ZN (normalizedWires[1108]), .A1 (n_0_48), .A2 (n_0_4));
NOR2_X1 i_0_578 (.ZN (normalizedWires[1107]), .A1 (n_0_48), .A2 (n_0_3));
NOR2_X1 i_0_577 (.ZN (normalizedWires[1106]), .A1 (n_0_48), .A2 (n_0_2));
NOR2_X1 i_0_576 (.ZN (normalizedWires[1105]), .A1 (n_0_48), .A2 (n_0_73));
INV_X4 i_0_575 (.ZN (n_0_48), .A (B[17]));
NOR2_X1 i_0_574 (.ZN (normalizedWires[1070]), .A1 (CLOCK_slo__n2299), .A2 (slo__n785));
NOR2_X1 i_0_573 (.ZN (normalizedWires[1069]), .A1 (CLOCK_slo__n2299), .A2 (slo__n332));
NOR2_X1 i_0_572 (.ZN (normalizedWires[1068]), .A1 (sgo__n131), .A2 (n_0_47));
NOR2_X2 slo__sro_c939 (.ZN (normalizedWires[1243]), .A1 (n_0_50), .A2 (n_0_9));
NOR2_X1 i_0_567 (.ZN (normalizedWires[1063]), .A1 (opt_ipo_n1532), .A2 (n_0_47));
NOR2_X1 i_0_565 (.ZN (normalizedWires[1061]), .A1 (CLOCK_slo__n2299), .A2 (n_0_22));
NOR2_X1 i_0_564 (.ZN (normalizedWires[1060]), .A1 (n_0_47), .A2 (n_0_21));
NOR2_X1 i_0_563 (.ZN (normalizedWires[1059]), .A1 (n_0_47), .A2 (n_0_20));
NOR2_X4 i_0_562 (.ZN (normalizedWires[1058]), .A1 (n_0_47), .A2 (n_0_19));
NOR2_X4 i_0_561 (.ZN (normalizedWires[1057]), .A1 (n_0_47), .A2 (slo___n436));
NOR2_X4 i_0_560 (.ZN (normalizedWires[1056]), .A1 (n_0_47), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_559 (.ZN (normalizedWires[1055]), .A1 (n_0_47), .A2 (n_0_16));
NOR2_X1 i_0_558 (.ZN (normalizedWires[1054]), .A1 (n_0_47), .A2 (n_0_15));
NOR2_X1 i_0_557 (.ZN (normalizedWires[1053]), .A1 (n_0_47), .A2 (n_0_14));
NOR2_X1 i_0_556 (.ZN (normalizedWires[1052]), .A1 (n_0_47), .A2 (slo__n1127));
NOR2_X1 i_0_555 (.ZN (normalizedWires[1051]), .A1 (n_0_47), .A2 (n_0_12));
NOR2_X1 i_0_554 (.ZN (normalizedWires[1050]), .A1 (n_0_47), .A2 (n_0_11));
NOR2_X1 i_0_553 (.ZN (normalizedWires[1049]), .A1 (n_0_47), .A2 (n_0_10));
NOR2_X1 i_0_552 (.ZN (normalizedWires[1048]), .A1 (n_0_47), .A2 (n_0_9));
NOR2_X1 i_0_551 (.ZN (normalizedWires[1047]), .A1 (n_0_47), .A2 (n_0_76));
NOR2_X1 i_0_550 (.ZN (normalizedWires[1046]), .A1 (n_0_47), .A2 (n_0_67));
NOR2_X1 i_0_549 (.ZN (normalizedWires[1045]), .A1 (n_0_47), .A2 (sgo__n175));
NOR2_X1 i_0_548 (.ZN (normalizedWires[1044]), .A1 (n_0_47), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_547 (.ZN (normalizedWires[1043]), .A1 (n_0_47), .A2 (CLOCK_slo___n3081));
NOR2_X1 i_0_546 (.ZN (normalizedWires[1042]), .A1 (n_0_47), .A2 (n_0_3));
NOR2_X2 CLOCK_slo__sro_c2168 (.ZN (normalizedWires[1194]), .A1 (n_0_25), .A2 (n_0_49));
NOR2_X1 i_0_544 (.ZN (normalizedWires[1040]), .A1 (n_0_47), .A2 (n_0_73));
NOR2_X1 i_0_542 (.ZN (normalizedWires[1005]), .A1 (n_0_46), .A2 (slo__n785));
NOR2_X2 i_0_541 (.ZN (normalizedWires[1004]), .A1 (n_0_46), .A2 (slo__n332));
NOR2_X4 i_0_540 (.ZN (normalizedWires[1003]), .A1 (n_0_46), .A2 (n_0_29));
NOR2_X2 i_0_537 (.ZN (normalizedWires[1000]), .A1 (CLOCK_slo__n3096), .A2 (n_0_46));
NOR2_X1 i_0_536 (.ZN (normalizedWires[999]), .A1 (n_0_46), .A2 (slo__n1158));
NOR2_X2 i_0_535 (.ZN (normalizedWires[998]), .A1 (n_0_46), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_533 (.ZN (normalizedWires[996]), .A1 (slo__n1004), .A2 (n_0_22));
NOR2_X2 i_0_532 (.ZN (normalizedWires[995]), .A1 (slo__n1004), .A2 (n_0_21));
NOR2_X1 i_0_531 (.ZN (normalizedWires[994]), .A1 (n_0_46), .A2 (n_0_20));
NOR2_X2 i_0_530 (.ZN (normalizedWires[993]), .A1 (n_0_46), .A2 (n_0_19));
NOR2_X2 i_0_529 (.ZN (normalizedWires[992]), .A1 (n_0_46), .A2 (slo___n436));
NOR2_X1 i_0_528 (.ZN (normalizedWires[991]), .A1 (n_0_46), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_527 (.ZN (normalizedWires[990]), .A1 (CLOCK_slo__n3319), .A2 (n_0_16));
NOR2_X1 i_0_526 (.ZN (normalizedWires[989]), .A1 (CLOCK_slo__n3319), .A2 (n_0_15));
NOR2_X1 i_0_525 (.ZN (normalizedWires[988]), .A1 (n_0_46), .A2 (n_0_14));
NOR2_X1 i_0_524 (.ZN (normalizedWires[987]), .A1 (n_0_46), .A2 (n_0_13));
NOR2_X2 slo__mro_c454 (.ZN (normalizedWires[591]), .A1 (n_0_67), .A2 (n_0_40));
NOR2_X1 i_0_522 (.ZN (normalizedWires[985]), .A1 (n_0_46), .A2 (n_0_11));
NOR2_X1 i_0_521 (.ZN (normalizedWires[984]), .A1 (slo__n1004), .A2 (n_0_10));
NOR2_X1 i_0_520 (.ZN (normalizedWires[983]), .A1 (slo__n1004), .A2 (n_0_9));
NOR2_X1 i_0_519 (.ZN (normalizedWires[982]), .A1 (CLOCK_slo__n3319), .A2 (n_0_76));
NOR2_X1 i_0_518 (.ZN (normalizedWires[981]), .A1 (CLOCK_slo__n3319), .A2 (n_0_67));
NOR2_X4 i_0_517 (.ZN (normalizedWires[980]), .A1 (n_0_46), .A2 (sgo__n175));
NOR2_X1 i_0_516 (.ZN (normalizedWires[979]), .A1 (n_0_46), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_515 (.ZN (normalizedWires[978]), .A1 (n_0_46), .A2 (CLOCK_slo___n3081));
NOR2_X1 i_0_514 (.ZN (normalizedWires[977]), .A1 (n_0_46), .A2 (n_0_3));
NOR2_X1 i_0_513 (.ZN (normalizedWires[976]), .A1 (n_0_46), .A2 (n_0_2));
NOR2_X1 i_0_512 (.ZN (normalizedWires[975]), .A1 (n_0_46), .A2 (n_0_73));
NOR2_X1 i_0_510 (.ZN (normalizedWires[940]), .A1 (n_0_45), .A2 (slo__n785));
NOR2_X1 i_0_509 (.ZN (normalizedWires[939]), .A1 (n_0_45), .A2 (slo__n332));
NOR2_X1 i_0_508 (.ZN (normalizedWires[938]), .A1 (n_0_45), .A2 (CLOCK_slo__n3235));
NOR2_X4 i_0_507 (.ZN (normalizedWires[937]), .A1 (n_0_45), .A2 (opt_ipo_n1675));
NOR2_X1 i_0_506 (.ZN (normalizedWires[936]), .A1 (n_0_45), .A2 (n_0_27));
NOR2_X1 i_0_505 (.ZN (normalizedWires[935]), .A1 (n_0_45), .A2 (n_0_26));
NOR2_X1 i_0_504 (.ZN (normalizedWires[934]), .A1 (n_0_45), .A2 (opt_ipo_n1677));
NOR2_X1 i_0_503 (.ZN (normalizedWires[933]), .A1 (n_0_45), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_502 (.ZN (normalizedWires[932]), .A1 (n_0_45), .A2 (n_0_23));
NOR2_X1 i_0_501 (.ZN (normalizedWires[931]), .A1 (n_0_45), .A2 (n_0_22));
NOR2_X1 i_0_500 (.ZN (normalizedWires[930]), .A1 (n_0_45), .A2 (n_0_21));
NOR2_X1 i_0_499 (.ZN (normalizedWires[929]), .A1 (n_0_45), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_498 (.ZN (normalizedWires[928]), .A1 (n_0_45), .A2 (n_0_19));
NOR2_X1 i_0_497 (.ZN (normalizedWires[927]), .A1 (n_0_45), .A2 (slo__n298));
NOR2_X1 i_0_496 (.ZN (normalizedWires[926]), .A1 (n_0_45), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_495 (.ZN (normalizedWires[925]), .A1 (n_0_45), .A2 (n_0_16));
NOR2_X1 i_0_494 (.ZN (normalizedWires[924]), .A1 (n_0_45), .A2 (CLOCK_sgo__n1891));
NOR2_X1 i_0_493 (.ZN (normalizedWires[923]), .A1 (n_0_45), .A2 (n_0_14));
NOR2_X1 i_0_492 (.ZN (normalizedWires[922]), .A1 (n_0_45), .A2 (CLOCK_sgo__n1896));
NOR2_X1 i_0_491 (.ZN (normalizedWires[921]), .A1 (n_0_45), .A2 (opt_ipo_n1525));
NOR2_X1 i_0_490 (.ZN (normalizedWires[920]), .A1 (n_0_45), .A2 (n_0_11));
NOR2_X1 i_0_489 (.ZN (normalizedWires[919]), .A1 (n_0_45), .A2 (opt_ipo_n1556));
NOR2_X1 i_0_488 (.ZN (normalizedWires[918]), .A1 (n_0_45), .A2 (n_0_9));
NOR2_X1 i_0_487 (.ZN (normalizedWires[917]), .A1 (n_0_45), .A2 (slo__n1013));
NOR2_X1 i_0_486 (.ZN (normalizedWires[916]), .A1 (n_0_45), .A2 (n_0_67));
NOR2_X1 i_0_485 (.ZN (normalizedWires[915]), .A1 (n_0_45), .A2 (sgo__n175));
NOR2_X1 i_0_484 (.ZN (normalizedWires[914]), .A1 (n_0_45), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_483 (.ZN (normalizedWires[913]), .A1 (n_0_45), .A2 (n_0_4));
NOR2_X1 i_0_482 (.ZN (normalizedWires[912]), .A1 (n_0_45), .A2 (n_0_3));
NOR2_X1 i_0_481 (.ZN (normalizedWires[911]), .A1 (n_0_45), .A2 (n_0_2));
NOR2_X1 i_0_480 (.ZN (normalizedWires[910]), .A1 (n_0_45), .A2 (n_0_73));
INV_X4 i_0_479 (.ZN (n_0_45), .A (B[14]));
NOR2_X1 i_0_478 (.ZN (normalizedWires[875]), .A1 (n_0_44), .A2 (slo__n785));
NOR2_X1 slo__sro_c1094 (.ZN (normalizedWires[464]), .A1 (n_0_38), .A2 (slo__n1191));
NOR2_X2 i_0_476 (.ZN (normalizedWires[873]), .A1 (n_0_44), .A2 (n_0_29));
NOR2_X4 i_0_475 (.ZN (normalizedWires[872]), .A1 (n_0_44), .A2 (n_0_28));
NOR2_X2 i_0_474 (.ZN (normalizedWires[871]), .A1 (n_0_44), .A2 (n_0_27));
NOR2_X1 i_0_473 (.ZN (normalizedWires[870]), .A1 (n_0_44), .A2 (n_0_26));
NOR2_X4 slo__sro_c1080 (.ZN (normalizedWires[874]), .A1 (n_0_30), .A2 (n_0_44));
NOR2_X1 i_0_471 (.ZN (normalizedWires[868]), .A1 (n_0_44), .A2 (opt_ipo_n1532));
NOR2_X2 i_0_470 (.ZN (normalizedWires[867]), .A1 (n_0_44), .A2 (n_0_23));
NOR2_X1 i_0_469 (.ZN (normalizedWires[866]), .A1 (n_0_44), .A2 (n_0_22));
NOR2_X1 i_0_468 (.ZN (normalizedWires[865]), .A1 (n_0_44), .A2 (n_0_21));
NOR2_X1 i_0_467 (.ZN (normalizedWires[864]), .A1 (n_0_44), .A2 (n_0_20));
NOR2_X4 i_0_466 (.ZN (normalizedWires[863]), .A1 (n_0_44), .A2 (n_0_19));
NOR2_X1 i_0_465 (.ZN (normalizedWires[862]), .A1 (n_0_44), .A2 (slo___n436));
NOR2_X1 i_0_464 (.ZN (normalizedWires[861]), .A1 (n_0_44), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_463 (.ZN (normalizedWires[860]), .A1 (n_0_44), .A2 (n_0_16));
NOR2_X1 i_0_462 (.ZN (normalizedWires[859]), .A1 (n_0_44), .A2 (n_0_15));
NOR2_X1 i_0_461 (.ZN (normalizedWires[858]), .A1 (n_0_44), .A2 (n_0_14));
NOR2_X1 i_0_460 (.ZN (normalizedWires[857]), .A1 (n_0_44), .A2 (slo__n1127));
NOR2_X1 i_0_459 (.ZN (normalizedWires[856]), .A1 (n_0_44), .A2 (n_0_12));
NOR2_X1 i_0_458 (.ZN (normalizedWires[855]), .A1 (n_0_44), .A2 (n_0_11));
NOR2_X1 i_0_457 (.ZN (normalizedWires[854]), .A1 (n_0_44), .A2 (n_0_10));
NOR2_X1 i_0_456 (.ZN (normalizedWires[853]), .A1 (n_0_44), .A2 (n_0_9));
NOR2_X1 i_0_455 (.ZN (normalizedWires[852]), .A1 (n_0_44), .A2 (n_0_76));
NOR2_X1 i_0_454 (.ZN (normalizedWires[851]), .A1 (n_0_44), .A2 (n_0_67));
NOR2_X1 i_0_453 (.ZN (normalizedWires[850]), .A1 (n_0_44), .A2 (sgo__n175));
NOR2_X1 i_0_452 (.ZN (normalizedWires[849]), .A1 (n_0_44), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_451 (.ZN (normalizedWires[848]), .A1 (n_0_44), .A2 (n_0_4));
NOR2_X1 i_0_450 (.ZN (normalizedWires[847]), .A1 (n_0_44), .A2 (n_0_3));
NOR2_X1 i_0_449 (.ZN (normalizedWires[846]), .A1 (n_0_44), .A2 (n_0_2));
NOR2_X1 i_0_448 (.ZN (normalizedWires[845]), .A1 (n_0_44), .A2 (n_0_73));
INV_X8 i_0_447 (.ZN (n_0_44), .A (B[13]));
NOR2_X1 CLOCK_slo__sro_c2257 (.ZN (normalizedWires[145]), .A1 (n_0_16), .A2 (n_0_33));
NOR2_X4 i_0_445 (.ZN (normalizedWires[809]), .A1 (CLOCK_slo__n2241), .A2 (n_0_30));
NOR2_X1 i_0_444 (.ZN (normalizedWires[808]), .A1 (n_0_43), .A2 (n_0_29));
NOR2_X2 i_0_443 (.ZN (normalizedWires[807]), .A1 (n_0_43), .A2 (n_0_28));
NOR2_X4 i_0_442 (.ZN (normalizedWires[806]), .A1 (n_0_43), .A2 (n_0_27));
NOR2_X2 i_0_441 (.ZN (normalizedWires[805]), .A1 (n_0_43), .A2 (n_0_26));
NOR2_X1 slo__sro_c784 (.ZN (normalizedWires[798]), .A1 (CLOCK_slo__n2241), .A2 (n_0_19));
NOR2_X1 i_0_439 (.ZN (normalizedWires[803]), .A1 (CLOCK_slo__n2241), .A2 (opt_ipo_n1532));
NOR2_X2 i_0_438 (.ZN (normalizedWires[802]), .A1 (n_0_43), .A2 (n_0_23));
NOR2_X1 i_0_437 (.ZN (normalizedWires[801]), .A1 (n_0_43), .A2 (n_0_22));
NOR2_X1 i_0_436 (.ZN (normalizedWires[800]), .A1 (CLOCK_slo__n2241), .A2 (n_0_21));
NOR2_X1 i_0_435 (.ZN (normalizedWires[799]), .A1 (n_0_43), .A2 (n_0_20));
BUF_X2 slo___L1_c794 (.Z (slo___n867), .A (n_0_49));
NOR2_X1 i_0_433 (.ZN (normalizedWires[797]), .A1 (n_0_43), .A2 (slo___n436));
NOR2_X1 i_0_432 (.ZN (normalizedWires[796]), .A1 (n_0_43), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_431 (.ZN (normalizedWires[795]), .A1 (CLOCK_slo__n2241), .A2 (n_0_16));
NOR2_X1 i_0_430 (.ZN (normalizedWires[794]), .A1 (n_0_43), .A2 (n_0_15));
NOR2_X1 i_0_429 (.ZN (normalizedWires[793]), .A1 (CLOCK_slo__n2241), .A2 (n_0_14));
NOR2_X1 i_0_428 (.ZN (normalizedWires[792]), .A1 (n_0_43), .A2 (n_0_13));
NOR2_X1 i_0_427 (.ZN (normalizedWires[791]), .A1 (CLOCK_slo__n2241), .A2 (n_0_12));
NOR2_X1 i_0_426 (.ZN (normalizedWires[790]), .A1 (n_0_43), .A2 (n_0_11));
NOR2_X1 i_0_425 (.ZN (normalizedWires[789]), .A1 (n_0_43), .A2 (n_0_10));
NOR2_X1 i_0_424 (.ZN (normalizedWires[788]), .A1 (n_0_43), .A2 (n_0_9));
NOR2_X1 i_0_423 (.ZN (normalizedWires[787]), .A1 (n_0_43), .A2 (n_0_76));
NOR2_X1 i_0_422 (.ZN (normalizedWires[786]), .A1 (n_0_43), .A2 (n_0_67));
NOR2_X1 i_0_421 (.ZN (normalizedWires[785]), .A1 (n_0_43), .A2 (sgo__n175));
NOR2_X1 i_0_420 (.ZN (normalizedWires[784]), .A1 (n_0_43), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_419 (.ZN (normalizedWires[783]), .A1 (n_0_43), .A2 (n_0_4));
NOR2_X1 i_0_418 (.ZN (normalizedWires[782]), .A1 (n_0_43), .A2 (n_0_3));
NOR2_X1 i_0_417 (.ZN (normalizedWires[781]), .A1 (n_0_43), .A2 (n_0_2));
NOR2_X1 i_0_416 (.ZN (normalizedWires[780]), .A1 (n_0_43), .A2 (n_0_73));
INV_X8 i_0_415 (.ZN (n_0_43), .A (B[12]));
NOR2_X1 i_0_414 (.ZN (normalizedWires[745]), .A1 (n_0_42), .A2 (slo__n785));
NOR2_X1 i_0_413 (.ZN (normalizedWires[744]), .A1 (n_0_42), .A2 (slo__n332));
NOR2_X1 i_0_412 (.ZN (normalizedWires[743]), .A1 (n_0_42), .A2 (sgo__n131));
NOR2_X1 i_0_411 (.ZN (normalizedWires[742]), .A1 (n_0_42), .A2 (opt_ipo_n1675));
NOR2_X1 i_0_410 (.ZN (normalizedWires[741]), .A1 (n_0_42), .A2 (n_0_27));
NOR2_X1 i_0_409 (.ZN (normalizedWires[740]), .A1 (n_0_42), .A2 (n_0_26));
NOR2_X1 i_0_408 (.ZN (normalizedWires[739]), .A1 (n_0_42), .A2 (opt_ipo_n1677));
NOR2_X1 i_0_407 (.ZN (normalizedWires[738]), .A1 (n_0_42), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_406 (.ZN (normalizedWires[737]), .A1 (n_0_42), .A2 (n_0_23));
NOR2_X1 i_0_405 (.ZN (normalizedWires[736]), .A1 (n_0_42), .A2 (n_0_22));
NOR2_X1 i_0_404 (.ZN (normalizedWires[735]), .A1 (n_0_42), .A2 (n_0_21));
NOR2_X1 i_0_403 (.ZN (normalizedWires[734]), .A1 (n_0_42), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_402 (.ZN (normalizedWires[733]), .A1 (n_0_42), .A2 (n_0_19));
NOR2_X1 i_0_401 (.ZN (normalizedWires[732]), .A1 (n_0_42), .A2 (slo__n298));
NOR2_X1 i_0_400 (.ZN (normalizedWires[731]), .A1 (n_0_42), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_399 (.ZN (normalizedWires[730]), .A1 (n_0_42), .A2 (n_0_16));
NOR2_X1 i_0_398 (.ZN (normalizedWires[729]), .A1 (n_0_42), .A2 (n_0_15));
NOR2_X1 i_0_397 (.ZN (normalizedWires[728]), .A1 (n_0_42), .A2 (n_0_14));
NOR2_X1 i_0_396 (.ZN (normalizedWires[727]), .A1 (n_0_42), .A2 (n_0_13));
NOR2_X1 i_0_395 (.ZN (normalizedWires[726]), .A1 (n_0_42), .A2 (opt_ipo_n1525));
NOR2_X1 i_0_394 (.ZN (normalizedWires[725]), .A1 (n_0_42), .A2 (n_0_11));
NOR2_X1 i_0_393 (.ZN (normalizedWires[724]), .A1 (n_0_42), .A2 (opt_ipo_n1556));
NOR2_X1 i_0_392 (.ZN (normalizedWires[723]), .A1 (n_0_42), .A2 (n_0_9));
NOR2_X1 i_0_391 (.ZN (normalizedWires[722]), .A1 (n_0_42), .A2 (slo__n1013));
NOR2_X1 i_0_390 (.ZN (normalizedWires[721]), .A1 (n_0_42), .A2 (n_0_67));
NOR2_X2 i_0_389 (.ZN (normalizedWires[720]), .A1 (n_0_42), .A2 (sgo__n175));
NOR2_X1 i_0_388 (.ZN (normalizedWires[719]), .A1 (n_0_42), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_387 (.ZN (normalizedWires[718]), .A1 (n_0_42), .A2 (n_0_4));
NOR2_X1 i_0_386 (.ZN (normalizedWires[717]), .A1 (n_0_42), .A2 (n_0_3));
NOR2_X1 i_0_385 (.ZN (normalizedWires[716]), .A1 (n_0_42), .A2 (n_0_2));
NOR2_X1 i_0_384 (.ZN (normalizedWires[715]), .A1 (n_0_42), .A2 (n_0_73));
INV_X8 i_0_383 (.ZN (n_0_42), .A (B[11]));
NOR2_X1 i_0_382 (.ZN (normalizedWires[680]), .A1 (opt_ipo_n1647), .A2 (slo__n785));
NOR2_X1 i_0_381 (.ZN (normalizedWires[679]), .A1 (n_0_30), .A2 (opt_ipo_n1649));
NOR2_X2 i_0_380 (.ZN (normalizedWires[678]), .A1 (slo__n1036), .A2 (n_0_29));
BUF_X4 opt_ipo_c1385 (.Z (opt_ipo_n1525), .A (n_0_12));
NOR2_X2 i_0_378 (.ZN (normalizedWires[676]), .A1 (opt_ipo_n1649), .A2 (n_0_27));
NOR2_X1 slo__sro_c693 (.ZN (normalizedWires[804]), .A1 (n_0_43), .A2 (slo__n1158));
NOR2_X1 i_0_376 (.ZN (normalizedWires[674]), .A1 (opt_ipo_n1649), .A2 (slo__n1158));
NOR2_X2 CLOCK_slo__sro_c2752 (.ZN (normalizedWires[1258]), .A1 (n_0_50), .A2 (opt_ipo_n1532));
NOR2_X2 i_0_374 (.ZN (normalizedWires[672]), .A1 (opt_ipo_n1649), .A2 (slo__n616));
NOR2_X1 i_0_373 (.ZN (normalizedWires[671]), .A1 (n_0_22), .A2 (opt_ipo_n1649));
NOR2_X4 i_0_372 (.ZN (normalizedWires[670]), .A1 (opt_ipo_n1649), .A2 (n_0_21));
NOR2_X1 i_0_371 (.ZN (normalizedWires[669]), .A1 (opt_ipo_n1649), .A2 (n_0_20));
NOR2_X1 i_0_370 (.ZN (normalizedWires[668]), .A1 (opt_ipo_n1649), .A2 (n_0_19));
NOR2_X1 i_0_369 (.ZN (normalizedWires[667]), .A1 (opt_ipo_n1649), .A2 (slo__n381));
NOR2_X2 CLOCK_slo__sro_c2915 (.ZN (normalizedWires[1182]), .A1 (n_0_49), .A2 (n_0_13));
NOR2_X1 CLOCK_slo__mro_c1983 (.ZN (normalizedWires[268]), .A1 (slo__n907), .A2 (n_0_35));
NOR2_X1 i_0_366 (.ZN (normalizedWires[664]), .A1 (slo__n1036), .A2 (n_0_15));
NOR2_X2 i_0_365 (.ZN (normalizedWires[663]), .A1 (opt_ipo_n1649), .A2 (n_0_14));
NOR2_X1 i_0_364 (.ZN (normalizedWires[662]), .A1 (opt_ipo_n1649), .A2 (slo__n1127));
NOR2_X1 slo__sro_c688 (.ZN (normalizedWires[675]), .A1 (n_0_26), .A2 (opt_ipo_n1649));
NOR2_X1 i_0_362 (.ZN (normalizedWires[660]), .A1 (opt_ipo_n1649), .A2 (n_0_11));
NOR2_X1 i_0_361 (.ZN (normalizedWires[659]), .A1 (opt_ipo_n1649), .A2 (n_0_10));
NOR2_X1 i_0_360 (.ZN (normalizedWires[658]), .A1 (opt_ipo_n1649), .A2 (n_0_9));
NOR2_X2 i_0_359 (.ZN (normalizedWires[657]), .A1 (CLOCK_slo__n2250), .A2 (n_0_76));
NOR2_X2 i_0_358 (.ZN (normalizedWires[656]), .A1 (CLOCK_slo__n2250), .A2 (n_0_67));
NOR2_X2 i_0_357 (.ZN (normalizedWires[655]), .A1 (opt_ipo_n1649), .A2 (n_0_68));
NOR2_X2 i_0_356 (.ZN (normalizedWires[654]), .A1 (opt_ipo_n1649), .A2 (n_0_5));
NOR2_X1 i_0_352 (.ZN (normalizedWires[650]), .A1 (slo__n1036), .A2 (n_0_73));
NOR2_X1 i_0_350 (.ZN (normalizedWires[615]), .A1 (n_0_40), .A2 (n_0_31));
NOR2_X2 i_0_349 (.ZN (normalizedWires[614]), .A1 (n_0_40), .A2 (n_0_30));
NOR2_X2 i_0_348 (.ZN (normalizedWires[613]), .A1 (n_0_40), .A2 (n_0_29));
NOR2_X1 i_0_347 (.ZN (normalizedWires[612]), .A1 (n_0_40), .A2 (n_0_28));
NOR2_X1 i_0_346 (.ZN (normalizedWires[611]), .A1 (n_0_27), .A2 (n_0_40));
NOR2_X2 CLOCK_slo__mro_c2603 (.ZN (normalizedWires[285]), .A1 (n_0_26), .A2 (n_0_35));
NOR2_X1 i_0_344 (.ZN (normalizedWires[609]), .A1 (n_0_40), .A2 (slo__n1158));
NOR2_X1 i_0_343 (.ZN (normalizedWires[608]), .A1 (n_0_40), .A2 (opt_ipo_n1532));
NOR2_X2 i_0_342 (.ZN (normalizedWires[607]), .A1 (n_0_40), .A2 (slo__n616));
NOR2_X1 i_0_341 (.ZN (normalizedWires[606]), .A1 (n_0_40), .A2 (n_0_22));
NOR2_X1 i_0_340 (.ZN (normalizedWires[605]), .A1 (n_0_40), .A2 (n_0_21));
NOR2_X1 i_0_339 (.ZN (normalizedWires[604]), .A1 (n_0_40), .A2 (n_0_20));
NOR2_X1 i_0_338 (.ZN (normalizedWires[603]), .A1 (n_0_40), .A2 (n_0_19));
NOR2_X2 i_0_337 (.ZN (normalizedWires[602]), .A1 (n_0_40), .A2 (slo___n436));
NOR2_X1 i_0_336 (.ZN (normalizedWires[601]), .A1 (n_0_40), .A2 (n_0_17));
NOR2_X1 i_0_335 (.ZN (normalizedWires[600]), .A1 (n_0_40), .A2 (n_0_16));
NOR2_X1 i_0_334 (.ZN (normalizedWires[599]), .A1 (n_0_40), .A2 (n_0_15));
NOR2_X1 i_0_333 (.ZN (normalizedWires[598]), .A1 (n_0_14), .A2 (n_0_40));
NOR2_X1 i_0_332 (.ZN (normalizedWires[597]), .A1 (n_0_40), .A2 (n_0_13));
NOR2_X1 i_0_331 (.ZN (normalizedWires[596]), .A1 (n_0_12), .A2 (n_0_40));
NOR2_X1 i_0_330 (.ZN (normalizedWires[595]), .A1 (n_0_40), .A2 (n_0_11));
NOR2_X1 i_0_329 (.ZN (normalizedWires[594]), .A1 (n_0_40), .A2 (n_0_10));
NOR2_X2 i_0_328 (.ZN (normalizedWires[593]), .A1 (n_0_40), .A2 (n_0_9));
NOR2_X4 i_0_327 (.ZN (normalizedWires[592]), .A1 (n_0_40), .A2 (n_0_76));
BUF_X8 opt_ipo_c1531 (.Z (opt_ipo_n1677), .A (n_0_25));
NOR2_X1 i_0_325 (.ZN (normalizedWires[590]), .A1 (n_0_40), .A2 (n_0_68));
NOR2_X1 i_0_322 (.ZN (normalizedWires[587]), .A1 (n_0_40), .A2 (n_0_3));
NOR2_X1 i_0_321 (.ZN (normalizedWires[586]), .A1 (n_0_40), .A2 (n_0_2));
NOR2_X1 i_0_320 (.ZN (normalizedWires[585]), .A1 (n_0_40), .A2 (n_0_73));
NOR2_X1 i_0_318 (.ZN (normalizedWires[550]), .A1 (n_0_39), .A2 (slo__n785));
NOR2_X1 i_0_317 (.ZN (normalizedWires[549]), .A1 (n_0_39), .A2 (slo__n332));
NOR2_X1 i_0_316 (.ZN (normalizedWires[548]), .A1 (n_0_39), .A2 (sgo__n131));
NOR2_X1 i_0_315 (.ZN (normalizedWires[547]), .A1 (n_0_39), .A2 (opt_ipo_n1675));
NOR2_X1 i_0_314 (.ZN (normalizedWires[546]), .A1 (n_0_39), .A2 (n_0_27));
NOR2_X1 i_0_313 (.ZN (normalizedWires[545]), .A1 (n_0_39), .A2 (n_0_26));
NOR2_X1 i_0_312 (.ZN (normalizedWires[544]), .A1 (n_0_39), .A2 (opt_ipo_n1677));
NOR2_X1 i_0_311 (.ZN (normalizedWires[543]), .A1 (n_0_39), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_310 (.ZN (normalizedWires[542]), .A1 (n_0_39), .A2 (sgo__n110));
NOR2_X1 i_0_309 (.ZN (normalizedWires[541]), .A1 (n_0_39), .A2 (slo__n302));
NOR2_X1 i_0_308 (.ZN (normalizedWires[540]), .A1 (n_0_39), .A2 (n_0_21));
NOR2_X1 i_0_307 (.ZN (normalizedWires[539]), .A1 (n_0_39), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_306 (.ZN (normalizedWires[538]), .A1 (n_0_39), .A2 (n_0_19));
NOR2_X1 i_0_305 (.ZN (normalizedWires[537]), .A1 (n_0_39), .A2 (slo__n298));
NOR2_X1 i_0_304 (.ZN (normalizedWires[536]), .A1 (n_0_39), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_303 (.ZN (normalizedWires[535]), .A1 (n_0_39), .A2 (n_0_16));
NOR2_X1 i_0_302 (.ZN (normalizedWires[534]), .A1 (n_0_39), .A2 (n_0_15));
NOR2_X1 i_0_301 (.ZN (normalizedWires[533]), .A1 (n_0_39), .A2 (n_0_14));
NOR2_X1 i_0_300 (.ZN (normalizedWires[532]), .A1 (n_0_39), .A2 (CLOCK_sgo__n1896));
NOR2_X1 i_0_299 (.ZN (normalizedWires[531]), .A1 (n_0_39), .A2 (opt_ipo_n1525));
NOR2_X1 i_0_298 (.ZN (normalizedWires[530]), .A1 (n_0_39), .A2 (n_0_11));
NOR2_X1 i_0_297 (.ZN (normalizedWires[529]), .A1 (n_0_39), .A2 (slo__n1191));
NOR2_X1 i_0_296 (.ZN (normalizedWires[528]), .A1 (n_0_39), .A2 (n_0_9));
NOR2_X1 i_0_295 (.ZN (normalizedWires[527]), .A1 (n_0_39), .A2 (n_0_76));
NOR2_X1 i_0_294 (.ZN (normalizedWires[526]), .A1 (n_0_39), .A2 (n_0_67));
NOR2_X1 i_0_293 (.ZN (normalizedWires[525]), .A1 (n_0_39), .A2 (sgo__n175));
NOR2_X1 i_0_292 (.ZN (normalizedWires[524]), .A1 (n_0_39), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_291 (.ZN (normalizedWires[523]), .A1 (n_0_39), .A2 (n_0_4));
NOR2_X1 i_0_290 (.ZN (normalizedWires[522]), .A1 (n_0_39), .A2 (n_0_3));
NOR2_X4 i_0_289 (.ZN (normalizedWires[521]), .A1 (n_0_39), .A2 (n_0_2));
NOR2_X1 i_0_288 (.ZN (normalizedWires[520]), .A1 (n_0_39), .A2 (n_0_73));
INV_X4 i_0_287 (.ZN (n_0_39), .A (B[8]));
NOR2_X1 i_0_286 (.ZN (normalizedWires[485]), .A1 (n_0_38), .A2 (slo__n785));
NOR2_X1 i_0_285 (.ZN (normalizedWires[484]), .A1 (n_0_38), .A2 (slo__n332));
NOR2_X1 i_0_284 (.ZN (normalizedWires[483]), .A1 (n_0_38), .A2 (n_0_29));
NOR2_X2 i_0_283 (.ZN (normalizedWires[482]), .A1 (n_0_38), .A2 (n_0_28));
NOR2_X2 i_0_282 (.ZN (normalizedWires[481]), .A1 (n_0_38), .A2 (n_0_27));
NOR2_X1 i_0_281 (.ZN (normalizedWires[480]), .A1 (n_0_38), .A2 (n_0_26));
NOR2_X1 i_0_280 (.ZN (normalizedWires[479]), .A1 (n_0_38), .A2 (n_0_25));
NOR2_X1 i_0_279 (.ZN (normalizedWires[478]), .A1 (n_0_38), .A2 (opt_ipo_n1532));
NOR2_X2 i_0_278 (.ZN (normalizedWires[477]), .A1 (slo__n616), .A2 (n_0_38));
NOR2_X1 i_0_277 (.ZN (normalizedWires[476]), .A1 (n_0_38), .A2 (n_0_22));
NOR2_X1 i_0_276 (.ZN (normalizedWires[475]), .A1 (n_0_38), .A2 (n_0_21));
NOR2_X1 i_0_275 (.ZN (normalizedWires[474]), .A1 (n_0_38), .A2 (n_0_20));
NOR2_X1 i_0_274 (.ZN (normalizedWires[473]), .A1 (n_0_38), .A2 (n_0_19));
NOR2_X1 i_0_273 (.ZN (normalizedWires[472]), .A1 (n_0_38), .A2 (n_0_18));
NOR2_X1 i_0_272 (.ZN (normalizedWires[471]), .A1 (n_0_38), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_271 (.ZN (normalizedWires[470]), .A1 (n_0_38), .A2 (n_0_16));
NOR2_X1 i_0_270 (.ZN (normalizedWires[469]), .A1 (n_0_38), .A2 (n_0_15));
NOR2_X1 i_0_269 (.ZN (normalizedWires[468]), .A1 (n_0_38), .A2 (n_0_14));
NOR2_X1 i_0_268 (.ZN (normalizedWires[467]), .A1 (n_0_38), .A2 (n_0_13));
NOR2_X1 i_0_267 (.ZN (normalizedWires[466]), .A1 (n_0_12), .A2 (n_0_38));
NOR2_X4 i_0_266 (.ZN (normalizedWires[465]), .A1 (n_0_38), .A2 (n_0_11));
BUF_X1 slo___L1_c1110 (.Z (slo___n1215), .A (opt_ipo_n1532));
NOR2_X2 i_0_264 (.ZN (normalizedWires[463]), .A1 (n_0_38), .A2 (slo__n907));
NOR2_X2 i_0_263 (.ZN (normalizedWires[462]), .A1 (n_0_38), .A2 (n_0_76));
NOR2_X2 i_0_262 (.ZN (normalizedWires[461]), .A1 (n_0_38), .A2 (n_0_67));
NOR2_X1 i_0_261 (.ZN (normalizedWires[460]), .A1 (n_0_38), .A2 (sgo__n175));
NOR2_X1 i_0_260 (.ZN (normalizedWires[459]), .A1 (n_0_38), .A2 (n_0_5));
NOR2_X2 i_0_258 (.ZN (normalizedWires[457]), .A1 (n_0_38), .A2 (n_0_3));
NOR2_X1 i_0_257 (.ZN (normalizedWires[456]), .A1 (n_0_38), .A2 (n_0_2));
NOR2_X1 i_0_256 (.ZN (normalizedWires[455]), .A1 (n_0_38), .A2 (n_0_73));
NOR2_X1 i_0_254 (.ZN (normalizedWires[420]), .A1 (spw__n3569), .A2 (slo__n785));
NOR2_X1 i_0_253 (.ZN (normalizedWires[419]), .A1 (n_0_30), .A2 (spw__n3569));
NOR2_X1 i_0_252 (.ZN (normalizedWires[418]), .A1 (spw__n3569), .A2 (n_0_29));
NOR2_X2 i_0_251 (.ZN (normalizedWires[417]), .A1 (spw__n3570), .A2 (n_0_28));
NOR2_X1 i_0_250 (.ZN (normalizedWires[416]), .A1 (spw__n3569), .A2 (n_0_27));
NOR2_X2 i_0_249 (.ZN (normalizedWires[415]), .A1 (spw__n3571), .A2 (n_0_26));
NOR2_X1 i_0_248 (.ZN (normalizedWires[414]), .A1 (spw__n3569), .A2 (n_0_25));
NOR2_X1 i_0_247 (.ZN (normalizedWires[413]), .A1 (spw__n3569), .A2 (opt_ipo_n1532));
NOR2_X2 i_0_246 (.ZN (normalizedWires[412]), .A1 (spw__n3573), .A2 (n_0_23));
NOR2_X1 i_0_245 (.ZN (normalizedWires[411]), .A1 (spw__n3572), .A2 (n_0_22));
NOR2_X1 i_0_244 (.ZN (normalizedWires[410]), .A1 (spw__n3569), .A2 (n_0_21));
NOR2_X1 i_0_243 (.ZN (normalizedWires[409]), .A1 (spw__n3569), .A2 (n_0_20));
NOR2_X1 i_0_242 (.ZN (normalizedWires[408]), .A1 (spw__n3569), .A2 (n_0_19));
NOR2_X1 i_0_241 (.ZN (normalizedWires[407]), .A1 (spw__n3569), .A2 (n_0_18));
NOR2_X1 i_0_240 (.ZN (normalizedWires[406]), .A1 (spw__n3569), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_239 (.ZN (normalizedWires[405]), .A1 (spw__n3569), .A2 (n_0_16));
NOR2_X1 i_0_238 (.ZN (normalizedWires[404]), .A1 (spw__n3569), .A2 (n_0_15));
NOR2_X1 i_0_237 (.ZN (normalizedWires[403]), .A1 (spw__n3569), .A2 (n_0_14));
NOR2_X1 i_0_236 (.ZN (normalizedWires[402]), .A1 (spw__n3574), .A2 (n_0_13));
NOR2_X4 i_0_235 (.ZN (normalizedWires[401]), .A1 (spw__n3575), .A2 (n_0_12));
NOR2_X2 CLOCK_slo__sro_c2877 (.ZN (normalizedWires[666]), .A1 (opt_ipo_n1550), .A2 (opt_ipo_n1649));
NOR2_X2 i_0_233 (.ZN (normalizedWires[399]), .A1 (spw__n3574), .A2 (n_0_10));
NOR2_X1 i_0_232 (.ZN (normalizedWires[398]), .A1 (spw__n3574), .A2 (slo__n907));
NOR2_X2 i_0_231 (.ZN (normalizedWires[397]), .A1 (spw__n3574), .A2 (n_0_76));
NOR2_X1 i_0_230 (.ZN (normalizedWires[396]), .A1 (spw__n3574), .A2 (n_0_67));
NOR2_X1 i_0_226 (.ZN (normalizedWires[392]), .A1 (spw__n3574), .A2 (n_0_3));
NOR2_X1 i_0_225 (.ZN (normalizedWires[391]), .A1 (spw__n3574), .A2 (n_0_2));
NOR2_X1 i_0_224 (.ZN (normalizedWires[390]), .A1 (spw__n3574), .A2 (n_0_73));
NOR2_X1 i_0_222 (.ZN (normalizedWires[355]), .A1 (n_0_36), .A2 (slo__n785));
NOR2_X1 i_0_221 (.ZN (normalizedWires[354]), .A1 (n_0_36), .A2 (slo__n332));
NOR2_X1 i_0_220 (.ZN (normalizedWires[353]), .A1 (n_0_36), .A2 (n_0_29));
NOR2_X1 i_0_219 (.ZN (normalizedWires[352]), .A1 (n_0_36), .A2 (opt_ipo_n1675));
NOR2_X1 i_0_218 (.ZN (normalizedWires[351]), .A1 (n_0_36), .A2 (sgo__n168));
NOR2_X1 i_0_217 (.ZN (normalizedWires[350]), .A1 (n_0_36), .A2 (sgo__n27));
NOR2_X1 i_0_216 (.ZN (normalizedWires[349]), .A1 (n_0_36), .A2 (opt_ipo_n1677));
NOR2_X1 i_0_215 (.ZN (normalizedWires[348]), .A1 (n_0_36), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_214 (.ZN (normalizedWires[347]), .A1 (n_0_36), .A2 (sgo__n110));
NOR2_X1 i_0_213 (.ZN (normalizedWires[346]), .A1 (n_0_36), .A2 (slo__n302));
NOR2_X1 i_0_212 (.ZN (normalizedWires[345]), .A1 (n_0_36), .A2 (n_0_21));
NOR2_X1 i_0_211 (.ZN (normalizedWires[344]), .A1 (n_0_36), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_210 (.ZN (normalizedWires[343]), .A1 (n_0_36), .A2 (n_0_19));
NOR2_X1 i_0_209 (.ZN (normalizedWires[342]), .A1 (n_0_36), .A2 (slo__n298));
NOR2_X1 i_0_208 (.ZN (normalizedWires[341]), .A1 (n_0_36), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_207 (.ZN (normalizedWires[340]), .A1 (n_0_36), .A2 (n_0_16));
NOR2_X2 i_0_206 (.ZN (normalizedWires[339]), .A1 (n_0_36), .A2 (CLOCK_sgo__n1891));
NOR2_X1 i_0_205 (.ZN (normalizedWires[338]), .A1 (n_0_36), .A2 (n_0_14));
NOR2_X1 i_0_204 (.ZN (normalizedWires[337]), .A1 (n_0_36), .A2 (CLOCK_sgo__n1896));
NOR2_X1 i_0_203 (.ZN (normalizedWires[336]), .A1 (n_0_36), .A2 (CLOCK_slo__n2695));
NOR2_X1 i_0_202 (.ZN (normalizedWires[335]), .A1 (n_0_36), .A2 (n_0_11));
NOR2_X1 i_0_201 (.ZN (normalizedWires[334]), .A1 (n_0_36), .A2 (opt_ipo_n1556));
NOR2_X1 i_0_200 (.ZN (normalizedWires[333]), .A1 (n_0_36), .A2 (n_0_9));
NOR2_X1 i_0_199 (.ZN (normalizedWires[332]), .A1 (n_0_36), .A2 (n_0_76));
NOR2_X1 i_0_198 (.ZN (normalizedWires[331]), .A1 (n_0_36), .A2 (n_0_67));
NOR2_X1 i_0_197 (.ZN (normalizedWires[330]), .A1 (n_0_36), .A2 (sgo__n175));
NOR2_X1 i_0_196 (.ZN (normalizedWires[329]), .A1 (n_0_36), .A2 (opt_ipo_n1710));
NOR2_X1 i_0_195 (.ZN (normalizedWires[328]), .A1 (n_0_36), .A2 (n_0_4));
NOR2_X1 i_0_194 (.ZN (normalizedWires[327]), .A1 (n_0_36), .A2 (n_0_3));
NOR2_X1 i_0_193 (.ZN (normalizedWires[326]), .A1 (n_0_36), .A2 (n_0_2));
NOR2_X1 i_0_192 (.ZN (normalizedWires[325]), .A1 (n_0_36), .A2 (n_0_73));
INV_X4 i_0_191 (.ZN (n_0_36), .A (B[5]));
NOR2_X1 i_0_190 (.ZN (normalizedWires[290]), .A1 (n_0_35), .A2 (n_0_31));
NOR2_X1 i_0_189 (.ZN (normalizedWires[289]), .A1 (n_0_35), .A2 (n_0_30));
NOR2_X1 i_0_188 (.ZN (normalizedWires[288]), .A1 (n_0_35), .A2 (n_0_29));
NOR2_X1 i_0_187 (.ZN (normalizedWires[287]), .A1 (n_0_35), .A2 (n_0_28));
NOR2_X2 i_0_186 (.ZN (normalizedWires[286]), .A1 (n_0_35), .A2 (n_0_27));
NOR2_X4 CLOCK_slo__mro_c2627 (.ZN (normalizedWires[1645]), .A1 (n_0_56), .A2 (n_0_21));
NOR2_X1 i_0_184 (.ZN (normalizedWires[284]), .A1 (n_0_35), .A2 (n_0_25));
NOR2_X1 i_0_183 (.ZN (normalizedWires[283]), .A1 (n_0_35), .A2 (opt_ipo_n1532));
INV_X4 CLOCK_slo__c2678 (.ZN (CLOCK_slo__n2927), .A (n_0_68));
NOR2_X1 i_0_181 (.ZN (normalizedWires[281]), .A1 (n_0_35), .A2 (n_0_22));
NOR2_X1 i_0_180 (.ZN (normalizedWires[280]), .A1 (n_0_35), .A2 (n_0_21));
NOR2_X1 i_0_179 (.ZN (normalizedWires[279]), .A1 (n_0_35), .A2 (n_0_20));
NOR2_X1 i_0_178 (.ZN (normalizedWires[278]), .A1 (n_0_35), .A2 (n_0_19));
NOR2_X1 i_0_177 (.ZN (normalizedWires[277]), .A1 (n_0_35), .A2 (n_0_18));
NOR2_X1 i_0_176 (.ZN (normalizedWires[276]), .A1 (n_0_35), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_175 (.ZN (normalizedWires[275]), .A1 (n_0_35), .A2 (n_0_16));
NOR2_X1 i_0_174 (.ZN (normalizedWires[274]), .A1 (n_0_35), .A2 (n_0_15));
NOR2_X4 i_0_173 (.ZN (normalizedWires[273]), .A1 (n_0_35), .A2 (n_0_14));
NOR2_X2 i_0_172 (.ZN (normalizedWires[272]), .A1 (n_0_35), .A2 (CLOCK_slo__n3242));
BUF_X8 slo__c344 (.Z (slo__n298), .A (slo__n317));
NOR2_X1 i_0_170 (.ZN (normalizedWires[270]), .A1 (n_0_35), .A2 (slo__n1353));
NOR2_X1 i_0_169 (.ZN (normalizedWires[269]), .A1 (n_0_35), .A2 (slo__n791));
NOR2_X2 slo__sro_c858 (.ZN (normalizedWires[1064]), .A1 (n_0_25), .A2 (n_0_47));
NOR2_X1 i_0_165 (.ZN (normalizedWires[265]), .A1 (n_0_35), .A2 (sgo__n175));
BUF_X2 spw__L1_c3185 (.Z (spw__n3533), .A (opt_ipo_n1675));
NOR2_X1 i_0_163 (.ZN (normalizedWires[263]), .A1 (n_0_35), .A2 (n_0_4));
NOR2_X1 i_0_162 (.ZN (normalizedWires[262]), .A1 (n_0_35), .A2 (n_0_3));
NOR2_X1 i_0_161 (.ZN (normalizedWires[261]), .A1 (n_0_35), .A2 (n_0_2));
NOR2_X1 i_0_160 (.ZN (normalizedWires[260]), .A1 (n_0_35), .A2 (n_0_73));
NOR2_X1 i_0_158 (.ZN (normalizedWires[225]), .A1 (n_0_34), .A2 (n_0_31));
NOR2_X2 i_0_157 (.ZN (normalizedWires[224]), .A1 (n_0_34), .A2 (n_0_30));
NOR2_X1 i_0_156 (.ZN (normalizedWires[223]), .A1 (n_0_34), .A2 (n_0_29));
NOR2_X1 i_0_155 (.ZN (normalizedWires[222]), .A1 (n_0_28), .A2 (n_0_34));
NOR2_X1 i_0_154 (.ZN (normalizedWires[221]), .A1 (n_0_34), .A2 (n_0_27));
NOR2_X1 i_0_153 (.ZN (normalizedWires[220]), .A1 (n_0_26), .A2 (n_0_34));
NOR2_X1 i_0_152 (.ZN (normalizedWires[219]), .A1 (n_0_34), .A2 (n_0_25));
NOR2_X1 i_0_151 (.ZN (normalizedWires[218]), .A1 (n_0_34), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_150 (.ZN (normalizedWires[217]), .A1 (n_0_34), .A2 (n_0_23));
NOR2_X1 i_0_148 (.ZN (normalizedWires[215]), .A1 (n_0_34), .A2 (n_0_21));
NOR2_X1 i_0_147 (.ZN (normalizedWires[214]), .A1 (n_0_34), .A2 (n_0_20));
NOR2_X1 i_0_146 (.ZN (normalizedWires[213]), .A1 (n_0_34), .A2 (n_0_19));
NOR2_X1 i_0_145 (.ZN (normalizedWires[212]), .A1 (n_0_34), .A2 (n_0_18));
NOR2_X1 i_0_144 (.ZN (normalizedWires[211]), .A1 (n_0_34), .A2 (opt_ipo_n1550));
NOR2_X1 i_0_143 (.ZN (normalizedWires[210]), .A1 (n_0_34), .A2 (n_0_16));
NOR2_X2 CLOCK_slo__mro_c1947 (.ZN (normalizedWires[665]), .A1 (n_0_16), .A2 (slo__n1036));
NOR2_X1 CLOCK_slo__sro_c2034 (.ZN (normalizedWires[1178]), .A1 (n_0_49), .A2 (n_0_9));
NOR2_X4 CLOCK_slo__sro_c2794 (.ZN (normalizedWires[5]), .A1 (n_0_68), .A2 (n_0_0));
NOR2_X4 i_0_139 (.ZN (normalizedWires[206]), .A1 (n_0_12), .A2 (n_0_34));
NOR2_X2 i_0_138 (.ZN (normalizedWires[205]), .A1 (n_0_34), .A2 (slo__n1353));
NOR2_X1 i_0_137 (.ZN (normalizedWires[204]), .A1 (slo__n791), .A2 (n_0_34));
NOR2_X1 i_0_136 (.ZN (normalizedWires[203]), .A1 (n_0_34), .A2 (n_0_9));
INV_X2 CLOCK_slo__c2093 (.ZN (CLOCK_slo__n2250), .A (B[10]));
NOR2_X1 i_0_132 (.ZN (normalizedWires[199]), .A1 (n_0_34), .A2 (n_0_5));
NOR2_X1 i_0_131 (.ZN (normalizedWires[198]), .A1 (n_0_34), .A2 (n_0_4));
NOR2_X1 i_0_130 (.ZN (normalizedWires[197]), .A1 (n_0_34), .A2 (n_0_3));
NOR2_X1 i_0_129 (.ZN (normalizedWires[196]), .A1 (n_0_34), .A2 (n_0_2));
NOR2_X1 i_0_128 (.ZN (normalizedWires[195]), .A1 (n_0_34), .A2 (n_0_73));
NOR2_X1 i_0_126 (.ZN (normalizedWires[160]), .A1 (n_0_33), .A2 (n_0_31));
NOR2_X1 i_0_125 (.ZN (normalizedWires[159]), .A1 (n_0_33), .A2 (n_0_30));
NOR2_X1 i_0_124 (.ZN (normalizedWires[158]), .A1 (n_0_33), .A2 (sgo__n131));
NOR2_X1 i_0_123 (.ZN (normalizedWires[157]), .A1 (n_0_33), .A2 (opt_ipo_n1675));
NOR2_X1 i_0_122 (.ZN (normalizedWires[156]), .A1 (n_0_33), .A2 (sgo__n168));
NOR2_X1 i_0_121 (.ZN (normalizedWires[155]), .A1 (n_0_33), .A2 (sgo__n27));
NOR2_X1 i_0_120 (.ZN (normalizedWires[154]), .A1 (n_0_33), .A2 (opt_ipo_n1677));
NOR2_X1 i_0_119 (.ZN (normalizedWires[153]), .A1 (n_0_33), .A2 (opt_ipo_n1532));
NOR2_X1 i_0_118 (.ZN (normalizedWires[152]), .A1 (n_0_33), .A2 (n_0_23));
NOR2_X1 i_0_117 (.ZN (normalizedWires[151]), .A1 (n_0_33), .A2 (slo__n302));
NOR2_X1 i_0_116 (.ZN (normalizedWires[150]), .A1 (n_0_33), .A2 (n_0_21));
NOR2_X1 i_0_115 (.ZN (normalizedWires[149]), .A1 (n_0_33), .A2 (opt_ipo_n1658));
NOR2_X1 i_0_114 (.ZN (normalizedWires[148]), .A1 (n_0_33), .A2 (n_0_19));
NOR2_X1 i_0_113 (.ZN (normalizedWires[147]), .A1 (n_0_33), .A2 (slo__n317));
NOR2_X1 i_0_112 (.ZN (normalizedWires[146]), .A1 (n_0_33), .A2 (opt_ipo_n1550));
CLKBUF_X1 CLOCK_slo___L3_c3_c2318 (.Z (CLOCK_slo_n2535), .A (CLOCK_slo___n2514));
NOR2_X2 i_0_110 (.ZN (normalizedWires[144]), .A1 (n_0_33), .A2 (n_0_15));
NOR2_X4 i_0_109 (.ZN (normalizedWires[143]), .A1 (n_0_33), .A2 (n_0_14));
NOR2_X2 i_0_108 (.ZN (normalizedWires[142]), .A1 (n_0_33), .A2 (slo__n1127));
NOR2_X2 i_0_107 (.ZN (normalizedWires[141]), .A1 (n_0_33), .A2 (n_0_12));
NOR2_X1 i_0_106 (.ZN (normalizedWires[140]), .A1 (n_0_33), .A2 (n_0_11));
NOR2_X1 i_0_105 (.ZN (normalizedWires[139]), .A1 (n_0_33), .A2 (n_0_10));
NOR2_X1 i_0_102 (.ZN (normalizedWires[136]), .A1 (n_0_33), .A2 (n_0_67));
NOR2_X1 i_0_101 (.ZN (normalizedWires[135]), .A1 (n_0_33), .A2 (n_0_68));
NOR2_X1 i_0_100 (.ZN (normalizedWires[134]), .A1 (n_0_33), .A2 (n_0_5));
NOR2_X1 i_0_99 (.ZN (normalizedWires[133]), .A1 (n_0_33), .A2 (n_0_4));
NOR2_X1 i_0_98 (.ZN (normalizedWires[132]), .A1 (n_0_33), .A2 (n_0_3));
NOR2_X1 i_0_97 (.ZN (normalizedWires[131]), .A1 (n_0_33), .A2 (n_0_2));
NOR2_X1 i_0_96 (.ZN (normalizedWires[130]), .A1 (n_0_33), .A2 (n_0_73));
NOR2_X1 i_0_94 (.ZN (normalizedWires[95]), .A1 (n_0_32), .A2 (n_0_31));
NOR2_X1 i_0_93 (.ZN (normalizedWires[94]), .A1 (n_0_32), .A2 (n_0_30));
NOR2_X1 i_0_92 (.ZN (normalizedWires[93]), .A1 (n_0_32), .A2 (sgo__n131));
NOR2_X1 i_0_91 (.ZN (normalizedWires[92]), .A1 (n_0_32), .A2 (opt_ipo_n1675));
NOR2_X1 i_0_90 (.ZN (normalizedWires[91]), .A1 (n_0_32), .A2 (n_0_27));
NOR2_X1 i_0_89 (.ZN (normalizedWires[90]), .A1 (n_0_32), .A2 (n_0_26));
NOR2_X1 i_0_88 (.ZN (normalizedWires[89]), .A1 (n_0_32), .A2 (n_0_25));
NOR2_X1 i_0_87 (.ZN (normalizedWires[88]), .A1 (n_0_32), .A2 (opt_ipo_n1532));
NOR2_X2 i_0_84 (.ZN (normalizedWires[85]), .A1 (n_0_32), .A2 (n_0_21));
NOR2_X4 i_0_83 (.ZN (normalizedWires[84]), .A1 (n_0_32), .A2 (n_0_20));
NOR2_X4 i_0_82 (.ZN (normalizedWires[83]), .A1 (n_0_32), .A2 (n_0_19));
NOR2_X4 i_0_80 (.ZN (normalizedWires[81]), .A1 (n_0_32), .A2 (n_0_17));
NOR2_X1 i_0_68 (.ZN (normalizedWires[69]), .A1 (n_0_32), .A2 (n_0_5));
NOR2_X4 i_0_67 (.ZN (normalizedWires[68]), .A1 (n_0_32), .A2 (n_0_4));
NOR2_X1 i_0_66 (.ZN (normalizedWires[67]), .A1 (n_0_32), .A2 (n_0_3));
NOR2_X1 i_0_65 (.ZN (normalizedWires[66]), .A1 (n_0_32), .A2 (n_0_2));
NOR2_X1 i_0_64 (.ZN (normalizedWires[65]), .A1 (n_0_32), .A2 (n_0_73));
NOR2_X1 i_0_62 (.ZN (normalizedWires[30]), .A1 (n_0_0), .A2 (n_0_31));
INV_X4 i_0_61 (.ZN (n_0_31), .A (A[30]));
NOR2_X1 i_0_60 (.ZN (normalizedWires[29]), .A1 (n_0_0), .A2 (slo__n332));
INV_X8 i_0_59 (.ZN (n_0_30), .A (A[29]));
NOR2_X1 i_0_58 (.ZN (normalizedWires[28]), .A1 (n_0_0), .A2 (sgo__n131));
INV_X8 i_0_57 (.ZN (n_0_29), .A (A[28]));
NOR2_X1 i_0_56 (.ZN (normalizedWires[27]), .A1 (n_0_0), .A2 (n_0_28));
NOR2_X2 i_0_54 (.ZN (normalizedWires[26]), .A1 (n_0_0), .A2 (n_0_27));
NOR2_X2 i_0_52 (.ZN (normalizedWires[25]), .A1 (n_0_0), .A2 (n_0_26));
NOR2_X2 CLOCK_slo__mro_c2555 (.ZN (normalizedWires[1247]), .A1 (n_0_50), .A2 (slo__n1127));
INV_X8 i_0_49 (.ZN (n_0_25), .A (A[24]));
NOR2_X2 i_0_48 (.ZN (normalizedWires[23]), .A1 (n_0_0), .A2 (opt_ipo_n1532));
NOR2_X2 CLOCK_slo__sro_c1996 (.ZN (normalizedWires[208]), .A1 (n_0_14), .A2 (n_0_34));
NOR2_X2 i_0_44 (.ZN (normalizedWires[21]), .A1 (n_0_0), .A2 (n_0_22));
NOR2_X2 i_0_40 (.ZN (normalizedWires[19]), .A1 (n_0_0), .A2 (n_0_20));
INV_X8 i_0_39 (.ZN (n_0_20), .A (A[19]));
NOR2_X4 i_0_36 (.ZN (normalizedWires[17]), .A1 (CLOCK_slo__n2403), .A2 (n_0_0));
BUF_X1 CLOCK_slo___L1_c2802 (.Z (CLOCK_slo___n3081), .A (n_0_4));
NOR2_X1 i_0_10 (.ZN (normalizedWires[4]), .A1 (n_0_0), .A2 (n_0_5));
NOR2_X1 i_0_8 (.ZN (normalizedWires[3]), .A1 (n_0_0), .A2 (CLOCK_slo___n3081));
NOR2_X1 i_0_6 (.ZN (normalizedWires[2]), .A1 (n_0_0), .A2 (n_0_3));
NOR2_X1 i_0_4 (.ZN (normalizedWires[1]), .A1 (n_0_0), .A2 (n_0_2));
NOR2_X1 i_0_2 (.ZN (normalizedWires[0]), .A1 (n_0_0), .A2 (n_0_73));
NOR2_X2 slo__mro_c309 (.ZN (normalizedWires[1644]), .A1 (n_0_20), .A2 (n_0_56));
INV_X1 CLOCK_slo___L2_c2_c2319 (.ZN (CLOCK_slo___n2514), .A (CLOCK_slo___n2515));
BUF_X4 slo__c348 (.Z (slo__n302), .A (n_0_22));
BUF_X4 slo__c378 (.Z (slo__n332), .A (n_0_30));
BUF_X2 slo__c363 (.Z (slo__n317), .A (CLOCK_slo__n2403));
NOR2_X2 slo__mro_c397 (.ZN (normalizedWires[677]), .A1 (n_0_28), .A2 (opt_ipo_n1649));
BUF_X2 slo__c424 (.Z (slo__n381), .A (CLOCK_slo__n2403));
NOR2_X2 slo__mro_c448 (.ZN (normalizedWires[986]), .A1 (n_0_12), .A2 (n_0_46));
BUF_X4 slo___L1_c471 (.Z (slo___n436), .A (CLOCK_slo__n2403));
INV_X2 CLOCK_slo__c2982 (.ZN (CLOCK_slo__n3319), .A (B[15]));
INV_X1 slo__c742 (.ZN (slo__n791), .A (A[9]));
NOR2_X2 slo__sro_c810 (.ZN (normalizedWires[1180]), .A1 (n_0_49), .A2 (n_0_11));
BUF_X2 slo__c524 (.Z (slo__n494), .A (B[19]));
NOR2_X1 slo__sro_c1055 (.ZN (normalizedWires[869]), .A1 (slo__n1158), .A2 (n_0_44));
INV_X4 slo__c604 (.ZN (slo__n616), .A (A[22]));
NOR2_X1 slo__sro_c627 (.ZN (normalizedWires[1834]), .A1 (n_0_64), .A2 (n_0_15));
NOR2_X1 slo__sro_c673 (.ZN (normalizedWires[1374]), .A1 (n_0_52), .A2 (n_0_10));
BUF_X4 slo__c733 (.Z (slo__n785), .A (n_0_31));
INV_X1 slo__c826 (.ZN (slo__n907), .A (A[8]));
INV_X2 slo__c923 (.ZN (slo__n1004), .A (B[15]));
BUF_X2 CLOCK_sgo__c1766 (.Z (CLOCK_sgo__n1896), .A (CLOCK_slo__n3242));
INV_X32 CLOCK_slo__c2680 (.ZN (sgo__n175), .A (CLOCK_slo__n2927));
BUF_X2 slo__c935 (.Z (slo__n1013), .A (n_0_76));
AND2_X2 slo__sro_c1049 (.ZN (normalizedWires[87]), .A1 (A[22]), .A2 (B[1]));
INV_X2 slo__c1041 (.ZN (slo__n1127), .A (A[12]));
INV_X4 slo__c1068 (.ZN (slo__n1158), .A (A[24]));
NOR2_X2 slo__sro_c1178 (.ZN (normalizedWires[1181]), .A1 (n_0_12), .A2 (n_0_49));
INV_X2 slo__c1220 (.ZN (slo__n1353), .A (A[10]));
NOR2_X1 CLOCK_slo__sro_c2120 (.ZN (normalizedWires[1041]), .A1 (n_0_47), .A2 (n_0_2));
BUF_X2 slo__c1195 (.Z (slo__n1306), .A (n_0_55));
INV_X2 CLOCK_slo__c2084 (.ZN (CLOCK_slo__n2241), .A (B[12]));
INV_X1 opt_ipo_c1504 (.ZN (opt_ipo_n1648), .A (opt_ipo_n1649));
NOR2_X4 CLOCK_slo__sro_c2252 (.ZN (normalizedWires[810]), .A1 (n_0_31), .A2 (n_0_43));
BUF_X4 opt_ipo_c1529 (.Z (opt_ipo_n1675), .A (n_0_28));
BUF_X16 opt_ipo_c1410 (.Z (opt_ipo_n1550), .A (n_0_17));
INV_X1 CLOCK_slo___L1_c1_c2320 (.ZN (CLOCK_slo___n2515), .A (B_4_PP_0));
NOR2_X1 CLOCK_slo__sro_c2341 (.ZN (normalizedWires[264]), .A1 (n_0_5), .A2 (CLOCK_slo__n2545));
BUF_X4 opt_ipo_c1416 (.Z (opt_ipo_n1556), .A (n_0_10));
BUF_X1 spw__L2_c3186 (.Z (spw__n3534), .A (spw__n3533));
BUF_X4 spw__L1_c3214 (.Z (spw__n3569), .A (spw__n3498));
BUF_X2 spw__L2_c3215 (.Z (spw__n3570), .A (spw__n3569));
INV_X1 CLOCK_slo__c2930 (.ZN (CLOCK_slo__n3242), .A (A[12]));
INV_X1 CLOCK_slo__c2338 (.ZN (CLOCK_slo__n2545), .A (B[4]));
BUF_X2 spw__L2_c3216 (.Z (spw__n3571), .A (spw__n3569));
BUF_X1 spw__L2_c3217 (.Z (spw__n3572), .A (spw__n3569));
BUF_X4 CLOCK_slo___L1_c2803 (.Z (CLOCK_slo___n3082), .A (n_0_4));
BUF_X4 opt_ipo_c1564 (.Z (opt_ipo_n1710), .A (n_0_5));
BUF_X2 spw__L2_c3218 (.Z (spw__n3573), .A (spw__n3569));
NOR2_X4 CLOCK_slo__sro_c2873 (.ZN (normalizedWires[400]), .A1 (n_0_11), .A2 (spw__n3574));
BUF_X8 spw__L1_c3219 (.Z (spw__n3574), .A (spw__n3498));
INV_X2 CLOCK_slo__c2820 (.ZN (CLOCK_slo__n3096), .A (A[25]));
BUF_X2 spw__L2_c3220 (.Z (spw__n3575), .A (spw__n3574));

endmodule //multiplyAllBits

module FA__4_247 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_247

module FA__4_243 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_243

module FA__4_239 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_239

module FA__4_235 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_235

module FA__4_231 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_231

module FA__4_227 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_227

module FA__4_223 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_223

module FA__4_219 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_219

module FA__4_215 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_215

module FA__4_211 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_211

module FA__4_207 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__sro_n10;
wire n_0_0;
wire CLOCK_slo__sro_n3;
wire CLOCK_slo__sro_n11;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n10), .B2 (CIN));
INV_X1 CLOCK_slo__sro_c7 (.ZN (CLOCK_slo__sro_n11), .A (B));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n3), .A (CIN));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (SUM), .A (CLOCK_slo__sro_n10), .B (CLOCK_slo__sro_n3));
XNOR2_X1 CLOCK_slo__sro_c8 (.ZN (CLOCK_slo__sro_n10), .A (A), .B (CLOCK_slo__sro_n11));

endmodule //FA__4_207

module FA__4_203 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n9;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X2 CLOCK_slo__mro_c6 (.ZN (CLOCK_slo__mro_n9), .A (A));
XNOR2_X2 CLOCK_slo__mro_c7 (.ZN (temp), .A (CLOCK_slo__mro_n9), .B (B));

endmodule //FA__4_203

module FA__4_199 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__mro_n10;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
INV_X1 CLOCK_slo__mro_c7 (.ZN (CLOCK_slo__mro_n10), .A (B));
INV_X1 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n3), .A (CIN));
XNOR2_X1 CLOCK_slo__mro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__mro_n3));
XNOR2_X2 CLOCK_slo__mro_c8 (.ZN (temp), .A (A), .B (CLOCK_slo__mro_n10));

endmodule //FA__4_199

module FA__4_195 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n1), .A (B));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (temp), .A (CLOCK_slo__sro_n1), .B (A));

endmodule //FA__4_195

module FA__4_191 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_191

module FA__4_187 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__sro_n27;
wire temp;
wire slo__sro_n9;
wire CLOCK_slo__sro_n28;


INV_X1 i_0_3 (.ZN (COUT), .A (CLOCK_slo__sro_n27));
AND2_X1 CLOCK_slo__sro_c14 (.ZN (CLOCK_slo__sro_n28), .A1 (A), .A2 (B));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n9), .A (CIN));
XNOR2_X2 slo__sro_c4 (.ZN (SUM), .A (temp), .B (slo__sro_n9));
AOI21_X1 CLOCK_slo__sro_c15 (.ZN (CLOCK_slo__sro_n27), .A (CLOCK_slo__sro_n28), .B1 (temp), .B2 (CIN));

endmodule //FA__4_187

module FA__4_183 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n4;
wire slo__mro_n8;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
INV_X1 slo__mro_c8 (.ZN (slo__mro_n8), .A (CIN));
INV_X1 slo__mro_c2 (.ZN (slo__mro_n4), .A (B));
XNOR2_X2 slo__mro_c3 (.ZN (temp), .A (slo__mro_n4), .B (A));
XNOR2_X2 slo__mro_c9 (.ZN (SUM), .A (temp), .B (slo__mro_n8));

endmodule //FA__4_183

module FA__4_179 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__mro_n22;
wire CLOCK_slo__mro_n23;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__mro_n22), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__mro_n22), .B (CIN));
INV_X2 CLOCK_slo__mro_c8 (.ZN (CLOCK_slo__mro_n23), .A (B));
XNOR2_X2 CLOCK_slo__mro_c9 (.ZN (CLOCK_slo__mro_n22), .A (CLOCK_slo__mro_n23), .B (A));

endmodule //FA__4_179

module FA__4_175 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_opt_ipo_n12;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (CLOCK_opt_ipo_n12), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (CLOCK_opt_ipo_n12));
INV_X2 CLOCK_opt_ipo_c8 (.ZN (CLOCK_opt_ipo_n12), .A (B));

endmodule //FA__4_175

module FA__4_171 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__mro_n37;
wire temp;
wire slo__sro_n10;
wire slo__sro_n11;
wire slo__sro_n18;


INV_X1 i_0_3 (.ZN (COUT), .A (slo__sro_n10));
INV_X1 slo__sro_c10 (.ZN (slo__sro_n18), .A (CIN));
INV_X2 CLOCK_slo__mro_c20 (.ZN (CLOCK_slo__mro_n37), .A (A));
AND2_X1 slo__sro_c4 (.ZN (slo__sro_n11), .A1 (B), .A2 (A));
AOI21_X2 slo__sro_c5 (.ZN (slo__sro_n10), .A (slo__sro_n11), .B1 (temp), .B2 (CIN));
XNOR2_X2 slo__sro_c11 (.ZN (SUM), .A (temp), .B (slo__sro_n18));
XNOR2_X2 CLOCK_slo__mro_c21 (.ZN (temp), .A (CLOCK_slo__mro_n37), .B (B));

endmodule //FA__4_171

module FA__4_167 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire CLOCK_slo__sro_n74;
wire CLOCK_slo__sro_n73;


INV_X2 i_0_3 (.ZN (COUT), .A (CLOCK_slo__sro_n73));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AOI21_X1 CLOCK_slo__sro_c46 (.ZN (CLOCK_slo__sro_n73), .A (CLOCK_slo__sro_n74), .B1 (temp), .B2 (CIN));
AND2_X1 CLOCK_slo__sro_c45 (.ZN (CLOCK_slo__sro_n74), .A1 (A), .A2 (B));

endmodule //FA__4_167

module FA__4_163 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo_n23;
wire n_0_0;
wire CLOCK_slo__sro_n26;
wire CLOCK_slo__sro_n27;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (CLOCK_slo_n23), .A2 (B), .B1 (CLOCK_slo__sro_n26), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n26), .B (CIN));
CLKBUF_X1 CLOCK_slo___L1_c1_c5 (.Z (CLOCK_slo_n23), .A (A));
INV_X1 CLOCK_slo__sro_c10 (.ZN (CLOCK_slo__sro_n27), .A (A));
XNOR2_X2 CLOCK_slo__sro_c11 (.ZN (CLOCK_slo__sro_n26), .A (CLOCK_slo__sro_n27), .B (B));

endmodule //FA__4_163

module FA__4_159 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire slo__mro_n10;
wire n_0_0;
wire slo__mro_n3;
wire slo__mro_n11;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__mro_n10), .B2 (CIN));
INV_X1 slo__mro_c7 (.ZN (slo__mro_n11), .A (B));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n3), .A (CIN));
XNOR2_X2 slo__mro_c2 (.ZN (SUM), .A (slo__mro_n10), .B (slo__mro_n3));
XNOR2_X2 slo__mro_c8 (.ZN (slo__mro_n10), .A (slo__mro_n11), .B (A));

endmodule //FA__4_159

module FA__4_155 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__mro_n9;
wire CLOCK_slo__mro_n10;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__mro_n9), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__mro_n9), .B (CIN));
INV_X2 CLOCK_slo__mro_c5 (.ZN (CLOCK_slo__mro_n10), .A (B));
XNOR2_X2 CLOCK_slo__mro_c6 (.ZN (CLOCK_slo__mro_n9), .A (CLOCK_slo__mro_n10), .B (A));

endmodule //FA__4_155

module FA__4_151 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n21;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 CLOCK_slo__sro_c10 (.Z (temp), .A (B), .B (A));
INV_X1 CLOCK_slo__mro_c4 (.ZN (CLOCK_slo__mro_n21), .A (CIN));
XNOR2_X1 CLOCK_slo__mro_c5 (.ZN (SUM), .A (temp), .B (CLOCK_slo__mro_n21));

endmodule //FA__4_151

module FA__4_147 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X4 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X2 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (CIN), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (B), .A2 (A));

endmodule //FA__4_147

module FA__4_143 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (SUM), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (CIN), .B1 (n_0_3), .B2 (n_0_0));
AND3_X2 i_0_5 (.ZN (n_0_4), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_0));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_1));
OAI21_X1 i_0_3 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (CIN));
NOR2_X2 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__4_143

module FA__4_139 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire opt_ipo_n13;


INV_X2 opt_ipo_c22 (.ZN (opt_ipo_n13), .A (B));
NAND2_X4 i_0_7 (.ZN (SUM), .A1 (n_0_4), .A2 (n_0_5));
OR3_X2 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_2), .A3 (CIN));
OAI21_X2 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_3), .B2 (n_0_2));
INV_X2 i_0_4 (.ZN (n_0_3), .A (n_0_1));
NOR2_X2 i_0_3 (.ZN (n_0_2), .A1 (opt_ipo_n13), .A2 (A));
NAND2_X2 i_0_2 (.ZN (n_0_1), .A1 (A), .A2 (opt_ipo_n13));
OAI21_X1 i_0_1 (.ZN (COUT), .A (n_0_1), .B1 (n_0_2), .B2 (n_0_0));
INV_X1 i_0_0 (.ZN (n_0_0), .A (CIN));

endmodule //FA__4_139

module FA__4_135 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (A));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (n_0_10), .A2 (B));
INV_X1 i_0_10 (.ZN (n_0_8), .A (B));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (A), .A2 (n_0_8));
NAND3_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_9), .A2 (CIN), .A3 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (CIN));
NOR2_X1 i_0_6 (.ZN (n_0_4), .A1 (A), .A2 (n_0_8));
INV_X1 i_0_5 (.ZN (n_0_3), .A (n_0_7));
OAI21_X2 i_0_4 (.ZN (n_0_2), .A (n_0_5), .B1 (n_0_3), .B2 (n_0_4));
NAND2_X2 i_0_3 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_6));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (A), .A2 (B));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
NOR2_X2 i_0_0 (.ZN (COUT), .A1 (n_0_0), .A2 (n_0_1));

endmodule //FA__4_135

module FA__4_131 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X2 i_0_7 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_6 (.ZN (n_0_4), .A (A), .B1 (n_0_1), .B2 (n_0_2));
AND3_X1 i_0_5 (.ZN (n_0_3), .A1 (A), .A2 (n_0_1), .A3 (n_0_2));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (B), .A2 (CIN));
OR2_X1 i_0_1 (.ZN (n_0_1), .A1 (B), .A2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));

endmodule //FA__4_131

module FA__4_127 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (SUM), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (B), .B1 (n_0_3), .B2 (n_0_0));
AND3_X1 i_0_5 (.ZN (n_0_4), .A1 (B), .A2 (n_0_3), .A3 (n_0_0));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
OAI21_X1 i_0_3 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
NOR2_X2 i_0_2 (.ZN (n_0_2), .A1 (A), .A2 (CIN));
INV_X1 i_0_1 (.ZN (n_0_1), .A (B));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (CIN));

endmodule //FA__4_127

module FA__4_123 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;


OAI22_X1 i_0_3 (.ZN (SUM), .A1 (n_0_0), .A2 (B), .B1 (A), .B2 (n_0_1));
NOR2_X2 i_0_2 (.ZN (COUT), .A1 (n_0_0), .A2 (n_0_1));
INV_X1 i_0_1 (.ZN (n_0_1), .A (B));
INV_X1 i_0_0 (.ZN (n_0_0), .A (A));

endmodule //FA__4_123

module FA__4_119 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_119

module FA__4_115 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;


OAI22_X1 i_0_3 (.ZN (SUM), .A1 (n_0_0), .A2 (B), .B1 (A), .B2 (n_0_1));
INV_X1 i_0_2 (.ZN (n_0_1), .A (B));
INV_X1 i_0_0 (.ZN (n_0_0), .A (A));
AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));

endmodule //FA__4_115

module FA__4_111 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;


OAI22_X2 i_0_3 (.ZN (SUM), .A1 (n_0_0), .A2 (B), .B1 (A), .B2 (n_0_1));
NOR2_X1 i_0_2 (.ZN (COUT), .A1 (n_0_0), .A2 (n_0_1));
INV_X1 i_0_1 (.ZN (n_0_1), .A (B));
INV_X2 i_0_0 (.ZN (n_0_0), .A (A));

endmodule //FA__4_111

module FA__4_107 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire slo__sro_n3;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XNOR2_X2 CLOCK_slo__sro_c9 (.ZN (SUM), .A (A), .B (slo__sro_n3));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n3), .A (B));

endmodule //FA__4_107

module FA__4_103 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire slo__mro_n5;


AND2_X4 i_0_1 (.ZN (COUT), .A1 (A), .A2 (B));
INV_X1 slo__mro_c6 (.ZN (slo__mro_n5), .A (B));
XNOR2_X2 slo__mro_c7 (.ZN (SUM), .A (A), .B (slo__mro_n5));

endmodule //FA__4_103

module FA__4_99 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;


OAI22_X1 i_0_3 (.ZN (SUM), .A1 (n_0_0), .A2 (B), .B1 (A), .B2 (n_0_1));
INV_X1 i_0_2 (.ZN (n_0_1), .A (B));
INV_X1 i_0_0 (.ZN (n_0_0), .A (A));
AND2_X2 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));

endmodule //FA__4_99

module FA__4_95 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (B), .A2 (A));
INV_X1 i_0_5 (.ZN (n_0_3), .A (B));
INV_X1 i_0_4 (.ZN (n_0_2), .A (A));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X2 i_0_2 (.ZN (n_0_0), .A1 (n_0_1), .A2 (n_0_4));
INV_X2 i_0_1 (.ZN (SUM), .A (n_0_0));
INV_X1 i_0_0 (.ZN (COUT), .A (n_0_4));

endmodule //FA__4_95

module FA__4_91 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_91

module FA__4_87 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_87

module FA__4_83 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_83

module FA__4_79 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire slo__mro_n3;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XNOR2_X2 slo__sro_c7 (.ZN (SUM), .A (A), .B (slo__mro_n3));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n3), .A (B));

endmodule //FA__4_79

module FA__4_75 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_75

module FA__4_71 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_71

module FA__4_67 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_67

module FA__4_63 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire opt_ipo_n2;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (opt_ipo_n2), .A (A), .B (B));
CLKBUF_X3 opt_ipo_c1 (.Z (SUM), .A (opt_ipo_n2));

endmodule //FA__4_63

module FA__4_59 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_59

module FA__4_55 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_55

module FA__4_51 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_51

module FA__4_47 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_47

module FA__4_43 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_43

module FA__4_39 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_39

module FA__4_35 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X2 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_35

module CSAlike (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__4_247 genblk1_61_fa (.COUT (carry[62]), .SUM (result[61]), .A (A[61]), .CIN (C[61]));
FA__4_243 genblk1_60_fa (.COUT (carry[61]), .SUM (result[60]), .A (A[60]), .B (B[60]), .CIN (C[60]));
FA__4_239 genblk1_59_fa (.COUT (carry[60]), .SUM (result[59]), .A (A[59]), .B (B[59]), .CIN (C[59]));
FA__4_235 genblk1_58_fa (.COUT (carry[59]), .SUM (result[58]), .A (A[58]), .B (B[58]), .CIN (C[58]));
FA__4_231 genblk1_57_fa (.COUT (carry[58]), .SUM (result[57]), .A (A[57]), .B (B[57]), .CIN (C[57]));
FA__4_227 genblk1_56_fa (.COUT (carry[57]), .SUM (result[56]), .A (A[56]), .B (B[56]), .CIN (C[56]));
FA__4_223 genblk1_55_fa (.COUT (carry[56]), .SUM (result[55]), .A (A[55]), .B (B[55]), .CIN (C[55]));
FA__4_219 genblk1_54_fa (.COUT (carry[55]), .SUM (result[54]), .A (A[54]), .B (B[54]), .CIN (C[54]));
FA__4_215 genblk1_53_fa (.COUT (carry[54]), .SUM (result[53]), .A (A[53]), .B (B[53]), .CIN (C[53]));
FA__4_211 genblk1_52_fa (.COUT (carry[53]), .SUM (result[52]), .A (A[52]), .B (B[52]), .CIN (C[52]));
FA__4_207 genblk1_51_fa (.COUT (carry[52]), .SUM (result[51]), .A (A[51]), .B (B[51]), .CIN (C[51]));
FA__4_203 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .B (B[50]), .CIN (C[50]));
FA__4_199 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .B (B[49]), .CIN (C[49]));
FA__4_195 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__4_191 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__4_187 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__4_183 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__4_179 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__4_175 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__4_171 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__4_167 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__4_163 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40])
    , .CIN (C[40]));
FA__4_159 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__4_155 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__4_151 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37])
    , .CIN (C[37]));
FA__4_147 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__4_143 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__4_139 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__4_135 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__4_131 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__4_127 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__4_123 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]));
FA__4_119 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]));
FA__4_115 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]));
FA__4_111 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]));
FA__4_107 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]));
FA__4_103 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]));
FA__4_99 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]));
FA__4_95 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]));
FA__4_91 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]));
FA__4_87 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]));
FA__4_83 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]));
FA__4_79 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]));
FA__4_75 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]));
FA__4_71 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]));
FA__4_67 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16]));
FA__4_63 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]));
FA__4_59 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]));
FA__4_55 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]));
FA__4_51 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12]));
FA__4_47 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]));
FA__4_43 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10]));
FA__4_39 genblk1_9_fa (.COUT (carry[10]), .SUM (result[9]), .A (A[9]), .B (B[9]));
FA__4_35 genblk1_8_fa (.COUT (carry[9]), .SUM (result[8]), .A (A[8]), .B (B[8]));

endmodule //CSAlike

module FA__4_1781 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_1781

module FA__4_1785 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_1785

module FA__4_1789 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_1789

module FA__4_1793 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_1793

module FA__4_1797 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_1797

module FA__4_1801 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1801

module FA__4_1805 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1805

module FA__4_1809 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1809

module FA__4_1813 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1813

module FA__4_1817 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1817

module FA__4_1821 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n3), .A (CIN));
XNOR2_X1 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n3));

endmodule //FA__4_1821

module FA__4_1825 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
XOR2_X1 slo__c1 (.Z (slo__n1), .A (A), .B (B));

endmodule //FA__4_1825

module FA__4_1829 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1829

module FA__4_1833 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n21;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X1 CLOCK_slo__sro_c9 (.ZN (CLOCK_slo__sro_n21), .A1 (A), .A2 (B));
AOI21_X1 CLOCK_slo__sro_c10 (.ZN (n_0_0), .A (CLOCK_slo__sro_n21), .B1 (temp), .B2 (CIN));

endmodule //FA__4_1833

module FA__4_1837 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1837

module FA__4_1841 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__mro_n4;
wire slo__mro_n5;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__mro_n4), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__mro_n4), .B (CIN));
INV_X1 slo__mro_c2 (.ZN (slo__mro_n5), .A (B));
XNOR2_X2 slo__mro_c3 (.ZN (slo__mro_n4), .A (A), .B (slo__mro_n5));

endmodule //FA__4_1841

module FA__4_1845 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1845

module FA__4_1849 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire CLOCK_opt_ipo_n15;
wire sgo__sro_n8;
wire CLOCK_slo__mro_n18;


INV_X2 CLOCK_slo__mro_c11 (.ZN (CLOCK_slo__mro_n18), .A (CIN));
INV_X2 CLOCK_opt_ipo_c10 (.ZN (CLOCK_opt_ipo_n15), .A (B));
XOR2_X2 i_0_0 (.Z (temp), .A (CLOCK_opt_ipo_n15), .B (A));
AND2_X1 sgo__sro_c3 (.ZN (sgo__sro_n8), .A1 (A), .A2 (CLOCK_opt_ipo_n15));
AOI21_X2 sgo__sro_c4 (.ZN (COUT), .A (sgo__sro_n8), .B1 (temp), .B2 (CIN));
XNOR2_X2 CLOCK_slo__mro_c12 (.ZN (SUM), .A (temp), .B (CLOCK_slo__mro_n18));

endmodule //FA__4_1849

module FA__4_1853 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire CLOCK_sgo__sro_n24;
wire CLOCK_sgo__sro_n25;


INV_X1 i_0_3 (.ZN (COUT), .A (CLOCK_sgo__sro_n24));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X1 CLOCK_sgo__sro_c10 (.ZN (CLOCK_sgo__sro_n25), .A1 (A), .A2 (B));
AOI21_X1 CLOCK_sgo__sro_c11 (.ZN (CLOCK_sgo__sro_n24), .A (CLOCK_sgo__sro_n25), .B1 (temp), .B2 (CIN));

endmodule //FA__4_1853

module FA__4_1857 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__mro_n82;
wire temp;
wire n_0_0;
wire slo__sro_n28;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
INV_X1 CLOCK_slo__mro_c50 (.ZN (CLOCK_slo__mro_n82), .A (B));
INV_X1 slo__sro_c16 (.ZN (slo__sro_n28), .A (CIN));
XNOR2_X1 slo__sro_c17 (.ZN (SUM), .A (temp), .B (slo__sro_n28));
XNOR2_X2 CLOCK_slo__mro_c51 (.ZN (temp), .A (CLOCK_slo__mro_n82), .B (A));

endmodule //FA__4_1857

module FA__4_1861 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));
AOI22_X1 slo__sro_c10 (.ZN (n_0_0), .A1 (temp), .A2 (CIN), .B1 (B), .B2 (A));

endmodule //FA__4_1861

module FA__4_1865 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n16;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 slo__sro_c12 (.ZN (slo__sro_n16), .A (B));
XNOR2_X2 slo__sro_c13 (.ZN (temp), .A (slo__sro_n16), .B (A));

endmodule //FA__4_1865

module FA__4_1869 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__mro_n16;
wire temp;
wire n_0_0;
wire slo__sro_n7;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
INV_X1 CLOCK_slo__mro_c9 (.ZN (CLOCK_slo__mro_n16), .A (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n7), .A (CIN));
XNOR2_X2 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n7));
XNOR2_X2 CLOCK_slo__mro_c10 (.ZN (temp), .A (CLOCK_slo__mro_n16), .B (A));

endmodule //FA__4_1869

module FA__4_1873 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (B), .A2 (A));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_6), .B2 (n_0_3));
NOR2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__4_1873

module FA__4_1877 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (SUM), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (CIN), .B1 (n_0_3), .B2 (n_0_0));
AND3_X2 i_0_5 (.ZN (n_0_4), .A1 (n_0_3), .A2 (n_0_0), .A3 (CIN));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_1));
OAI21_X1 i_0_3 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (CIN));
NOR2_X2 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__4_1877

module FA__4_1881 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NOR2_X2 i_0_7 (.ZN (SUM), .A1 (n_0_4), .A2 (n_0_5));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (CIN), .B1 (n_0_3), .B2 (n_0_0));
AND3_X2 i_0_5 (.ZN (n_0_4), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_0));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_1));
OAI21_X1 i_0_3 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (CIN));
NOR2_X2 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__4_1881

module FA__4_1885 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__sro_n38;
wire temp;
wire slo__n16;
wire slo__sro_n21;


AND2_X1 CLOCK_slo__sro_c25 (.ZN (CLOCK_slo__sro_n38), .A1 (A), .A2 (B));
AOI21_X2 CLOCK_slo__sro_c26 (.ZN (COUT), .A (CLOCK_slo__sro_n38), .B1 (slo__n16), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
XOR2_X1 slo__c9 (.Z (slo__n16), .A (A), .B (B));
INV_X1 slo__sro_c12 (.ZN (slo__sro_n21), .A (CIN));
XNOR2_X2 slo__sro_c13 (.ZN (SUM), .A (temp), .B (slo__sro_n21));

endmodule //FA__4_1885

module FA__4_1889 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X2 i_0_8 (.ZN (SUM), .A1 (n_0_5), .A2 (n_0_6));
AOI21_X2 i_0_7 (.ZN (n_0_6), .A (A), .B1 (n_0_3), .B2 (n_0_4));
AND3_X4 i_0_6 (.ZN (n_0_5), .A1 (A), .A2 (n_0_3), .A3 (n_0_4));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (B), .A2 (CIN));
OR2_X2 i_0_4 (.ZN (n_0_3), .A1 (B), .A2 (CIN));
INV_X1 i_0_3 (.ZN (n_0_2), .A (B));
INV_X1 i_0_2 (.ZN (n_0_1), .A (A));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
AOI21_X4 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_1));

endmodule //FA__4_1889

module FA__4_1893 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X2 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (A), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (A), .A3 (n_0_1));
NAND2_X2 i_0_1 (.ZN (n_0_1), .A1 (B), .A2 (CIN));
OR2_X2 i_0_0 (.ZN (n_0_0), .A1 (B), .A2 (CIN));

endmodule //FA__4_1893

module FA__4_1897 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X2 i_0_7 (.ZN (SUM), .A1 (n_0_4), .A2 (n_0_5));
OR3_X4 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (n_0_1), .A3 (CIN));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_3), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X1 i_0_3 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (CIN));
NOR2_X2 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__4_1897

module FA__4_1901 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


INV_X1 i_0_8 (.ZN (n_0_6), .A (CIN));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (A), .A2 (B));
NOR2_X2 i_0_6 (.ZN (n_0_4), .A1 (A), .A2 (B));
OAI21_X1 i_0_5 (.ZN (COUT), .A (n_0_5), .B1 (n_0_4), .B2 (n_0_6));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_4));
NAND3_X1 i_0_3 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_5));
INV_X1 i_0_2 (.ZN (n_0_1), .A (n_0_2));
AOI21_X2 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_5));
NOR2_X2 i_0_0 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));

endmodule //FA__4_1901

module FA__4_1905 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


XNOR2_X1 i_0_7 (.ZN (n_0_5), .A (B), .B (CIN));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (A), .A2 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_3), .A (A));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_5));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_2 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (B), .A2 (CIN));
OAI21_X1 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_3), .B2 (n_0_5));

endmodule //FA__4_1905

module FA__4_1909 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X4 i_0_6 (.ZN (SUM), .A1 (n_0_4), .A2 (n_0_3));
AOI21_X2 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X2 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X2 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (CIN), .A3 (n_0_1));
NAND2_X2 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
OR2_X4 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__4_1909

module FA__4_1913 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


NAND2_X2 i_0_7 (.ZN (SUM), .A1 (n_0_4), .A2 (n_0_5));
OAI21_X1 i_0_6 (.ZN (n_0_5), .A (A), .B1 (n_0_3), .B2 (n_0_2));
OR3_X4 i_0_5 (.ZN (n_0_4), .A1 (A), .A2 (n_0_3), .A3 (n_0_2));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_0));
OAI21_X2 i_0_3 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_2), .A1 (B), .A2 (CIN));
INV_X1 i_0_1 (.ZN (n_0_1), .A (A));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (B), .A2 (CIN));

endmodule //FA__4_1913

module FA__4_1917 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire CLOCK_slo__mro_n3;
wire CLOCK_slo__mro_n4;


INV_X1 i_0_5 (.ZN (n_0_2), .A (B));
INV_X1 i_0_4 (.ZN (n_0_1), .A (CIN));
OAI21_X1 i_0_3 (.ZN (n_0_0), .A (A), .B1 (B), .B2 (CIN));
OAI21_X1 i_0_2 (.ZN (COUT), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_1));
INV_X2 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n4), .A (CIN));
XNOR2_X2 CLOCK_slo__mro_c2 (.ZN (CLOCK_slo__mro_n3), .A (n_0_2), .B (CLOCK_slo__mro_n4));
XNOR2_X2 CLOCK_slo__mro_c3 (.ZN (SUM), .A (CLOCK_slo__mro_n3), .B (A));

endmodule //FA__4_1917

module FA__4_1921 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (CIN));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (B), .A2 (n_0_9));
INV_X1 i_0_9 (.ZN (n_0_7), .A (B));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (CIN));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (A), .A2 (n_0_8), .A3 (n_0_6));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_6), .A2 (n_0_8));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (n_0_4));
NAND2_X1 i_0_3 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_5));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (A), .A2 (B));
NOR2_X1 i_0_1 (.ZN (n_0_0), .A1 (A), .A2 (B));
OAI21_X2 i_0_0 (.ZN (COUT), .A (n_0_1), .B1 (n_0_0), .B2 (n_0_9));

endmodule //FA__4_1921

module FA__4_1925 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


NOR2_X1 i_0_9 (.ZN (n_0_7), .A1 (B), .A2 (CIN));
INV_X1 i_0_8 (.ZN (n_0_6), .A (n_0_7));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (B), .A2 (CIN));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (A), .A2 (n_0_4));
INV_X1 i_0_4 (.ZN (n_0_2), .A (A));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_4));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_0), .A2 (n_0_3));
AOI21_X1 i_0_0 (.ZN (COUT), .A (n_0_7), .B1 (n_0_2), .B2 (n_0_5));

endmodule //FA__4_1925

module FA__4_1929 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire sgo__sro_n9;
wire sgo__sro_n10;


AOI21_X2 i_0_8 (.ZN (SUM), .A (n_0_4), .B1 (A), .B2 (n_0_5));
OR2_X2 i_0_7 (.ZN (n_0_5), .A1 (n_0_2), .A2 (n_0_3));
NOR3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_2), .A2 (A), .A3 (n_0_3));
NOR2_X1 i_0_5 (.ZN (n_0_3), .A1 (B), .A2 (n_0_1));
AND2_X1 i_0_4 (.ZN (n_0_2), .A1 (B), .A2 (n_0_1));
INV_X1 i_0_1 (.ZN (n_0_1), .A (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X2 i_0_3 (.ZN (COUT), .A (sgo__sro_n9));
AND2_X1 sgo__sro_c8 (.ZN (sgo__sro_n10), .A1 (B), .A2 (A));
AOI21_X1 sgo__sro_c9 (.ZN (sgo__sro_n9), .A (sgo__sro_n10), .B1 (temp), .B2 (CIN));

endmodule //FA__4_1929

module FA__4_1933 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1933

module FA__4_1937 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire slo__sro_n3;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n3), .A (B));
XNOR2_X2 slo__sro_c2 (.ZN (SUM), .A (A), .B (slo__sro_n3));

endmodule //FA__4_1937

module FA__4_1941 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (B), .B (A));

endmodule //FA__4_1941

module FA__4_1945 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire slo__mro_n3;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n3), .A (A));
XNOR2_X2 slo__mro_c2 (.ZN (SUM), .A (slo__mro_n3), .B (B));

endmodule //FA__4_1945

module FA__4_1949 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1949

module FA__4_1953 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1953

module FA__4_1957 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1957

module FA__4_1961 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1961

module FA__4_1965 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (A));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (B));
INV_X1 i_0_3 (.ZN (n_0_1), .A (B));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (n_0_1));
NAND2_X1 i_0_0 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_0));
AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));

endmodule //FA__4_1965

module FA__4_1969 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1969

module FA__4_1973 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1973

module FA__4_1977 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1977

module FA__4_1981 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1981

module FA__4_1985 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X2 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1985

module FA__4_1989 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1989

module CSAlike__4_2018 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__4_1781 genblk1_59_fa (.COUT (carry[60]), .SUM (result[59]), .A (A[59]), .CIN (C[59]));
FA__4_1785 genblk1_58_fa (.COUT (carry[59]), .SUM (result[58]), .A (A[58]), .CIN (C[58]));
FA__4_1789 genblk1_57_fa (.COUT (carry[58]), .SUM (result[57]), .A (A[57]), .CIN (C[57]));
FA__4_1793 genblk1_56_fa (.COUT (carry[57]), .SUM (result[56]), .A (A[56]), .CIN (C[56]));
FA__4_1797 genblk1_55_fa (.COUT (carry[56]), .SUM (result[55]), .A (A[55]), .CIN (C[55]));
FA__4_1801 genblk1_54_fa (.COUT (carry[55]), .SUM (result[54]), .A (A[54]), .B (B[54]), .CIN (C[54]));
FA__4_1805 genblk1_53_fa (.COUT (carry[54]), .SUM (result[53]), .A (A[53]), .B (B[53]), .CIN (C[53]));
FA__4_1809 genblk1_52_fa (.COUT (carry[53]), .SUM (result[52]), .A (A[52]), .B (B[52]), .CIN (C[52]));
FA__4_1813 genblk1_51_fa (.COUT (carry[52]), .SUM (result[51]), .A (A[51]), .B (B[51]), .CIN (C[51]));
FA__4_1817 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .B (B[50]), .CIN (C[50]));
FA__4_1821 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .B (B[49]), .CIN (C[49]));
FA__4_1825 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__4_1829 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__4_1833 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__4_1837 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__4_1841 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__4_1845 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__4_1849 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__4_1853 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__4_1857 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__4_1861 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__4_1865 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__4_1869 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__4_1873 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__4_1877 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__4_1881 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__4_1885 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__4_1889 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__4_1893 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__4_1897 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__4_1901 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__4_1905 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__4_1909 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27])
    , .CIN (C[27]));
FA__4_1913 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__4_1917 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__4_1921 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__4_1925 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__4_1929 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__4_1933 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]));
FA__4_1937 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]));
FA__4_1941 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]));
FA__4_1945 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]));
FA__4_1949 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]));
FA__4_1953 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16]));
FA__4_1957 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]));
FA__4_1961 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]));
FA__4_1965 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]));
FA__4_1969 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12]));
FA__4_1973 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]));
FA__4_1977 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10]));
FA__4_1981 genblk1_9_fa (.COUT (carry[10]), .SUM (result[9]), .A (A[9]), .B (B[9]));
FA__4_1985 genblk1_8_fa (.COUT (carry[9]), .SUM (result[8]), .A (A[8]), .B (B[8]));
FA__4_1989 genblk1_7_fa (.COUT (carry[8]), .SUM (result[7]), .A (A[7]), .B (B[7]));

endmodule //CSAlike__4_2018

module FA__4_1552 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X2 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_1552

module FA__4_1556 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_1556

module FA__4_1560 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_1560

module FA__4_1564 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_1564

module FA__4_1568 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (CIN), .B (A));

endmodule //FA__4_1568

module FA__4_1572 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire slo__sro_n3;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n3), .A (A));
XNOR2_X2 slo__sro_c2 (.ZN (SUM), .A (CIN), .B (slo__sro_n3));

endmodule //FA__4_1572

module FA__4_1576 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (CIN), .B (A));

endmodule //FA__4_1576

module FA__4_1580 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X2 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (CIN), .B (A));

endmodule //FA__4_1580

module FA__4_1584 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1584

module FA__4_1588 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire sgo__sro_n7;
wire sgo__sro_n8;


INV_X1 i_0_3 (.ZN (COUT), .A (sgo__sro_n7));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X1 sgo__sro_c3 (.ZN (sgo__sro_n8), .A1 (B), .A2 (A));
AOI21_X1 sgo__sro_c4 (.ZN (sgo__sro_n7), .A (sgo__sro_n8), .B1 (CIN), .B2 (temp));

endmodule //FA__4_1588

module FA__4_1592 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire slo__sro_n10;
wire slo__sro_n11;


INV_X1 i_0_3 (.ZN (COUT), .A (slo__sro_n10));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X1 slo__sro_c4 (.ZN (slo__sro_n11), .A1 (A), .A2 (B));
AOI21_X1 slo__sro_c5 (.ZN (slo__sro_n10), .A (slo__sro_n11), .B1 (temp), .B2 (CIN));

endmodule //FA__4_1592

module FA__4_1596 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1596

module FA__4_1600 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;


AOI22_X2 i_0_2 (.ZN (COUT), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1600

module FA__4_1604 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n1;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n1), .A (B));
XNOR2_X2 slo__mro_c2 (.ZN (temp), .A (A), .B (slo__mro_n1));

endmodule //FA__4_1604

module FA__4_1608 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_opt_ipo_n12;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (CLOCK_opt_ipo_n12), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (CLOCK_opt_ipo_n12));
INV_X1 CLOCK_opt_ipo_c9 (.ZN (CLOCK_opt_ipo_n12), .A (B));

endmodule //FA__4_1608

module FA__4_1612 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n3;
wire CLOCK_slo__sro_n4;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n3), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n3), .B (CIN));
INV_X2 CLOCK_slo__sro_c3 (.ZN (CLOCK_slo__sro_n4), .A (B));
XNOR2_X2 CLOCK_slo__sro_c4 (.ZN (CLOCK_slo__sro_n3), .A (CLOCK_slo__sro_n4), .B (A));

endmodule //FA__4_1612

module FA__4_1616 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire CLOCK_slo__sro_n18;
wire CLOCK_slo__sro_n19;


INV_X1 i_0_3 (.ZN (COUT), .A (CLOCK_slo__sro_n18));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X1 CLOCK_slo__sro_c11 (.ZN (CLOCK_slo__sro_n19), .A1 (A), .A2 (B));
AOI21_X1 CLOCK_slo__sro_c12 (.ZN (CLOCK_slo__sro_n18), .A (CLOCK_slo__sro_n19), .B1 (temp), .B2 (CIN));

endmodule //FA__4_1616

module FA__4_1620 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire sgo__sro_n7;
wire sgo__sro_n8;


INV_X1 i_0_3 (.ZN (COUT), .A (sgo__sro_n7));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X1 sgo__sro_c3 (.ZN (sgo__sro_n8), .A1 (A), .A2 (B));
AOI21_X1 sgo__sro_c4 (.ZN (sgo__sro_n7), .A (sgo__sro_n8), .B1 (temp), .B2 (CIN));

endmodule //FA__4_1620

module FA__4_1624 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (B), .A2 (A));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X2 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__4_1624

module FA__4_1628 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire CLOCK_sgo__sro_n32;
wire opt_ipo_n21;
wire CLOCK_sgo__sro_n33;


INV_X1 i_0_3 (.ZN (COUT), .A (CLOCK_sgo__sro_n32));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (opt_ipo_n21));
AND2_X1 CLOCK_sgo__sro_c16 (.ZN (CLOCK_sgo__sro_n33), .A1 (A), .A2 (opt_ipo_n21));
INV_X1 opt_ipo_c9 (.ZN (opt_ipo_n21), .A (B));
AOI21_X1 CLOCK_sgo__sro_c17 (.ZN (CLOCK_sgo__sro_n32), .A (CLOCK_sgo__sro_n33), .B1 (temp), .B2 (CIN));

endmodule //FA__4_1628

module FA__4_1632 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1632

module FA__4_1636 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (B));
INV_X1 i_0_10 (.ZN (n_0_8), .A (CIN));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (B), .A2 (CIN));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (A), .A2 (n_0_7), .A3 (n_0_6));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (n_0_5));
INV_X2 i_0_2 (.ZN (SUM), .A (n_0_1));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
AOI21_X2 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_9), .B2 (n_0_4));

endmodule //FA__4_1636

module FA__4_1640 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (B), .A2 (A));
INV_X1 i_0_8 (.ZN (n_0_6), .A (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (A));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN));
AOI21_X2 i_0_3 (.ZN (n_0_1), .A (CIN), .B1 (B), .B2 (A));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_1), .A2 (n_0_4));
NAND2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_0));
AOI21_X2 i_0_0 (.ZN (COUT), .A (n_0_1), .B1 (n_0_6), .B2 (n_0_5));

endmodule //FA__4_1640

module FA__4_1644 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X2 i_0_12 (.ZN (n_0_10), .A (CIN));
NAND2_X2 i_0_11 (.ZN (n_0_9), .A1 (B), .A2 (n_0_10));
INV_X1 i_0_10 (.ZN (n_0_8), .A (B));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_8), .A2 (CIN));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_9));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (A));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_9), .A3 (n_0_7));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (n_0_5));
INV_X2 i_0_3 (.ZN (SUM), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (A), .A2 (B));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (A), .A2 (B));
OAI21_X2 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_10));

endmodule //FA__4_1644

module FA__4_1648 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (B));
INV_X1 i_0_9 (.ZN (n_0_7), .A (CIN));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (B), .A2 (CIN));
NAND3_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (A), .A3 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_3), .A (n_0_4));
AOI21_X1 i_0_4 (.ZN (n_0_2), .A (A), .B1 (n_0_6), .B2 (n_0_5));
NOR2_X2 i_0_3 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_1), .A (A));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
OAI21_X1 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_8), .B2 (n_0_1));

endmodule //FA__4_1648

module FA__4_1652 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (B));
INV_X1 i_0_9 (.ZN (n_0_7), .A (CIN));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (CIN), .A2 (B));
AOI21_X1 i_0_6 (.ZN (n_0_4), .A (A), .B1 (n_0_6), .B2 (n_0_5));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_6), .A2 (A), .A3 (n_0_5));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_3));
NOR2_X1 i_0_3 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_4));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (A), .A2 (B));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
NOR2_X2 i_0_0 (.ZN (COUT), .A1 (n_0_0), .A2 (n_0_1));

endmodule //FA__4_1652

module FA__4_1656 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


INV_X2 i_0_9 (.ZN (n_0_7), .A (CIN));
INV_X1 i_0_8 (.ZN (n_0_6), .A (B));
INV_X2 i_0_7 (.ZN (n_0_5), .A (A));
NAND2_X2 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_6));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (A), .A2 (B));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
AOI21_X2 i_0_3 (.ZN (n_0_1), .A (n_0_7), .B1 (A), .B2 (B));
AOI22_X2 i_0_2 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_7), .B1 (n_0_1), .B2 (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_4), .A2 (CIN));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_0), .A2 (n_0_3));

endmodule //FA__4_1656

module FA__4_1660 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (A), .A2 (B));
NAND2_X2 i_0_8 (.ZN (n_0_6), .A1 (n_0_2), .A2 (n_0_3));
NAND2_X2 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (CIN));
NAND2_X1 i_0_6 (.ZN (COUT), .A1 (n_0_5), .A2 (n_0_7));
NAND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_6), .A2 (CIN), .A3 (n_0_7));
INV_X1 i_0_4 (.ZN (n_0_3), .A (B));
INV_X1 i_0_3 (.ZN (n_0_2), .A (A));
INV_X1 i_0_2 (.ZN (n_0_1), .A (n_0_4));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (n_0_6), .B2 (n_0_7));
NOR2_X2 i_0_0 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));

endmodule //FA__4_1660

module FA__4_1664 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire CLOCK_sgo__n18;


NOR2_X4 i_0_8 (.ZN (SUM), .A1 (n_0_5), .A2 (n_0_6));
AOI21_X1 i_0_7 (.ZN (n_0_6), .A (B), .B1 (n_0_4), .B2 (n_0_3));
AND3_X2 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (B), .A3 (n_0_4));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (A), .A2 (CIN));
NAND2_X1 i_0_3 (.ZN (n_0_2), .A1 (B), .A2 (A));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (B), .A2 (A));
OAI21_X1 i_0_1 (.ZN (COUT), .A (n_0_2), .B1 (n_0_1), .B2 (n_0_0));
INV_X1 i_0_0 (.ZN (n_0_0), .A (CIN));
NOR2_X1 CLOCK_sgo__c36 (.ZN (CLOCK_sgo__n18), .A1 (A), .A2 (CIN));
INV_X1 CLOCK_sgo__c38 (.ZN (n_0_3), .A (CLOCK_sgo__n18));

endmodule //FA__4_1664

module FA__4_1668 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__4_1668

module FA__4_1672 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__mro_n20;
wire CLOCK_slo__mro_n21;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__mro_n20), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (CLOCK_slo__mro_n20), .B (CIN));
INV_X2 CLOCK_slo__mro_c12 (.ZN (CLOCK_slo__mro_n21), .A (A));
XNOR2_X2 CLOCK_slo__mro_c13 (.ZN (CLOCK_slo__mro_n20), .A (CLOCK_slo__mro_n21), .B (B));

endmodule //FA__4_1672

module FA__4_1676 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire opt_ipo_n4;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (opt_ipo_n4), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (opt_ipo_n4), .B (A));
INV_X1 opt_ipo_c2 (.ZN (opt_ipo_n4), .A (B));

endmodule //FA__4_1676

module FA__4_1680 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire sgo__sro_n7;
wire sgo__sro_n8;


INV_X1 i_0_3 (.ZN (COUT), .A (sgo__sro_n7));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X1 sgo__sro_c3 (.ZN (sgo__sro_n8), .A1 (A), .A2 (B));
AOI21_X2 sgo__sro_c4 (.ZN (sgo__sro_n7), .A (sgo__sro_n8), .B1 (temp), .B2 (CIN));

endmodule //FA__4_1680

module FA__4_1684 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__4_1684

module FA__4_1688 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


NAND2_X2 i_0_9 (.ZN (SUM), .A1 (n_0_5), .A2 (n_0_7));
NAND3_X1 i_0_8 (.ZN (n_0_7), .A1 (n_0_6), .A2 (n_0_2), .A3 (n_0_0));
INV_X1 i_0_7 (.ZN (n_0_6), .A (n_0_1));
OAI221_X1 i_0_6 (.ZN (n_0_5), .A (CIN), .B1 (A), .B2 (n_0_3), .C1 (n_0_4), .C2 (B));
INV_X1 i_0_5 (.ZN (n_0_4), .A (A));
INV_X1 i_0_4 (.ZN (n_0_3), .A (B));
OAI21_X1 i_0_3 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (CIN));
NOR2_X2 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
NAND2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__4_1688

module FA__4_1692 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire slo_n14;
wire n_0_0;
wire temp;
wire n_0_1;


XNOR2_X1 i_0_4 (.ZN (SUM), .A (slo_n14), .B (n_0_1));
XNOR2_X1 i_0_1 (.ZN (n_0_1), .A (B), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
CLKBUF_X1 slo___L1_c1_c3 (.Z (slo_n14), .A (A));

endmodule //FA__4_1692

module FA__4_1696 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1696

module FA__4_1700 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1700

module FA__4_1704 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X2 i_0_8 (.ZN (SUM), .A1 (n_0_5), .A2 (n_0_6));
AOI21_X1 i_0_7 (.ZN (n_0_6), .A (A), .B1 (n_0_3), .B2 (n_0_4));
AND3_X2 i_0_6 (.ZN (n_0_5), .A1 (A), .A2 (n_0_3), .A3 (n_0_4));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (B), .A2 (CIN));
OR2_X4 i_0_4 (.ZN (n_0_3), .A1 (B), .A2 (CIN));
NAND2_X1 i_0_3 (.ZN (n_0_2), .A1 (A), .A2 (B));
OR2_X1 i_0_2 (.ZN (n_0_1), .A1 (A), .A2 (B));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_1), .A2 (CIN));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_0), .A2 (n_0_2));

endmodule //FA__4_1704

module FA__4_1708 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1708

module FA__4_1712 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (A));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (B));
INV_X1 i_0_3 (.ZN (n_0_1), .A (B));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (n_0_1));
NAND2_X1 i_0_0 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_0));
AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));

endmodule //FA__4_1712

module FA__4_1716 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;


OAI22_X1 i_0_3 (.ZN (SUM), .A1 (n_0_0), .A2 (B), .B1 (A), .B2 (n_0_1));
INV_X1 i_0_2 (.ZN (n_0_1), .A (B));
INV_X1 i_0_0 (.ZN (n_0_0), .A (A));
AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));

endmodule //FA__4_1716

module FA__4_1720 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__mro_n3;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
INV_X2 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n3), .A (B));
XNOR2_X2 CLOCK_slo__mro_c2 (.ZN (SUM), .A (CLOCK_slo__mro_n3), .B (A));

endmodule //FA__4_1720

module FA__4_1724 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1724

module FA__4_1728 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1728

module FA__4_1732 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X2 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1732

module FA__4_1736 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1736

module FA__4_1740 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1740

module CSAlike__4_1765 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__4_1552 genblk1_53_fa (.COUT (carry[54]), .SUM (result[53]), .A (A[53]), .CIN (C[53]));
FA__4_1556 genblk1_52_fa (.COUT (carry[53]), .SUM (result[52]), .A (A[52]), .CIN (C[52]));
FA__4_1560 genblk1_51_fa (.COUT (carry[52]), .SUM (result[51]), .A (A[51]), .CIN (C[51]));
FA__4_1564 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .CIN (C[50]));
FA__4_1568 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .CIN (C[49]));
FA__4_1572 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .CIN (C[48]));
FA__4_1576 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .CIN (C[47]));
FA__4_1580 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .CIN (C[46]));
FA__4_1584 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__4_1588 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__4_1592 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__4_1596 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__4_1600 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41])
    , .CIN (C[41]));
FA__4_1604 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__4_1608 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__4_1612 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__4_1616 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__4_1620 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__4_1624 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__4_1628 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__4_1632 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__4_1636 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__4_1640 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__4_1644 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__4_1648 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__4_1652 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__4_1656 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27])
    , .CIN (C[27]));
FA__4_1660 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__4_1664 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__4_1668 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__4_1672 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__4_1676 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__4_1680 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__4_1684 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__4_1688 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__4_1692 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__4_1696 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]), .CIN (C[17]));
FA__4_1700 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16])
    , .CIN (C[16]));
FA__4_1704 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]), .CIN (C[15]));
FA__4_1708 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]));
FA__4_1712 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]));
FA__4_1716 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12]));
FA__4_1720 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]));
FA__4_1724 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10]));
FA__4_1728 genblk1_9_fa (.COUT (carry[10]), .SUM (result[9]), .A (A[9]), .B (B[9]));
FA__4_1732 genblk1_8_fa (.COUT (carry[9]), .SUM (result[8]), .A (A[8]), .B (B[8]));
FA__4_1736 genblk1_7_fa (.COUT (carry[8]), .SUM (result[7]), .A (A[7]), .B (B[7]));
FA__4_1740 genblk1_6_fa (.COUT (carry[7]), .SUM (result[6]), .A (A[6]), .B (B[6]));

endmodule //CSAlike__4_1765

module FA__4_1335 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_1335

module FA__4_1339 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_1339

module FA__4_1343 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (CIN), .B (A));

endmodule //FA__4_1343

module FA__4_1347 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (CIN), .B (A));

endmodule //FA__4_1347

module FA__4_1351 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__sro_n3;


AND2_X2 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n3), .A (A));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (SUM), .A (CIN), .B (CLOCK_slo__sro_n3));

endmodule //FA__4_1351

module FA__4_1355 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1355

module FA__4_1359 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;


AOI22_X2 i_0_2 (.ZN (COUT), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1359

module FA__4_1363 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n1;
wire CLOCK_slo__sro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n1), .B (CIN));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n2), .A (B));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (CLOCK_slo__sro_n1), .A (CLOCK_slo__sro_n2), .B (A));

endmodule //FA__4_1363

module FA__4_1367 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1367

module FA__4_1371 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n19;
wire CLOCK_slo__sro_n20;
wire slo__sro_n12;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n19), .B2 (CIN));
XNOR2_X2 CLOCK_slo__sro_c10 (.ZN (CLOCK_slo__sro_n19), .A (B), .B (CLOCK_slo__sro_n20));
INV_X1 CLOCK_slo__sro_c9 (.ZN (CLOCK_slo__sro_n20), .A (A));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n12), .A (CIN));
XNOR2_X2 slo__sro_c4 (.ZN (SUM), .A (slo__sro_n12), .B (CLOCK_slo__sro_n19));

endmodule //FA__4_1371

module FA__4_1375 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1375

module FA__4_1379 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;


XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AOI22_X1 slo__sro_c4 (.ZN (COUT), .A1 (temp), .A2 (CIN), .B1 (A), .B2 (B));

endmodule //FA__4_1379

module FA__4_1383 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (B), .A2 (A));
INV_X1 i_0_8 (.ZN (n_0_6), .A (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (A));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (CIN), .A3 (n_0_7));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_3));
AOI21_X1 i_0_3 (.ZN (n_0_1), .A (CIN), .B1 (n_0_4), .B2 (n_0_7));
NOR2_X2 i_0_2 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_1));
AOI21_X2 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
AOI21_X4 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_6), .B2 (n_0_5));

endmodule //FA__4_1383

module FA__4_1387 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (B));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (A), .A2 (CIN));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_3), .A2 (n_0_2));
NAND3_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_9), .A2 (n_0_8), .A3 (n_0_7));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (B));
NAND2_X1 i_0_5 (.ZN (SUM), .A1 (n_0_6), .A2 (n_0_4));
INV_X1 i_0_4 (.ZN (n_0_3), .A (A));
INV_X1 i_0_3 (.ZN (n_0_2), .A (CIN));
AOI21_X1 i_0_2 (.ZN (n_0_1), .A (CIN), .B1 (B), .B2 (A));
NOR2_X1 i_0_1 (.ZN (n_0_0), .A1 (B), .A2 (A));
NOR2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_1), .A2 (n_0_0));

endmodule //FA__4_1387

module FA__4_1391 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


NAND2_X1 i_0_12 (.ZN (n_0_10), .A1 (B), .A2 (CIN));
OAI21_X1 i_0_11 (.ZN (n_0_9), .A (n_0_10), .B1 (B), .B2 (CIN));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (n_0_9), .A2 (A));
INV_X1 i_0_9 (.ZN (n_0_7), .A (A));
INV_X1 i_0_8 (.ZN (n_0_6), .A (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (CIN));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_7), .A2 (n_0_10), .A3 (n_0_4));
NAND2_X1 i_0_4 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_8));
NOR2_X1 i_0_3 (.ZN (n_0_2), .A1 (A), .A2 (B));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (A), .A2 (B));
OAI21_X2 i_0_1 (.ZN (COUT), .A (n_0_1), .B1 (n_0_2), .B2 (n_0_5));

endmodule //FA__4_1391

module FA__4_1395 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


NOR2_X1 i_0_12 (.ZN (n_0_10), .A1 (B), .A2 (CIN));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (B), .A2 (CIN));
OAI21_X2 i_0_10 (.ZN (COUT), .A (n_0_9), .B1 (n_0_10), .B2 (n_0_2));
INV_X1 i_0_9 (.ZN (n_0_8), .A (B));
NOR2_X1 i_0_8 (.ZN (n_0_7), .A1 (A), .A2 (B));
NAND2_X1 i_0_7 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_6 (.ZN (n_0_5), .A (n_0_6));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_5), .B2 (n_0_7));
INV_X1 i_0_4 (.ZN (n_0_3), .A (CIN));
INV_X1 i_0_3 (.ZN (n_0_2), .A (A));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (n_0_2), .A2 (n_0_8));
NAND3_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_1), .A2 (n_0_3), .A3 (n_0_6));
NAND2_X1 i_0_0 (.ZN (SUM), .A1 (n_0_4), .A2 (n_0_0));

endmodule //FA__4_1395

module FA__4_1399 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__4_1399

module FA__4_1403 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire slo__sro_n6;
wire slo__sro_n7;
wire slo__sro_n8;


INV_X1 i_0_8 (.ZN (n_0_6), .A (CIN));
NOR2_X1 i_0_7 (.ZN (n_0_5), .A1 (B), .A2 (A));
NOR2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_0), .A2 (n_0_5));
NOR2_X1 slo__sro_c8 (.ZN (slo__sro_n8), .A1 (A), .A2 (B));
OAI21_X2 i_0_3 (.ZN (SUM), .A (slo__sro_n6), .B1 (n_0_4), .B2 (n_0_6));
NOR2_X1 i_0_2 (.ZN (COUT), .A1 (n_0_3), .A2 (n_0_5));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (B), .A2 (A));
INV_X1 i_0_0 (.ZN (n_0_0), .A (n_0_1));
AOI21_X2 slo__sro_c4 (.ZN (n_0_3), .A (CIN), .B1 (A), .B2 (B));
INV_X1 slo__sro_c9 (.ZN (slo__sro_n7), .A (slo__sro_n8));
NAND2_X2 slo__sro_c10 (.ZN (slo__sro_n6), .A1 (n_0_3), .A2 (slo__sro_n7));

endmodule //FA__4_1403

module FA__4_1407 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (A));
INV_X1 i_0_9 (.ZN (n_0_7), .A (CIN));
XNOR2_X2 i_0_8 (.ZN (n_0_6), .A (B), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (A), .A2 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
INV_X2 i_0_3 (.ZN (SUM), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (A), .A2 (B));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (A), .A2 (B));
OAI21_X2 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_7));

endmodule //FA__4_1407

module FA__4_1411 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n5;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 CLOCK_slo__mro_c5 (.ZN (CLOCK_slo__mro_n5), .A (B));
XNOR2_X2 CLOCK_slo__mro_c6 (.ZN (temp), .A (A), .B (CLOCK_slo__mro_n5));

endmodule //FA__4_1411

module FA__4_1415 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_11 (.ZN (n_0_8), .A (B));
INV_X1 i_0_10 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_9 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_5), .A1 (A), .A2 (B));
AOI21_X1 i_0_7 (.ZN (n_0_4), .A (CIN), .B1 (n_0_6), .B2 (n_0_5));
NAND3_X1 i_0_6 (.ZN (n_0_3), .A1 (n_0_6), .A2 (CIN), .A3 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_2), .A (n_0_3));
NOR2_X1 i_0_4 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_0 (.ZN (temp), .A (n_0_1));
INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));

endmodule //FA__4_1415

module FA__4_1419 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_11 (.ZN (n_0_8), .A (B));
INV_X1 i_0_10 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_9 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_5), .A1 (A), .A2 (B));
AOI21_X2 i_0_7 (.ZN (n_0_4), .A (CIN), .B1 (n_0_6), .B2 (n_0_5));
NAND3_X1 i_0_6 (.ZN (n_0_3), .A1 (n_0_6), .A2 (CIN), .A3 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_2), .A (n_0_3));
NOR2_X2 i_0_4 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_0 (.ZN (temp), .A (n_0_1));
INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));

endmodule //FA__4_1419

module FA__4_1423 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n16;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 slo__mro_c12 (.ZN (slo__mro_n16), .A (B));
XNOR2_X2 slo__mro_c13 (.ZN (temp), .A (slo__mro_n16), .B (A));

endmodule //FA__4_1423

module FA__4_1427 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire slo__mro_n10;
wire slo__mro_n11;


AOI22_X1 i_0_2 (.ZN (COUT), .A1 (A), .A2 (B), .B1 (slo__mro_n10), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__mro_n10), .B (CIN));
INV_X1 slo__mro_c4 (.ZN (slo__mro_n11), .A (B));
XNOR2_X2 slo__mro_c5 (.ZN (slo__mro_n10), .A (A), .B (slo__mro_n11));

endmodule //FA__4_1427

module FA__4_1431 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n3), .A (B));
XNOR2_X2 slo__sro_c4 (.ZN (temp), .A (A), .B (slo__sro_n3));

endmodule //FA__4_1431

module FA__4_1435 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__sro_n1;
wire slo__sro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__sro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__sro_n1), .B (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n2), .A (B));
XNOR2_X2 slo__sro_c2 (.ZN (slo__sro_n1), .A (slo__sro_n2), .B (A));

endmodule //FA__4_1435

module FA__4_1439 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n6;
wire CLOCK_slo__sro_n7;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n6), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n6), .B (CIN));
INV_X2 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n7), .A (B));
XNOR2_X2 CLOCK_slo__sro_c2 (.ZN (CLOCK_slo__sro_n6), .A (A), .B (CLOCK_slo__sro_n7));

endmodule //FA__4_1439

module FA__4_1443 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1443

module FA__4_1447 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__mro_n1;
wire slo__mro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__mro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__mro_n1), .B (CIN));
INV_X2 slo__mro_c1 (.ZN (slo__mro_n2), .A (B));
XNOR2_X2 slo__mro_c2 (.ZN (slo__mro_n1), .A (A), .B (slo__mro_n2));

endmodule //FA__4_1447

module FA__4_1451 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_sgo__sro_n30;
wire CLOCK_sgo__sro_n31;
wire CLOCK_slo__sro_n38;
wire CLOCK_slo__sro_n39;


INV_X1 i_0_3 (.ZN (COUT), .A (CLOCK_sgo__sro_n30));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n38), .B (CIN));
AND2_X1 CLOCK_sgo__sro_c16 (.ZN (CLOCK_sgo__sro_n31), .A1 (A), .A2 (B));
AOI21_X1 CLOCK_sgo__sro_c17 (.ZN (CLOCK_sgo__sro_n30), .A (CLOCK_sgo__sro_n31), .B1 (CLOCK_slo__sro_n38), .B2 (CIN));
INV_X1 CLOCK_slo__sro_c24 (.ZN (CLOCK_slo__sro_n39), .A (A));
XNOR2_X2 CLOCK_slo__sro_c25 (.ZN (CLOCK_slo__sro_n38), .A (CLOCK_slo__sro_n39), .B (B));

endmodule //FA__4_1451

module FA__4_1455 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X2 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND3_X2 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X2 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X2 CLOCK_slo__mro_c2 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__4_1455

module FA__4_1459 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;


AOI21_X1 i_0_8 (.ZN (SUM), .A (n_0_4), .B1 (A), .B2 (n_0_5));
OR2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_2), .A2 (n_0_3));
NOR3_X1 i_0_6 (.ZN (n_0_4), .A1 (A), .A2 (n_0_2), .A3 (n_0_3));
NOR2_X1 i_0_5 (.ZN (n_0_3), .A1 (B), .A2 (n_0_1));
AND2_X1 i_0_4 (.ZN (n_0_2), .A1 (B), .A2 (n_0_1));
INV_X1 i_0_1 (.ZN (n_0_1), .A (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));

endmodule //FA__4_1459

module FA__4_1463 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (B));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (A), .A2 (n_0_9));
INV_X1 i_0_9 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_7), .A2 (B));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (CIN), .A3 (n_0_8));
INV_X1 i_0_6 (.ZN (n_0_4), .A (CIN));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (A), .A2 (B));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_7), .A2 (n_0_9));
NAND3_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (n_0_4), .A3 (n_0_3));
NAND2_X1 i_0_2 (.ZN (SUM), .A1 (n_0_5), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_2), .A2 (CIN));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_0), .A2 (n_0_3));

endmodule //FA__4_1463

module FA__4_1467 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X2 i_0_8 (.ZN (SUM), .A1 (n_0_5), .A2 (n_0_6));
AOI21_X1 i_0_7 (.ZN (n_0_6), .A (A), .B1 (n_0_3), .B2 (n_0_4));
AND3_X2 i_0_6 (.ZN (n_0_5), .A1 (A), .A2 (n_0_3), .A3 (n_0_4));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (B), .A2 (CIN));
OR2_X2 i_0_4 (.ZN (n_0_3), .A1 (B), .A2 (CIN));
NAND2_X1 i_0_3 (.ZN (n_0_2), .A1 (A), .A2 (B));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (A), .A2 (B));
OAI21_X1 i_0_1 (.ZN (COUT), .A (n_0_2), .B1 (n_0_1), .B2 (n_0_0));
INV_X1 i_0_0 (.ZN (n_0_0), .A (CIN));

endmodule //FA__4_1467

module FA__4_1471 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X4 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X2 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X2 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X2 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (CIN), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__4_1471

module FA__4_1475 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (A));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (B), .A2 (n_0_3));
INV_X1 i_0_3 (.ZN (n_0_1), .A (B));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_1), .A2 (A));
NAND2_X2 i_0_0 (.ZN (SUM), .A1 (n_0_0), .A2 (n_0_2));
AND2_X4 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));

endmodule //FA__4_1475

module FA__4_1479 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire slo__sro_n3;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
INV_X2 slo__sro_c1 (.ZN (slo__sro_n3), .A (B));
XNOR2_X1 slo__sro_c2 (.ZN (SUM), .A (slo__sro_n3), .B (A));

endmodule //FA__4_1479

module FA__4_1483 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1483

module FA__4_1487 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1487

module FA__4_1491 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1491

module CSAlike__4_1512 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__4_1335 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .CIN (C[44]));
FA__4_1339 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .CIN (C[43]));
FA__4_1343 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .CIN (C[42]));
FA__4_1347 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .CIN (C[41]));
FA__4_1351 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .CIN (C[40]));
FA__4_1355 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__4_1359 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__4_1363 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__4_1367 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__4_1371 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35])
    , .CIN (C[35]));
FA__4_1375 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__4_1379 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33])
    , .CIN (C[33]));
FA__4_1383 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__4_1387 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__4_1391 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__4_1395 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__4_1399 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__4_1403 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27])
    , .CIN (C[27]));
FA__4_1407 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__4_1411 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__4_1415 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__4_1419 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__4_1423 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__4_1427 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__4_1431 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__4_1435 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__4_1439 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__4_1443 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]), .CIN (C[17]));
FA__4_1447 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16])
    , .CIN (C[16]));
FA__4_1451 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]), .CIN (C[15]));
FA__4_1455 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]), .CIN (C[14]));
FA__4_1459 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]), .CIN (C[13]));
FA__4_1463 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12]), .CIN (C[12]));
FA__4_1467 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]), .CIN (C[11]));
FA__4_1471 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10])
    , .CIN (C[10]));
FA__4_1475 genblk1_9_fa (.COUT (carry[10]), .SUM (result[9]), .A (A[9]), .B (B[9]));
FA__4_1479 genblk1_8_fa (.COUT (carry[9]), .SUM (result[8]), .A (A[8]), .B (B[8]));
FA__4_1483 genblk1_7_fa (.COUT (carry[8]), .SUM (result[7]), .A (A[7]), .B (B[7]));
FA__4_1487 genblk1_6_fa (.COUT (carry[7]), .SUM (result[6]), .A (A[6]), .B (B[6]));
FA__4_1491 genblk1_5_fa (.COUT (carry[6]), .SUM (result[5]), .A (A[5]), .B (B[5]));

endmodule //CSAlike__4_1512

module FA__4_1026 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_1026

module FA__4_1030 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_1030

module FA__4_1034 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_1034

module FA__4_1038 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_1038

module FA__4_1042 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_1042

module FA__4_1046 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X2 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_1046

module FA__4_1050 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X2 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_1050

module FA__4_1054 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_1054

module FA__4_1058 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1058

module FA__4_1062 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1062

module FA__4_1066 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__mro_n1;
wire CLOCK_slo__mro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__mro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__mro_n1), .B (CIN));
INV_X2 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n2), .A (A));
XNOR2_X2 CLOCK_slo__mro_c2 (.ZN (CLOCK_slo__mro_n1), .A (B), .B (CLOCK_slo__mro_n2));

endmodule //FA__4_1066

module FA__4_1070 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));
INV_X1 CLOCK_slo__sro_c5 (.ZN (CLOCK_slo__sro_n7), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c6 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n7));

endmodule //FA__4_1070

module FA__4_1074 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__4_1074

module FA__4_1078 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1078

module FA__4_1082 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1082

module FA__4_1086 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n1;
wire slo__mro_n5;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
INV_X1 slo__mro_c7 (.ZN (slo__mro_n5), .A (CIN));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n1), .A (A));
XNOR2_X2 slo__mro_c2 (.ZN (temp), .A (B), .B (slo__mro_n1));
XNOR2_X2 slo__mro_c8 (.ZN (SUM), .A (temp), .B (slo__mro_n5));

endmodule //FA__4_1086

module FA__4_1090 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n3;
wire slo__sro_n12;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n3), .A (CIN));
XNOR2_X2 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n3));
INV_X1 slo__sro_c9 (.ZN (slo__sro_n12), .A (A));
XNOR2_X2 slo__sro_c10 (.ZN (temp), .A (slo__sro_n12), .B (B));

endmodule //FA__4_1090

module FA__4_1094 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1094

module FA__4_1098 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1098

module FA__4_1102 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__sro_n10;
wire temp;
wire n_0_0;
wire slo__mro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
INV_X2 CLOCK_slo__sro_c7 (.ZN (CLOCK_slo__sro_n10), .A (A));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n3), .A (CIN));
XNOR2_X1 slo__mro_c2 (.ZN (SUM), .A (temp), .B (slo__mro_n3));
XNOR2_X2 CLOCK_slo__sro_c8 (.ZN (temp), .A (CLOCK_slo__sro_n10), .B (B));

endmodule //FA__4_1102

module FA__4_1106 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1106

module FA__4_1110 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n1;
wire CLOCK_slo__sro_n8;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
INV_X1 CLOCK_slo__sro_c10 (.ZN (CLOCK_slo__sro_n8), .A (CIN));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n1), .A (A));
XNOR2_X1 slo__mro_c2 (.ZN (temp), .A (slo__mro_n1), .B (B));
XNOR2_X1 CLOCK_slo__sro_c11 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n8));

endmodule //FA__4_1110

module FA__4_1114 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n1;
wire slo__sro_n6;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
INV_X1 slo__sro_c8 (.ZN (slo__sro_n6), .A (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n1), .A (A));
XNOR2_X2 slo__sro_c2 (.ZN (temp), .A (B), .B (slo__sro_n1));
XNOR2_X2 slo__sro_c9 (.ZN (SUM), .A (temp), .B (slo__sro_n6));

endmodule //FA__4_1114

module FA__4_1118 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n1), .A (A));
XNOR2_X2 slo__sro_c2 (.ZN (temp), .A (slo__sro_n1), .B (B));

endmodule //FA__4_1118

module FA__4_1122 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1122

module FA__4_1126 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1126

module FA__4_1130 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1130

module FA__4_1134 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1134

module FA__4_1138 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1138

module FA__4_1142 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1142

module FA__4_1146 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_1146

module FA__4_1150 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__mro_n1;
wire slo__mro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__mro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__mro_n1), .B (CIN));
INV_X2 slo__mro_c1 (.ZN (slo__mro_n2), .A (A));
XNOR2_X2 slo__mro_c2 (.ZN (slo__mro_n1), .A (B), .B (slo__mro_n2));

endmodule //FA__4_1150

module FA__4_1154 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n3), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n3));

endmodule //FA__4_1154

module FA__4_1158 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n3), .A (CIN));
XNOR2_X2 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n3));

endmodule //FA__4_1158

module FA__4_1162 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1162

module FA__4_1166 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1166

module FA__4_1170 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1170

module FA__4_1174 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_1174

module CSAlike__4_1259 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__4_1026 genblk1_58_fa (.COUT (carry[59]), .SUM (result[58]), .B (B[58]), .CIN (C[58]));
FA__4_1030 genblk1_57_fa (.COUT (carry[58]), .SUM (result[57]), .B (B[57]), .CIN (C[57]));
FA__4_1034 genblk1_56_fa (.COUT (carry[57]), .SUM (result[56]), .B (B[56]), .CIN (C[56]));
FA__4_1038 genblk1_55_fa (.COUT (carry[56]), .SUM (result[55]), .B (B[55]), .CIN (C[55]));
FA__4_1042 genblk1_54_fa (.COUT (carry[55]), .SUM (result[54]), .B (B[54]), .CIN (C[54]));
FA__4_1046 genblk1_53_fa (.COUT (carry[54]), .SUM (result[53]), .B (B[53]), .CIN (C[53]));
FA__4_1050 genblk1_52_fa (.COUT (carry[53]), .SUM (result[52]), .B (B[52]), .CIN (C[52]));
FA__4_1054 genblk1_51_fa (.COUT (carry[52]), .SUM (result[51]), .B (B[51]), .CIN (C[51]));
FA__4_1058 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .B (B[50])
    , .CIN (C[50]));
FA__4_1062 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .B (B[49]), .CIN (C[49]));
FA__4_1066 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__4_1070 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__4_1074 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__4_1078 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__4_1082 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__4_1086 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__4_1090 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__4_1094 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__4_1098 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__4_1102 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__4_1106 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__4_1110 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__4_1114 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__4_1118 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__4_1122 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__4_1126 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__4_1130 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__4_1134 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31])
    , .CIN (C[31]));
FA__4_1138 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__4_1142 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__4_1146 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__4_1150 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27])
    , .CIN (C[27]));
FA__4_1154 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__4_1158 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__4_1162 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]));
FA__4_1166 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]));
FA__4_1170 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]));
FA__4_1174 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]));

endmodule //CSAlike__4_1259

module FA__4_853 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_853

module FA__4_857 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__4_857

module FA__4_861 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n10;
wire CLOCK_slo__sro_n11;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
NAND2_X1 CLOCK_slo__sro_c4 (.ZN (CLOCK_slo__sro_n11), .A1 (A), .A2 (B));
INV_X1 CLOCK_slo__sro_c5 (.ZN (CLOCK_slo__sro_n10), .A (CLOCK_slo__sro_n11));
AOI21_X1 CLOCK_slo__sro_c6 (.ZN (n_0_0), .A (CLOCK_slo__sro_n10), .B1 (CIN), .B2 (temp));

endmodule //FA__4_861

module FA__4_865 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_865

module FA__4_869 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_869

module FA__4_873 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (B), .A2 (A));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X2 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__4_873

module FA__4_877 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (A), .A2 (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_5));
OAI21_X1 i_0_5 (.ZN (n_0_3), .A (CIN), .B1 (n_0_4), .B2 (n_0_6));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_6));
AOI21_X1 i_0_3 (.ZN (n_0_1), .A (CIN), .B1 (A), .B2 (B));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_0));
NOR2_X2 i_0_0 (.ZN (COUT), .A1 (n_0_1), .A2 (n_0_6));

endmodule //FA__4_877

module FA__4_881 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


INV_X1 i_0_12 (.ZN (n_0_10), .A (A));
INV_X1 i_0_11 (.ZN (n_0_9), .A (B));
INV_X1 i_0_10 (.ZN (n_0_8), .A (CIN));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (B), .A2 (CIN));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_10), .A2 (n_0_5));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (A), .A2 (n_0_7), .A3 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
INV_X1 i_0_3 (.ZN (SUM), .A (n_0_2));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (A), .A2 (B));
NOR2_X1 i_0_1 (.ZN (n_0_0), .A1 (A), .A2 (B));
OAI21_X2 i_0_0 (.ZN (COUT), .A (n_0_1), .B1 (n_0_0), .B2 (n_0_8));

endmodule //FA__4_881

module FA__4_885 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X1 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (A), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (A), .A2 (n_0_0), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (B), .A2 (CIN));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (B), .A2 (CIN));

endmodule //FA__4_885

module FA__4_889 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X1 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (A), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (A), .A2 (n_0_0), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (B), .A2 (CIN));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (B), .A2 (CIN));

endmodule //FA__4_889

module FA__4_893 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (A));
INV_X1 i_0_9 (.ZN (n_0_7), .A (CIN));
XNOR2_X1 i_0_8 (.ZN (n_0_6), .A (B), .B (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (A), .A2 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_4), .A2 (n_0_3));
INV_X1 i_0_3 (.ZN (SUM), .A (n_0_2));
NOR2_X1 i_0_2 (.ZN (n_0_1), .A1 (A), .A2 (B));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (A), .A2 (B));
OAI21_X1 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_7));

endmodule //FA__4_893

module FA__4_897 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


OR2_X2 i_0_10 (.ZN (n_0_8), .A1 (B), .A2 (CIN));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (B), .A2 (CIN));
NAND3_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (n_0_8), .A3 (n_0_7));
INV_X1 i_0_7 (.ZN (n_0_5), .A (A));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (n_0_6));
INV_X1 i_0_3 (.ZN (SUM), .A (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_1), .A (B));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
AOI21_X1 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_5));

endmodule //FA__4_897

module FA__4_901 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


AOI22_X2 i_0_6 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_3), .B1 (n_0_4), .B2 (A));
INV_X1 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X1 i_0_4 (.ZN (n_0_3), .A (CIN), .B (B));
INV_X1 i_0_2 (.ZN (n_0_2), .A (B));
INV_X1 i_0_1 (.ZN (n_0_1), .A (A));
OAI21_X1 i_0_0 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
OAI21_X4 CLOCK_slo__sro_c4 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));

endmodule //FA__4_901

module FA__4_905 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire opt_ipo_n7;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


AOI22_X2 i_0_6 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_3), .B1 (n_0_4), .B2 (A));
INV_X2 i_0_5 (.ZN (n_0_4), .A (n_0_3));
XNOR2_X2 i_0_4 (.ZN (n_0_3), .A (B), .B (CIN));
OAI21_X1 i_0_3 (.ZN (opt_ipo_n7), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (B));
INV_X1 i_0_1 (.ZN (n_0_1), .A (A));
OAI21_X1 i_0_0 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
BUF_X1 opt_ipo_c6 (.Z (COUT), .A (opt_ipo_n7));

endmodule //FA__4_905

module FA__4_909 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X2 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X2 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__4_909

module FA__4_913 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (A), .A2 (B));
INV_X1 i_0_8 (.ZN (n_0_6), .A (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (A));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_6));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (CIN), .A3 (n_0_7));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_3));
AOI21_X1 i_0_3 (.ZN (n_0_1), .A (CIN), .B1 (n_0_4), .B2 (n_0_7));
NOR2_X2 i_0_2 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_1));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
AOI21_X1 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_6), .B2 (n_0_5));

endmodule //FA__4_913

module FA__4_917 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X2 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__4_917

module FA__4_921 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire opt_ipo_n20;
wire temp;
wire n_0_0;
wire slo__mro_n17;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (opt_ipo_n20), .A (temp), .B (CIN));
BUF_X4 opt_ipo_c17 (.Z (SUM), .A (opt_ipo_n20));
INV_X1 slo__mro_c11 (.ZN (slo__mro_n17), .A (B));
XNOR2_X2 slo__mro_c12 (.ZN (temp), .A (slo__mro_n17), .B (A));

endmodule //FA__4_921

module FA__4_925 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire opt_ipo_n13;
wire temp;
wire n_0_0;
wire slo__mro_n10;
wire opt_ipo_n14;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (opt_ipo_n14), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (opt_ipo_n13), .A (temp), .B (CIN));
BUF_X4 opt_ipo_c10 (.Z (SUM), .A (opt_ipo_n13));
INV_X2 slo__mro_c4 (.ZN (slo__mro_n10), .A (A));
XNOR2_X2 slo__mro_c5 (.ZN (temp), .A (slo__mro_n10), .B (opt_ipo_n14));
INV_X1 opt_ipo_c11 (.ZN (opt_ipo_n14), .A (B));

endmodule //FA__4_925

module FA__4_929 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X2 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__4_929

module FA__4_933 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire opt_ipo_n5;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (opt_ipo_n5), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
BUF_X4 opt_ipo_c2 (.Z (SUM), .A (opt_ipo_n5));

endmodule //FA__4_933

module FA__4_937 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_937

module FA__4_941 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n15;
wire CLOCK_slo__sro_n16;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n15), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n15), .B (CIN));
INV_X2 CLOCK_slo__sro_c14 (.ZN (CLOCK_slo__sro_n16), .A (A));
XNOR2_X2 CLOCK_slo__sro_c15 (.ZN (CLOCK_slo__sro_n15), .A (CLOCK_slo__sro_n16), .B (B));

endmodule //FA__4_941

module FA__4_945 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo_n64;
wire temp;
wire n_0_0;
wire CLOCK_slo__n54;
wire opt_ipo_n23;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X4 i_0_2 (.ZN (n_0_0), .A1 (CLOCK_slo_n64), .A2 (opt_ipo_n23), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__n54), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (opt_ipo_n23));
XOR2_X2 CLOCK_slo__c31 (.Z (CLOCK_slo__n54), .A (A), .B (opt_ipo_n23));
INV_X2 opt_ipo_c13 (.ZN (opt_ipo_n23), .A (B));
CLKBUF_X1 CLOCK_slo___L1_c1_c34 (.Z (CLOCK_slo_n64), .A (A));

endmodule //FA__4_945

module FA__4_949 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_949

module FA__4_953 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (A));
NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (n_0_9), .A2 (B));
INV_X1 i_0_9 (.ZN (n_0_7), .A (B));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (n_0_7));
NAND3_X1 i_0_7 (.ZN (n_0_5), .A1 (CIN), .A2 (n_0_8), .A3 (n_0_6));
INV_X1 i_0_6 (.ZN (n_0_4), .A (CIN));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (n_0_6));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (n_0_4));
NAND2_X2 i_0_3 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_5));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (A), .A2 (B));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_3), .A2 (CIN));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_0), .A2 (n_0_1));

endmodule //FA__4_953

module FA__4_957 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X2 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (CIN), .A2 (n_0_0), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
OR2_X2 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__4_957

module FA__4_961 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__4_961

module FA__4_965 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X1 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (CIN), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
OR2_X2 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__4_965

module FA__4_969 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (A), .A2 (B));
NAND2_X2 i_0_8 (.ZN (n_0_6), .A1 (n_0_2), .A2 (n_0_3));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (CIN));
NAND2_X1 i_0_6 (.ZN (COUT), .A1 (n_0_5), .A2 (n_0_7));
NAND3_X1 i_0_5 (.ZN (n_0_4), .A1 (n_0_6), .A2 (CIN), .A3 (n_0_7));
INV_X1 i_0_4 (.ZN (n_0_3), .A (B));
INV_X1 i_0_3 (.ZN (n_0_2), .A (A));
INV_X1 i_0_2 (.ZN (n_0_1), .A (n_0_4));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (n_0_6), .B2 (n_0_7));
NOR2_X2 i_0_0 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));

endmodule //FA__4_969

module FA__4_973 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire opt_ipo_n6;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (opt_ipo_n6), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (opt_ipo_n6), .B (A));
INV_X1 opt_ipo_c4 (.ZN (opt_ipo_n6), .A (B));

endmodule //FA__4_973

module FA__4_977 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n12;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X2 CLOCK_slo__sro_c6 (.ZN (CLOCK_slo__sro_n12), .A (B));
XNOR2_X2 CLOCK_slo__sro_c7 (.ZN (temp), .A (CLOCK_slo__sro_n12), .B (A));

endmodule //FA__4_977

module FA__4_981 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_981

module FA__4_985 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_985

module FA__4_989 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_989

module CSAlike__4_1006 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__4_853 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .CIN (C[38]));
FA__4_857 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .CIN (C[37]));
FA__4_861 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36])
    , .CIN (C[36]));
FA__4_865 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__4_869 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__4_873 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__4_877 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__4_881 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__4_885 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__4_889 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__4_893 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__4_897 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__4_901 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__4_905 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__4_909 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__4_913 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__4_917 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__4_921 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__4_925 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__4_929 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__4_933 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__4_937 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]), .CIN (C[17]));
FA__4_941 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16])
    , .CIN (C[16]));
FA__4_945 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]), .CIN (C[15]));
FA__4_949 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]), .CIN (C[14]));
FA__4_953 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]), .CIN (C[13]));
FA__4_957 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12]), .CIN (C[12]));
FA__4_961 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]), .CIN (C[11]));
FA__4_965 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10]), .CIN (C[10]));
FA__4_969 genblk1_9_fa (.COUT (carry[10]), .SUM (result[9]), .A (A[9]), .B (B[9]), .CIN (C[9]));
FA__4_973 genblk1_8_fa (.COUT (carry[9]), .SUM (result[8]), .A (A[8]), .B (B[8]), .CIN (C[8]));
FA__4_977 genblk1_7_fa (.COUT (carry[8]), .SUM (result[7]), .A (A[7]), .B (B[7]), .CIN (C[7]));
FA__4_981 genblk1_6_fa (.COUT (carry[7]), .SUM (result[6]), .A (A[6]), .B (B[6]));
FA__4_985 genblk1_5_fa (.COUT (carry[6]), .SUM (result[5]), .A (A[5]), .B (B[5]));
FA__4_989 genblk1_4_fa (.COUT (carry[5]), .SUM (result[4]), .A (A[4]), .B (B[4]));

endmodule //CSAlike__4_1006

module FA__4_556 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_556

module FA__4_560 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_560

module FA__4_564 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_564

module FA__4_568 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_568

module FA__4_572 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_572

module FA__4_576 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__4_576

module FA__4_580 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_580

module FA__4_584 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__4_584

module FA__4_588 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_588

module FA__4_592 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_opt_ipo_n20;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (CLOCK_opt_ipo_n20), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (CLOCK_opt_ipo_n20), .B (B));
INV_X2 CLOCK_opt_ipo_c5 (.ZN (CLOCK_opt_ipo_n20), .A (A));

endmodule //FA__4_592

module FA__4_596 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_596

module FA__4_600 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_600

module FA__4_604 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_604

module FA__4_608 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n26;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X2 CLOCK_slo__mro_c7 (.ZN (CLOCK_slo__mro_n26), .A (A));
XNOR2_X2 CLOCK_slo__mro_c8 (.ZN (temp), .A (CLOCK_slo__mro_n26), .B (B));

endmodule //FA__4_608

module FA__4_612 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_612

module FA__4_616 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire opt_ipo_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (opt_ipo_n3), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (opt_ipo_n3), .B (B));
INV_X2 opt_ipo_c3 (.ZN (opt_ipo_n3), .A (A));

endmodule //FA__4_616

module FA__4_620 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_620

module FA__4_624 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_624

module FA__4_628 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire opt_ipo_n4;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (opt_ipo_n4), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (opt_ipo_n4), .B (B));
INV_X2 opt_ipo_c2 (.ZN (opt_ipo_n4), .A (A));

endmodule //FA__4_628

module FA__4_632 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_632

module FA__4_636 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__n1), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
XOR2_X2 CLOCK_slo__c1 (.Z (CLOCK_slo__n1), .A (A), .B (B));

endmodule //FA__4_636

module FA__4_640 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_640

module FA__4_644 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (CLOCK_slo__n1), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
XOR2_X1 CLOCK_slo__c1 (.Z (CLOCK_slo__n1), .A (A), .B (B));

endmodule //FA__4_644

module FA__4_648 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_648

module FA__4_652 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_652

module FA__4_656 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire opt_ipo_n25;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (opt_ipo_n25), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (opt_ipo_n25), .B (B));
INV_X2 opt_ipo_c9 (.ZN (opt_ipo_n25), .A (A));

endmodule //FA__4_656

module FA__4_660 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_660

module FA__4_664 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_664

module FA__4_668 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_668

module FA__4_672 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_672

module FA__4_676 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_676

module FA__4_680 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__4_680

module FA__4_684 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_684

module FA__4_688 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_688

module FA__4_692 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_692

module FA__4_696 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_696

module CSAlike__4_753 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__4_556 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .B (B[49]), .CIN (C[49]));
FA__4_560 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .B (B[48]), .CIN (C[48]));
FA__4_564 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .B (B[47]), .CIN (C[47]));
FA__4_568 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .B (B[46]), .CIN (C[46]));
FA__4_572 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .B (B[45]), .CIN (C[45]));
FA__4_576 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .B (B[44]), .CIN (C[44]));
FA__4_580 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__4_584 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__4_588 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__4_592 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40])
    , .CIN (C[40]));
FA__4_596 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__4_600 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38])
    , .CIN (C[38]));
FA__4_604 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__4_608 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36])
    , .CIN (C[36]));
FA__4_612 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__4_616 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__4_620 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33])
    , .CIN (C[33]));
FA__4_624 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__4_628 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__4_632 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__4_636 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__4_640 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__4_644 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__4_648 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__4_652 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__4_656 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24])
    , .CIN (C[24]));
FA__4_660 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__4_664 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__4_668 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__4_672 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__4_676 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__4_680 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__4_684 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]), .CIN (C[17]));
FA__4_688 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16]));
FA__4_692 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]));
FA__4_696 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]));

endmodule //CSAlike__4_753

module FA__4_271 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_271

module FA__4_275 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_275

module FA__4_279 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_279

module FA__4_283 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_283

module FA__4_287 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_287

module FA__4_291 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_291

module FA__4_295 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_295

module FA__4_299 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n7), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c2 (.ZN (SUM), .A (CLOCK_slo__sro_n7), .B (temp));

endmodule //FA__4_299

module FA__4_303 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_303

module FA__4_307 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n1), .A (B));
XNOR2_X2 slo__sro_c2 (.ZN (temp), .A (slo__sro_n1), .B (A));

endmodule //FA__4_307

module FA__4_311 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n5;
wire CLOCK_slo__sro_n6;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n5), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n5), .B (CIN));
INV_X1 CLOCK_slo__sro_c5 (.ZN (CLOCK_slo__sro_n6), .A (A));
XNOR2_X2 CLOCK_slo__sro_c6 (.ZN (CLOCK_slo__sro_n5), .A (CLOCK_slo__sro_n6), .B (B));

endmodule //FA__4_311

module FA__4_315 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_315

module FA__4_319 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__sro_n1;
wire slo__sro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__sro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__sro_n1), .B (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n2), .A (B));
XNOR2_X2 slo__sro_c2 (.ZN (slo__sro_n1), .A (slo__sro_n2), .B (A));

endmodule //FA__4_319

module FA__4_323 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_323

module FA__4_327 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n1), .A (A));
XNOR2_X2 slo__mro_c2 (.ZN (temp), .A (slo__mro_n1), .B (B));

endmodule //FA__4_327

module FA__4_331 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_331

module FA__4_335 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_335

module FA__4_339 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_339

module FA__4_343 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X2 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n3), .A (temp));
XNOR2_X2 CLOCK_slo__sro_c2 (.ZN (SUM), .A (CLOCK_slo__sro_n3), .B (CIN));

endmodule //FA__4_343

module FA__4_347 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_347

module FA__4_351 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_351

module FA__4_355 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_355

module FA__4_359 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__sro_n1;
wire slo__sro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__sro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__sro_n1), .B (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n2), .A (B));
XNOR2_X1 slo__sro_c2 (.ZN (slo__sro_n1), .A (A), .B (slo__sro_n2));

endmodule //FA__4_359

module FA__4_363 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_363

module FA__4_367 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__4_367

module FA__4_371 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_371

module FA__4_375 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n7), .A (CIN));
XNOR2_X2 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n7));

endmodule //FA__4_375

module FA__4_379 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_379

module FA__4_383 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_383

module FA__4_387 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__4_387

module FA__4_391 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__mro_n1;
wire slo__mro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__mro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__mro_n1), .B (CIN));
XNOR2_X2 slo__mro_c1 (.ZN (slo__mro_n2), .A (B), .B (A));
INV_X2 slo__mro_c2 (.ZN (slo__mro_n1), .A (slo__mro_n2));

endmodule //FA__4_391

module FA__4_395 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_395

module FA__4_399 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_399

module FA__4_403 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__4_403

module CSAlike__4_500 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__4_271 genblk1_57_fa (.COUT (carry[58]), .SUM (result[57]), .A (A[57]), .B (B[57]), .CIN (C[57]));
FA__4_275 genblk1_56_fa (.COUT (carry[57]), .SUM (result[56]), .A (A[56]), .B (B[56]), .CIN (C[56]));
FA__4_279 genblk1_55_fa (.COUT (carry[56]), .SUM (result[55]), .A (A[55]), .B (B[55]), .CIN (C[55]));
FA__4_283 genblk1_54_fa (.COUT (carry[55]), .SUM (result[54]), .A (A[54]), .B (B[54]), .CIN (C[54]));
FA__4_287 genblk1_53_fa (.COUT (carry[54]), .SUM (result[53]), .A (A[53]), .B (B[53]), .CIN (C[53]));
FA__4_291 genblk1_52_fa (.COUT (carry[53]), .SUM (result[52]), .A (A[52]), .B (B[52]), .CIN (C[52]));
FA__4_295 genblk1_51_fa (.COUT (carry[52]), .SUM (result[51]), .A (A[51]), .B (B[51]), .CIN (C[51]));
FA__4_299 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .B (B[50]), .CIN (C[50]));
FA__4_303 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .B (B[49])
    , .CIN (C[49]));
FA__4_307 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__4_311 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__4_315 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__4_319 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__4_323 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__4_327 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__4_331 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__4_335 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41])
    , .CIN (C[41]));
FA__4_339 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__4_343 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__4_347 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__4_351 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__4_355 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__4_359 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__4_363 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__4_367 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__4_371 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32])
    , .CIN (C[32]));
FA__4_375 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__4_379 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__4_383 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__4_387 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__4_391 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__4_395 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]));
FA__4_399 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]));
FA__4_403 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]));

endmodule //CSAlike__4_500

module FA__3_143 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__3_143

module FA__3_139 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (CIN));

endmodule //FA__3_139

module FA__3_135 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__3_135

module FA__3_131 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_11 (.ZN (n_0_8), .A (B));
INV_X1 i_0_10 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_9 (.ZN (n_0_6), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X1 i_0_8 (.ZN (n_0_5), .A1 (B), .A2 (A));
AOI21_X1 i_0_7 (.ZN (n_0_4), .A (CIN), .B1 (n_0_6), .B2 (n_0_5));
NAND3_X1 i_0_6 (.ZN (n_0_3), .A1 (n_0_6), .A2 (CIN), .A3 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_2), .A (n_0_3));
NOR2_X1 i_0_4 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_0 (.ZN (temp), .A (n_0_1));
INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));

endmodule //FA__3_131

module FA__3_127 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X1 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (CIN), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (B), .A2 (A));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (B), .A2 (A));

endmodule //FA__3_127

module FA__3_123 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


OR2_X1 i_0_9 (.ZN (n_0_7), .A1 (B), .A2 (CIN));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (B), .A2 (CIN));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (A), .A2 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_3), .A (A));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_5));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_2 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (A), .A2 (n_0_7));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_0), .A2 (n_0_6));

endmodule //FA__3_123

module FA__3_119 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


INV_X1 i_0_9 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (B), .A2 (CIN));
NOR2_X1 i_0_7 (.ZN (n_0_5), .A1 (B), .A2 (CIN));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_6));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_7), .A2 (n_0_2));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (n_0_3));
NAND2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
OAI21_X1 i_0_0 (.ZN (COUT), .A (n_0_6), .B1 (n_0_7), .B2 (n_0_5));

endmodule //FA__3_119

module FA__3_115 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


INV_X1 i_0_9 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (B), .A2 (CIN));
NOR2_X1 i_0_7 (.ZN (n_0_5), .A1 (B), .A2 (CIN));
INV_X1 i_0_6 (.ZN (n_0_4), .A (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_6));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_7), .A2 (n_0_2));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (n_0_3));
NAND2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
OAI21_X1 i_0_0 (.ZN (COUT), .A (n_0_6), .B1 (n_0_7), .B2 (n_0_5));

endmodule //FA__3_115

module FA__3_111 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n1), .A (B));
XNOR2_X1 CLOCK_slo__mro_c2 (.ZN (temp), .A (A), .B (CLOCK_slo__mro_n1));

endmodule //FA__3_111

module FA__3_107 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__n13;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__n13), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));
XOR2_X1 slo__c5 (.Z (slo__n13), .A (B), .B (A));

endmodule //FA__3_107

module FA__3_103 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_103

module FA__3_99 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n35;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X2 CLOCK_slo__mro_c14 (.ZN (CLOCK_slo__mro_n35), .A (A));
XNOR2_X2 CLOCK_slo__mro_c15 (.ZN (temp), .A (CLOCK_slo__mro_n35), .B (B));

endmodule //FA__3_99

module FA__3_95 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_95

module FA__3_91 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


INV_X1 i_0_9 (.ZN (n_0_7), .A (CIN));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_1), .A2 (n_0_2));
AOI21_X1 i_0_7 (.ZN (n_0_5), .A (n_0_7), .B1 (A), .B2 (B));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (A), .A2 (B));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_6), .A2 (n_0_4));
AOI22_X1 i_0_4 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_7), .B1 (n_0_6), .B2 (n_0_5));
INV_X1 i_0_3 (.ZN (n_0_2), .A (B));
INV_X1 i_0_2 (.ZN (n_0_1), .A (A));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
AOI21_X1 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_1));

endmodule //FA__3_91

module FA__3_87 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_87

module FA__3_83 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_83

module FA__3_79 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;


AOI22_X1 i_0_2 (.ZN (COUT), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__3_79

module FA__3_75 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X2 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__3_75

module FA__3_71 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__sro_n6;
wire slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CIN), .B2 (slo__sro_n6));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__sro_n6), .B (CIN));
INV_X2 slo__sro_c4 (.ZN (slo__sro_n7), .A (B));
XNOR2_X2 slo__sro_c5 (.ZN (slo__sro_n6), .A (A), .B (slo__sro_n7));

endmodule //FA__3_71

module FA__3_67 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__3_67

module FA__3_63 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__n75;
wire temp;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire slo__n29;
wire CLOCK_slo__sro_n69;
wire opt_ipo_n44;


INV_X1 i_0_11 (.ZN (n_0_8), .A (B));
INV_X2 i_0_10 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_9 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
AOI22_X1 CLOCK_slo__sro_c57 (.ZN (CLOCK_slo__sro_n69), .A1 (temp), .A2 (CIN), .B1 (B), .B2 (A));
AOI21_X4 i_0_7 (.ZN (n_0_4), .A (CIN), .B1 (n_0_6), .B2 (n_0_5));
NAND3_X2 i_0_6 (.ZN (n_0_3), .A1 (CLOCK_slo__n75), .A2 (CIN), .A3 (n_0_5));
NOR2_X4 i_0_4 (.ZN (SUM), .A1 (n_0_4), .A2 (opt_ipo_n44));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (slo__n29), .A2 (n_0_5));
INV_X1 i_0_0 (.ZN (temp), .A (n_0_1));
INV_X2 i_0_3 (.ZN (COUT), .A (CLOCK_slo__sro_n69));
NAND2_X1 CLOCK_slo__c63 (.ZN (CLOCK_slo__n75), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 slo__c28 (.ZN (slo__n29), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X2 CLOCK_slo__sro_c49 (.ZN (n_0_5), .A1 (B), .A2 (A));
INV_X2 opt_ipo_c41 (.ZN (opt_ipo_n44), .A (n_0_3));

endmodule //FA__3_63

module FA__3_59 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire CLOCK_sgo__sro_n5;


AND2_X1 CLOCK_sgo__sro_c2 (.ZN (CLOCK_sgo__sro_n5), .A1 (B), .A2 (A));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AOI21_X2 CLOCK_sgo__sro_c3 (.ZN (COUT), .A (CLOCK_sgo__sro_n5), .B1 (temp), .B2 (CIN));

endmodule //FA__3_59

module FA__3_55 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X1 i_0_8 (.ZN (SUM), .A1 (n_0_5), .A2 (n_0_6));
AOI21_X1 i_0_7 (.ZN (n_0_6), .A (A), .B1 (n_0_3), .B2 (n_0_4));
AND3_X1 i_0_6 (.ZN (n_0_5), .A1 (A), .A2 (n_0_3), .A3 (n_0_4));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (CIN), .A2 (B));
OR2_X2 i_0_4 (.ZN (n_0_3), .A1 (CIN), .A2 (B));
INV_X1 i_0_3 (.ZN (n_0_2), .A (B));
INV_X1 i_0_2 (.ZN (n_0_1), .A (A));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
AOI21_X2 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_1));

endmodule //FA__3_55

module FA__3_51 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


NOR2_X1 i_0_9 (.ZN (n_0_7), .A1 (A), .A2 (B));
INV_X1 i_0_8 (.ZN (n_0_6), .A (n_0_7));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (A), .A2 (B));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (CIN), .A2 (n_0_4));
INV_X1 i_0_4 (.ZN (n_0_2), .A (CIN));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_4));
NAND2_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1));
NAND2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_0), .A2 (n_0_3));
AOI21_X1 i_0_0 (.ZN (COUT), .A (n_0_7), .B1 (n_0_2), .B2 (n_0_5));

endmodule //FA__3_51

module FA__3_47 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X2 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X2 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (CIN), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__3_47

module FA__3_43 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


OR2_X2 i_0_12 (.ZN (n_0_10), .A1 (B), .A2 (A));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (B), .A2 (A));
NAND2_X2 i_0_10 (.ZN (n_0_8), .A1 (n_0_10), .A2 (n_0_9));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (CIN), .A2 (n_0_8));
INV_X1 i_0_8 (.ZN (n_0_6), .A (CIN));
INV_X1 i_0_7 (.ZN (n_0_5), .A (n_0_8));
NAND2_X2 i_0_6 (.ZN (n_0_4), .A1 (n_0_6), .A2 (n_0_5));
NAND2_X2 i_0_5 (.ZN (SUM), .A1 (n_0_4), .A2 (n_0_7));
INV_X1 i_0_2 (.ZN (n_0_1), .A (n_0_9));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (n_0_1), .B1 (CIN), .B2 (n_0_10));
INV_X1 i_0_0 (.ZN (COUT), .A (n_0_0));

endmodule //FA__3_43

module FA__3_39 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NOR2_X2 i_0_8 (.ZN (SUM), .A1 (n_0_5), .A2 (n_0_6));
AOI21_X2 i_0_7 (.ZN (n_0_6), .A (A), .B1 (n_0_3), .B2 (n_0_4));
AND3_X1 i_0_6 (.ZN (n_0_5), .A1 (n_0_3), .A2 (A), .A3 (n_0_4));
NAND2_X1 i_0_5 (.ZN (n_0_4), .A1 (CIN), .A2 (B));
OR2_X2 i_0_4 (.ZN (n_0_3), .A1 (CIN), .A2 (B));
OAI21_X1 i_0_3 (.ZN (COUT), .A (n_0_0), .B1 (n_0_1), .B2 (n_0_2));
INV_X1 i_0_2 (.ZN (n_0_2), .A (A));
INV_X1 i_0_1 (.ZN (n_0_1), .A (B));
OAI21_X1 i_0_0 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));

endmodule //FA__3_39

module FA__3_35 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


NOR2_X1 i_0_10 (.ZN (n_0_8), .A1 (A), .A2 (B));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (A), .A2 (B));
INV_X1 i_0_8 (.ZN (n_0_6), .A (n_0_7));
OAI21_X1 i_0_7 (.ZN (n_0_5), .A (CIN), .B1 (n_0_6), .B2 (n_0_8));
INV_X1 i_0_6 (.ZN (n_0_4), .A (CIN));
INV_X1 i_0_5 (.ZN (n_0_3), .A (B));
INV_X1 i_0_4 (.ZN (n_0_2), .A (A));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (n_0_3));
NAND3_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_1), .A2 (n_0_4), .A3 (n_0_7));
NAND2_X2 i_0_1 (.ZN (SUM), .A1 (n_0_5), .A2 (n_0_0));
OAI21_X1 i_0_0 (.ZN (COUT), .A (n_0_7), .B1 (n_0_8), .B2 (n_0_4));

endmodule //FA__3_35

module FA__3_31 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__n5;
wire temp;


XOR2_X1 CLOCK_slo__c4 (.Z (CLOCK_slo__n5), .A (A), .B (B));
AOI22_X1 i_0_2 (.ZN (COUT), .A1 (A), .A2 (B), .B1 (CLOCK_slo__n5), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_31

module FA__3_27 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__sro_n16;
wire sgo__sro_n7;
wire sgo__sro_n8;
wire CLOCK_slo__sro_n17;


INV_X2 i_0_3 (.ZN (COUT), .A (sgo__sro_n7));
INV_X1 CLOCK_slo__sro_c10 (.ZN (CLOCK_slo__sro_n17), .A (A));
XOR2_X1 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n16), .B (CIN));
AND2_X1 sgo__sro_c3 (.ZN (sgo__sro_n8), .A1 (B), .A2 (A));
AOI21_X2 sgo__sro_c4 (.ZN (sgo__sro_n7), .A (sgo__sro_n8), .B1 (CLOCK_slo__sro_n16), .B2 (CIN));
XNOR2_X2 CLOCK_slo__sro_c11 (.ZN (CLOCK_slo__sro_n16), .A (B), .B (CLOCK_slo__sro_n17));

endmodule //FA__3_27

module FA__3_23 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_23

module FA__3_19 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__3_19

module FA__3_15 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__3_15

module CSAlike__0_118 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__3_143 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .CIN (C[35]));
FA__3_139 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .CIN (C[34]));
FA__3_135 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__3_131 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__3_127 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__3_123 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__3_119 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__3_115 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__3_111 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__3_107 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__3_103 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__3_99 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24])
    , .CIN (C[24]));
FA__3_95 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__3_91 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__3_87 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__3_83 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__3_79 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__3_75 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__3_71 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17])
    , .CIN (C[17]));
FA__3_67 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16]), .CIN (C[16]));
FA__3_63 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]), .CIN (C[15]));
FA__3_59 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]), .CIN (C[14]));
FA__3_55 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]), .CIN (C[13]));
FA__3_51 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12]), .CIN (C[12]));
FA__3_47 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]), .CIN (C[11]));
FA__3_43 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10]), .CIN (C[10]));
FA__3_39 genblk1_9_fa (.COUT (carry[10]), .SUM (result[9]), .A (A[9]), .B (B[9]), .CIN (C[9]));
FA__3_35 genblk1_8_fa (.COUT (carry[9]), .SUM (result[8]), .A (A[8]), .B (B[8]), .CIN (C[8]));
FA__3_31 genblk1_7_fa (.COUT (carry[8]), .SUM (result[7]), .A (A[7]), .B (B[7]), .CIN (C[7]));
FA__3_27 genblk1_6_fa (.COUT (carry[7]), .SUM (result[6]), .A (A[6]), .B (B[6]), .CIN (C[6]));
FA__3_23 genblk1_5_fa (.COUT (carry[6]), .SUM (result[5]), .A (A[5]), .B (B[5]), .CIN (C[5]));
FA__3_19 genblk1_4_fa (.COUT (carry[5]), .SUM (result[4]), .A (A[4]), .B (B[4]));
FA__3_15 genblk1_3_fa (.COUT (carry[4]), .SUM (result[3]), .A (A[3]), .B (B[3]));

endmodule //CSAlike__0_118

module FA__3_1090 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__3_1090

module FA__3_1094 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__3_1094

module FA__3_1098 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__3_1098

module FA__3_1102 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__sro_n7;
wire CLOCK_slo__sro_n8;


INV_X2 CLOCK_slo__sro_c6 (.ZN (CLOCK_slo__sro_n8), .A (A));
AOI22_X1 i_0_2 (.ZN (COUT), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n7), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n7), .B (CIN));
XNOR2_X2 CLOCK_slo__sro_c7 (.ZN (CLOCK_slo__sro_n7), .A (B), .B (CLOCK_slo__sro_n8));

endmodule //FA__3_1102

module FA__3_1106 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1106

module FA__3_1110 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire sgo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X1 sgo__sro_c3 (.ZN (sgo__sro_n7), .A1 (B), .A2 (A));
AOI21_X1 sgo__sro_c4 (.ZN (n_0_0), .A (sgo__sro_n7), .B1 (temp), .B2 (CIN));

endmodule //FA__3_1110

module FA__3_1114 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n3;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n3), .A (CIN));
XNOR2_X2 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n3));

endmodule //FA__3_1114

module FA__3_1118 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1118

module FA__3_1122 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1122

module FA__3_1126 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;


AOI22_X1 i_0_2 (.ZN (COUT), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1126

module FA__3_1130 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__mro_n10;
wire slo__mro_n11;
wire CLOCK_slo__sro_n22;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__mro_n10), .B2 (CIN));
INV_X1 CLOCK_slo__sro_c17 (.ZN (CLOCK_slo__sro_n22), .A (CIN));
INV_X1 slo__mro_c7 (.ZN (slo__mro_n11), .A (A));
XNOR2_X2 slo__mro_c8 (.ZN (slo__mro_n10), .A (slo__mro_n11), .B (B));
XNOR2_X1 CLOCK_slo__sro_c18 (.ZN (SUM), .A (slo__mro_n10), .B (CLOCK_slo__sro_n22));

endmodule //FA__3_1130

module FA__3_1134 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__sro_n19;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n3;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AND2_X2 CLOCK_slo__sro_c10 (.ZN (CLOCK_slo__sro_n19), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n3), .A (CIN));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n3));
AOI21_X1 CLOCK_slo__sro_c11 (.ZN (n_0_0), .A (CLOCK_slo__sro_n19), .B1 (temp), .B2 (CIN));

endmodule //FA__3_1134

module FA__3_1138 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;


AOI22_X2 i_0_2 (.ZN (COUT), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1138

module FA__3_1142 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1142

module FA__3_1146 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n6;
wire CLOCK_slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
XOR2_X1 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n6), .B (CIN));
AOI22_X2 CLOCK_slo__sro_c12 (.ZN (n_0_0), .A1 (CLOCK_slo__sro_n6), .A2 (CIN), .B1 (A), .B2 (B));
INV_X2 CLOCK_slo__sro_c4 (.ZN (CLOCK_slo__sro_n7), .A (A));
XNOR2_X2 CLOCK_slo__sro_c5 (.ZN (CLOCK_slo__sro_n6), .A (B), .B (CLOCK_slo__sro_n7));

endmodule //FA__3_1146

module FA__3_1150 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1150

module FA__3_1154 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1154

module FA__3_1158 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1158

module FA__3_1162 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1162

module FA__3_1166 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;


AOI22_X1 i_0_2 (.ZN (COUT), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__3_1166

module FA__3_1170 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1170

module FA__3_1174 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1174

module FA__3_1178 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1178

module FA__3_1182 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1182

module FA__3_1186 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1186

module FA__3_1190 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n1;
wire CLOCK_slo__sro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n1), .B (CIN));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n2), .A (B));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (CLOCK_slo__sro_n1), .A (CLOCK_slo__sro_n2), .B (A));

endmodule //FA__3_1190

module FA__3_1194 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_1194

module FA__3_1198 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n3), .A (CIN));
XNOR2_X2 slo__mro_c2 (.ZN (SUM), .A (temp), .B (slo__mro_n3));

endmodule //FA__3_1198

module FA__3_1202 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo___n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo___n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
CLKBUF_X1 slo___L1_c1 (.Z (slo___n1), .A (temp));

endmodule //FA__3_1202

module FA__3_1206 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_11 (.ZN (n_0_8), .A (B));
INV_X1 i_0_10 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_9 (.ZN (n_0_6), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X1 i_0_8 (.ZN (n_0_5), .A1 (B), .A2 (A));
AOI21_X1 i_0_7 (.ZN (n_0_4), .A (CIN), .B1 (n_0_6), .B2 (n_0_5));
NAND3_X1 i_0_6 (.ZN (n_0_3), .A1 (n_0_6), .A2 (CIN), .A3 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_2), .A (n_0_3));
NOR2_X1 i_0_4 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_0 (.ZN (temp), .A (n_0_1));
INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));

endmodule //FA__3_1206

module FA__3_1210 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;


NAND2_X1 i_0_13 (.ZN (n_0_10), .A1 (B), .A2 (A));
INV_X1 i_0_12 (.ZN (n_0_9), .A (n_0_10));
NOR2_X1 i_0_11 (.ZN (n_0_8), .A1 (B), .A2 (A));
OAI21_X1 i_0_10 (.ZN (n_0_7), .A (CIN), .B1 (n_0_9), .B2 (n_0_8));
INV_X1 i_0_9 (.ZN (n_0_6), .A (CIN));
INV_X1 i_0_8 (.ZN (n_0_5), .A (B));
INV_X1 i_0_7 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND3_X1 i_0_5 (.ZN (n_0_2), .A1 (n_0_3), .A2 (n_0_6), .A3 (n_0_10));
NAND2_X1 i_0_4 (.ZN (SUM), .A1 (n_0_7), .A2 (n_0_2));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_10));
INV_X1 i_0_0 (.ZN (temp), .A (n_0_1));
INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));

endmodule //FA__3_1210

module FA__3_1214 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__3_1214

module FA__3_1218 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__3_1218

module FA__3_1222 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__3_1222

module CSAlike__3_1259 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__3_1090 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .B (B[42]), .CIN (C[42]));
FA__3_1094 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .B (B[41]), .CIN (C[41]));
FA__3_1098 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .B (B[40]), .CIN (C[40]));
FA__3_1102 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__3_1106 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__3_1110 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__3_1114 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__3_1118 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35])
    , .CIN (C[35]));
FA__3_1122 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__3_1126 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__3_1130 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__3_1134 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__3_1138 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__3_1142 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__3_1146 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__3_1150 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__3_1154 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__3_1158 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__3_1162 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__3_1166 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23])
    , .CIN (C[23]));
FA__3_1170 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__3_1174 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__3_1178 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__3_1182 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__3_1186 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__3_1190 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]), .CIN (C[17]));
FA__3_1194 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16])
    , .CIN (C[16]));
FA__3_1198 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]), .CIN (C[15]));
FA__3_1202 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]), .CIN (C[14]));
FA__3_1206 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]), .CIN (C[13]));
FA__3_1210 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12]), .CIN (C[12]));
FA__3_1214 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]));
FA__3_1218 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10]));
FA__3_1222 genblk1_9_fa (.COUT (carry[10]), .SUM (result[9]), .A (A[9]), .B (B[9]));

endmodule //CSAlike__3_1259

module FA__3_813 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__3_813

module FA__3_817 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_817

module FA__3_821 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_821

module FA__3_825 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_825

module FA__3_829 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_829

module FA__3_833 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire spw_n30;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (spw_n30), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));
CLKBUF_X1 spw__L1_c1_c23 (.Z (spw_n30), .A (A));

endmodule //FA__3_833

module FA__3_837 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__3_837

module FA__3_841 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_841

module FA__3_845 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n7), .A (CIN));
XNOR2_X1 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n7));

endmodule //FA__3_845

module FA__3_849 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_849

module FA__3_853 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n11;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c5 (.ZN (CLOCK_slo__sro_n11), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c6 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n11));

endmodule //FA__3_853

module FA__3_857 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_857

module FA__3_861 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n7;
wire CLOCK_slo__sro_n16;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n7), .A (CIN));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n7));
INV_X1 CLOCK_slo__sro_c9 (.ZN (CLOCK_slo__sro_n16), .A (B));
XNOR2_X1 CLOCK_slo__sro_c10 (.ZN (temp), .A (CLOCK_slo__sro_n16), .B (A));

endmodule //FA__3_861

module FA__3_865 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_865

module FA__3_869 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_869

module FA__3_873 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n5;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));
INV_X2 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n5), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n5));

endmodule //FA__3_873

module FA__3_877 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__3_877

module FA__3_881 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n3), .A (CIN));
XNOR2_X2 slo__mro_c2 (.ZN (SUM), .A (temp), .B (slo__mro_n3));

endmodule //FA__3_881

module FA__3_885 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_885

module FA__3_889 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_889

module FA__3_893 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n3), .A (CIN));
XNOR2_X1 CLOCK_slo__mro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__mro_n3));

endmodule //FA__3_893

module FA__3_897 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_897

module FA__3_901 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n3), .A (CIN));
XNOR2_X2 slo__mro_c2 (.ZN (SUM), .A (temp), .B (slo__mro_n3));

endmodule //FA__3_901

module FA__3_905 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_905

module FA__3_909 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n7), .A (CIN));
XNOR2_X1 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n7));

endmodule //FA__3_909

module FA__3_913 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_913

module FA__3_917 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_917

module FA__3_921 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_921

module FA__3_925 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_925

module FA__3_929 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_929

module FA__3_933 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n3), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n3));

endmodule //FA__3_933

module FA__3_937 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X2 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__3_937

module FA__3_941 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__3_941

module CSAlike__3_1006 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__3_813 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .B (B[48]), .CIN (C[48]));
FA__3_817 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__3_821 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__3_825 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__3_829 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__3_833 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__3_837 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__3_841 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__3_845 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__3_849 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__3_853 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__3_857 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__3_861 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__3_865 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__3_869 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__3_873 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__3_877 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__3_881 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__3_885 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__3_889 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__3_893 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__3_897 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__3_901 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__3_905 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25])
    , .CIN (C[25]));
FA__3_909 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__3_913 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__3_917 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__3_921 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__3_925 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__3_929 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__3_933 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__3_937 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]));
FA__3_941 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16]));

endmodule //CSAlike__3_1006

module FA__3_528 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__3_528

module FA__3_532 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__3_532

module FA__3_536 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__3_536

module FA__3_540 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__3_540

module FA__3_544 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__3_544

module FA__3_548 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_548

module FA__3_552 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_552

module FA__3_556 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n5;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n5), .A (CIN));
XNOR2_X2 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n5));

endmodule //FA__3_556

module FA__3_560 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire CLOCK_sgo__sro_n9;
wire CLOCK_sgo__sro_n10;
wire CLOCK_sgo__sro_n11;


INV_X2 i_0_3 (.ZN (COUT), .A (CLOCK_sgo__sro_n9));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
NAND2_X1 CLOCK_sgo__sro_c5 (.ZN (CLOCK_sgo__sro_n11), .A1 (B), .A2 (A));
INV_X1 CLOCK_sgo__sro_c6 (.ZN (CLOCK_sgo__sro_n10), .A (CLOCK_sgo__sro_n11));
AOI21_X1 CLOCK_sgo__sro_c7 (.ZN (CLOCK_sgo__sro_n9), .A (CLOCK_sgo__sro_n10), .B1 (temp), .B2 (CIN));

endmodule //FA__3_560

module FA__3_564 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__mro_n1;
wire CLOCK_slo__mro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__mro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__mro_n1), .B (CIN));
INV_X2 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n2), .A (B));
XNOR2_X2 CLOCK_slo__mro_c2 (.ZN (CLOCK_slo__mro_n1), .A (CLOCK_slo__mro_n2), .B (A));

endmodule //FA__3_564

module FA__3_568 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_568

module FA__3_572 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n1), .A (A));
XNOR2_X2 CLOCK_slo__mro_c2 (.ZN (temp), .A (CLOCK_slo__mro_n1), .B (B));

endmodule //FA__3_572

module FA__3_576 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_576

module FA__3_580 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_580

module FA__3_584 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_584

module FA__3_588 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X2 slo__mro_c3 (.ZN (slo__mro_n7), .A (A));
XNOR2_X2 slo__mro_c4 (.ZN (temp), .A (slo__mro_n7), .B (B));

endmodule //FA__3_588

module FA__3_592 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_592

module FA__3_596 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n1), .A (A));
XNOR2_X2 slo__mro_c2 (.ZN (temp), .A (slo__mro_n1), .B (B));

endmodule //FA__3_596

module FA__3_600 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_600

module FA__3_604 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_604

module FA__3_608 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_608

module FA__3_612 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_612

module FA__3_616 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n1), .A (A));
XNOR2_X2 slo__sro_c2 (.ZN (temp), .A (B), .B (slo__sro_n1));

endmodule //FA__3_616

module FA__3_620 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_620

module FA__3_624 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n24;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c9 (.ZN (CLOCK_slo__sro_n24), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c10 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n24));

endmodule //FA__3_624

module FA__3_628 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__n1;
wire opt_ipo_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (opt_ipo_n7), .A2 (B), .B1 (slo__n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (opt_ipo_n7), .B (B));
XOR2_X1 slo__c1 (.Z (slo__n1), .A (opt_ipo_n7), .B (B));
INV_X2 opt_ipo_c5 (.ZN (opt_ipo_n7), .A (A));

endmodule //FA__3_628

module FA__3_632 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_632

module FA__3_636 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n4;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 slo__sro_c4 (.ZN (slo__sro_n4), .A (B));
XNOR2_X2 slo__sro_c5 (.ZN (temp), .A (slo__sro_n4), .B (A));

endmodule //FA__3_636

module FA__3_640 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n3), .A (CIN));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n3));

endmodule //FA__3_640

module FA__3_644 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_644

module FA__3_648 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__n15;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__n15), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
XOR2_X1 CLOCK_slo__c8 (.Z (CLOCK_slo__n15), .A (A), .B (B));

endmodule //FA__3_648

module FA__3_652 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_652

module FA__3_656 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__3_656

module FA__3_660 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__3_660

module CSAlike__3_753 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__3_528 genblk1_56_fa (.COUT (carry[57]), .SUM (result[56]), .B (B[56]), .CIN (C[56]));
FA__3_532 genblk1_55_fa (.COUT (carry[56]), .SUM (result[55]), .B (B[55]), .CIN (C[55]));
FA__3_536 genblk1_54_fa (.COUT (carry[55]), .SUM (result[54]), .B (B[54]), .CIN (C[54]));
FA__3_540 genblk1_53_fa (.COUT (carry[54]), .SUM (result[53]), .B (B[53]), .CIN (C[53]));
FA__3_544 genblk1_52_fa (.COUT (carry[53]), .SUM (result[52]), .B (B[52]), .CIN (C[52]));
FA__3_548 genblk1_51_fa (.COUT (carry[52]), .SUM (result[51]), .A (A[51]), .B (B[51]), .CIN (C[51]));
FA__3_552 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .B (B[50]), .CIN (C[50]));
FA__3_556 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .B (B[49])
    , .CIN (C[49]));
FA__3_560 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__3_564 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__3_568 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__3_572 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__3_576 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__3_580 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__3_584 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__3_588 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41])
    , .CIN (C[41]));
FA__3_592 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__3_596 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__3_600 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__3_604 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__3_608 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__3_612 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__3_616 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__3_620 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__3_624 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32])
    , .CIN (C[32]));
FA__3_628 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__3_632 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__3_636 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__3_640 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__3_644 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__3_648 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__3_652 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__3_656 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]));
FA__3_660 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]));

endmodule //CSAlike__3_753

module FA__3_259 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_259

module FA__3_263 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_263

module FA__3_267 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_267

module FA__3_271 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_271

module FA__3_275 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_275

module FA__3_279 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_279

module FA__3_283 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_283

module FA__3_287 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_287

module FA__3_291 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_291

module FA__3_295 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_295

module FA__3_299 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_299

module FA__3_303 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_303

module FA__3_307 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_307

module FA__3_311 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_311

module FA__3_315 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_315

module FA__3_319 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_319

module FA__3_323 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_323

module FA__3_327 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_327

module FA__3_331 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_331

module FA__3_335 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_335

module FA__3_339 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_339

module FA__3_343 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_343

module FA__3_347 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_347

module FA__3_351 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_351

module FA__3_355 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_355

module FA__3_359 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_359

module FA__3_363 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_363

module FA__3_367 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_367

module FA__3_371 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_371

module FA__3_375 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__3_375

module FA__3_379 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__3_379

module CSAlike__3_500 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__3_259 genblk1_60_fa (.COUT (carry[61]), .SUM (result[60]), .A (A[60]), .B (B[60]), .CIN (C[60]));
FA__3_263 genblk1_59_fa (.COUT (carry[60]), .SUM (result[59]), .A (A[59]), .B (B[59]), .CIN (C[59]));
FA__3_267 genblk1_58_fa (.COUT (carry[59]), .SUM (result[58]), .A (A[58]), .B (B[58]), .CIN (C[58]));
FA__3_271 genblk1_57_fa (.COUT (carry[58]), .SUM (result[57]), .A (A[57]), .B (B[57]), .CIN (C[57]));
FA__3_275 genblk1_56_fa (.COUT (carry[57]), .SUM (result[56]), .A (A[56]), .B (B[56]), .CIN (C[56]));
FA__3_279 genblk1_55_fa (.COUT (carry[56]), .SUM (result[55]), .A (A[55]), .B (B[55]), .CIN (C[55]));
FA__3_283 genblk1_54_fa (.COUT (carry[55]), .SUM (result[54]), .A (A[54]), .B (B[54]), .CIN (C[54]));
FA__3_287 genblk1_53_fa (.COUT (carry[54]), .SUM (result[53]), .A (A[53]), .B (B[53]), .CIN (C[53]));
FA__3_291 genblk1_52_fa (.COUT (carry[53]), .SUM (result[52]), .A (A[52]), .B (B[52]), .CIN (C[52]));
FA__3_295 genblk1_51_fa (.COUT (carry[52]), .SUM (result[51]), .A (A[51]), .B (B[51]), .CIN (C[51]));
FA__3_299 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .B (B[50]), .CIN (C[50]));
FA__3_303 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .B (B[49]), .CIN (C[49]));
FA__3_307 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__3_311 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47])
    , .CIN (C[47]));
FA__3_315 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__3_319 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__3_323 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__3_327 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__3_331 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__3_335 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__3_339 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__3_343 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__3_347 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__3_351 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__3_355 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__3_359 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__3_363 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__3_367 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__3_371 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__3_375 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__3_379 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]));

endmodule //CSAlike__3_500

module FA__2_131 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_131

module FA__2_127 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (B), .A2 (A));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__2_127

module FA__2_123 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X1 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (CIN), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__2_123

module FA__2_119 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X1 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (CIN), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__2_119

module FA__2_115 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_115

module FA__2_111 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_111

module FA__2_107 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X2 CLOCK_slo__sro_c3 (.ZN (CLOCK_slo__sro_n3), .A (B));
XNOR2_X2 CLOCK_slo__sro_c4 (.ZN (temp), .A (A), .B (CLOCK_slo__sro_n3));

endmodule //FA__2_107

module FA__2_103 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__2_103

module FA__2_99 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n13;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c5 (.ZN (CLOCK_slo__sro_n13), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c6 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n13));

endmodule //FA__2_99

module FA__2_95 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n12;
wire CLOCK_slo__sro_n13;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n12), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n12), .B (CIN));
INV_X1 CLOCK_slo__sro_c6 (.ZN (CLOCK_slo__sro_n13), .A (A));
XNOR2_X1 CLOCK_slo__sro_c7 (.ZN (CLOCK_slo__sro_n12), .A (CLOCK_slo__sro_n13), .B (B));

endmodule //FA__2_95

module FA__2_91 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;


NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (A), .A2 (B));
INV_X1 i_0_8 (.ZN (n_0_6), .A (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (A));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_6));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (CIN), .A3 (n_0_7));
INV_X1 i_0_4 (.ZN (n_0_2), .A (n_0_3));
AOI21_X1 i_0_3 (.ZN (n_0_1), .A (CIN), .B1 (n_0_4), .B2 (n_0_7));
NOR2_X1 i_0_2 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_1));
AOI21_X1 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
AOI21_X1 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_6), .B2 (n_0_5));

endmodule //FA__2_91

module FA__2_87 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_87

module FA__2_83 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__2_83

module FA__2_79 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_79

module FA__2_75 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__2_75

module FA__2_71 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo___n37;
wire CLOCK_slo__mro_n53;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo___n37), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
CLKBUF_X1 CLOCK_slo___L1_c37 (.Z (CLOCK_slo___n37), .A (temp));
INV_X2 CLOCK_slo__mro_c49 (.ZN (CLOCK_slo__mro_n53), .A (B));
XNOR2_X2 CLOCK_slo__mro_c50 (.ZN (temp), .A (CLOCK_slo__mro_n53), .B (A));

endmodule //FA__2_71

module FA__2_67 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__n29;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__n29), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
XOR2_X1 CLOCK_slo__c16 (.Z (CLOCK_slo__n29), .A (A), .B (B));

endmodule //FA__2_67

module FA__2_63 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__n10;
wire CLOCK_slo__sro_n23;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));
XOR2_X1 slo__c3 (.Z (slo__n10), .A (B), .B (A));
INV_X1 CLOCK_slo__sro_c13 (.ZN (CLOCK_slo__sro_n23), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c14 (.ZN (SUM), .A (CLOCK_slo__sro_n23), .B (slo__n10));

endmodule //FA__2_63

module FA__2_59 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire slo__mro_n10;
wire temp;
wire slo__mro_n3;
wire slo__sro_n22;


INV_X2 i_0_3 (.ZN (COUT), .A (slo__sro_n22));
INV_X1 slo__mro_c7 (.ZN (slo__mro_n10), .A (A));
AOI22_X1 slo__sro_c17 (.ZN (slo__sro_n22), .A1 (temp), .A2 (CIN), .B1 (B), .B2 (A));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n3), .A (CIN));
XNOR2_X2 slo__mro_c2 (.ZN (SUM), .A (slo__mro_n3), .B (temp));
XNOR2_X1 slo__mro_c8 (.ZN (temp), .A (slo__mro_n10), .B (B));

endmodule //FA__2_59

module FA__2_55 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (n_0_1), .A2 (n_0_2));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (A), .A2 (B));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (CIN));
INV_X1 i_0_6 (.ZN (n_0_4), .A (CIN));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (n_0_4), .A3 (n_0_7));
NAND2_X1 i_0_4 (.ZN (SUM), .A1 (n_0_5), .A2 (n_0_3));
INV_X1 i_0_3 (.ZN (n_0_2), .A (B));
INV_X1 i_0_2 (.ZN (n_0_1), .A (A));
AOI21_X2 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
AOI21_X2 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_1));

endmodule //FA__2_55

module FA__2_51 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__2_51

module FA__2_47 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X1 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (CIN), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__2_47

module FA__2_43 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X1 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (CIN), .A2 (n_0_0), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__2_43

module FA__2_39 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire slo__n1;
wire opt_ipo_n7;


NOR2_X1 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X2 i_0_2 (.ZN (n_0_2), .A1 (CIN), .A2 (n_0_0), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (opt_ipo_n7));
NOR2_X2 slo__c1 (.ZN (slo__n1), .A1 (opt_ipo_n7), .A2 (A));
INV_X2 slo__c3 (.ZN (n_0_0), .A (slo__n1));
INV_X2 opt_ipo_c13 (.ZN (opt_ipo_n7), .A (B));

endmodule //FA__2_39

module FA__2_35 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (B), .A2 (A));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__2_35

module FA__2_31 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NOR2_X1 i_0_5 (.ZN (n_0_2), .A1 (A), .A2 (B));
AOI21_X1 i_0_4 (.ZN (n_0_1), .A (CIN), .B1 (A), .B2 (B));
NOR2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_1), .A2 (n_0_2));
XNOR2_X1 i_0_2 (.ZN (n_0_0), .A (A), .B (B));
INV_X2 i_0_0 (.ZN (temp), .A (n_0_0));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));

endmodule //FA__2_31

module FA__2_27 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__2_27

module FA__2_23 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_23

module FA__2_19 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_19

module FA__2_15 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_15

module FA__2_11 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__2_11

module CSAlike__0_113 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__2_131 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__2_127 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__2_123 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__2_119 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__2_115 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__2_111 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__2_107 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__2_103 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__2_99 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__2_95 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__2_91 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__2_87 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__2_83 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__2_79 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19])
    , .CIN (C[19]));
FA__2_75 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__2_71 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17])
    , .CIN (C[17]));
FA__2_67 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16]), .CIN (C[16]));
FA__2_63 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15])
    , .CIN (C[15]));
FA__2_59 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]), .CIN (C[14]));
FA__2_55 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]), .CIN (C[13]));
FA__2_51 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12]), .CIN (C[12]));
FA__2_47 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]), .CIN (C[11]));
FA__2_43 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10]), .CIN (C[10]));
FA__2_39 genblk1_9_fa (.COUT (carry[10]), .SUM (result[9]), .A (A[9]), .B (B[9]), .CIN (C[9]));
FA__2_35 genblk1_8_fa (.COUT (carry[9]), .SUM (result[8]), .A (A[8]), .B (B[8]), .CIN (C[8]));
FA__2_31 genblk1_7_fa (.COUT (carry[8]), .SUM (result[7]), .A (A[7]), .B (B[7]), .CIN (C[7]));
FA__2_27 genblk1_6_fa (.COUT (carry[7]), .SUM (result[6]), .A (A[6]), .B (B[6]), .CIN (C[6]));
FA__2_23 genblk1_5_fa (.COUT (carry[6]), .SUM (result[5]), .A (A[5]), .B (B[5]), .CIN (C[5]));
FA__2_19 genblk1_4_fa (.COUT (carry[5]), .SUM (result[4]), .A (A[4]), .B (B[4]), .CIN (C[4]));
FA__2_15 genblk1_3_fa (.COUT (carry[4]), .SUM (result[3]), .A (A[3]), .B (B[3]), .CIN (C[3]));
FA__2_11 genblk1_2_fa (.COUT (carry[3]), .SUM (result[2]), .A (A[2]), .B (B[2]));

endmodule //CSAlike__0_113

module FA__2_1612 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__2_1612

module FA__2_1616 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__2_1616

module FA__2_1620 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__2_1620

module FA__2_1624 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n7;
wire CLOCK_slo__sro_n8;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n7), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n7), .B (CIN));
INV_X1 CLOCK_slo__sro_c3 (.ZN (CLOCK_slo__sro_n8), .A (A));
XNOR2_X1 CLOCK_slo__sro_c4 (.ZN (CLOCK_slo__sro_n7), .A (B), .B (CLOCK_slo__sro_n8));

endmodule //FA__2_1624

module FA__2_1628 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__mro_n10;
wire n_0_0;
wire CLOCK_slo__mro_n3;
wire CLOCK_slo__mro_n11;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__mro_n10), .B2 (CIN));
INV_X2 CLOCK_slo__mro_c7 (.ZN (CLOCK_slo__mro_n11), .A (B));
INV_X2 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n3), .A (CIN));
XNOR2_X1 CLOCK_slo__mro_c2 (.ZN (SUM), .A (CLOCK_slo__mro_n10), .B (CLOCK_slo__mro_n3));
XNOR2_X2 CLOCK_slo__mro_c8 (.ZN (CLOCK_slo__mro_n10), .A (CLOCK_slo__mro_n11), .B (A));

endmodule //FA__2_1628

module FA__2_1632 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1632

module FA__2_1636 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1636

module FA__2_1640 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1640

module FA__2_1644 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1644

module FA__2_1648 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1648

module FA__2_1652 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1652

module FA__2_1656 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1656

module FA__2_1660 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1660

module FA__2_1664 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n20;
wire CLOCK_slo__sro_n21;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n20), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n20), .B (CIN));
INV_X1 CLOCK_slo__sro_c5 (.ZN (CLOCK_slo__sro_n21), .A (A));
XNOR2_X2 CLOCK_slo__sro_c6 (.ZN (CLOCK_slo__sro_n20), .A (CLOCK_slo__sro_n21), .B (B));

endmodule //FA__2_1664

module FA__2_1668 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_sgo__sro_n7;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X1 CLOCK_sgo__sro_c3 (.ZN (CLOCK_sgo__sro_n7), .A1 (A), .A2 (B));
AOI21_X1 CLOCK_sgo__sro_c4 (.ZN (n_0_0), .A (CLOCK_sgo__sro_n7), .B1 (temp), .B2 (CIN));

endmodule //FA__2_1668

module FA__2_1672 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1672

module FA__2_1676 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire opt_ipo_n6;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (opt_ipo_n6), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (opt_ipo_n6), .B (B));
INV_X2 opt_ipo_c4 (.ZN (opt_ipo_n6), .A (A));

endmodule //FA__2_1676

module FA__2_1680 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1680

module FA__2_1684 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1684

module FA__2_1688 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1688

module FA__2_1692 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1692

module FA__2_1696 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1696

module FA__2_1700 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1700

module FA__2_1704 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1704

module FA__2_1708 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__n6;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__n6), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));
XOR2_X1 CLOCK_slo__c4 (.Z (CLOCK_slo__n6), .A (B), .B (A));

endmodule //FA__2_1708

module FA__2_1712 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__mro_n13;
wire CLOCK_slo__mro_n14;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__mro_n13), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (CLOCK_slo__mro_n13), .B (CIN));
INV_X1 CLOCK_slo__mro_c5 (.ZN (CLOCK_slo__mro_n14), .A (A));
XNOR2_X1 CLOCK_slo__mro_c6 (.ZN (CLOCK_slo__mro_n13), .A (B), .B (CLOCK_slo__mro_n14));

endmodule //FA__2_1712

module FA__2_1716 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1716

module FA__2_1720 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1720

module FA__2_1724 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__sro_n1;
wire slo__sro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__sro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__sro_n1), .B (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n2), .A (A));
XNOR2_X2 slo__sro_c2 (.ZN (slo__sro_n1), .A (B), .B (slo__sro_n2));

endmodule //FA__2_1724

module FA__2_1728 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__2_1728

module FA__2_1732 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__2_1732

module FA__2_1736 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__2_1736

module FA__2_1740 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__2_1740

module CSAlike__2_1765 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__2_1612 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .B (B[38]), .CIN (C[38]));
FA__2_1616 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .B (B[37]), .CIN (C[37]));
FA__2_1620 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .B (B[36]), .CIN (C[36]));
FA__2_1624 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__2_1628 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__2_1632 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__2_1636 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32])
    , .CIN (C[32]));
FA__2_1640 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__2_1644 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__2_1648 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__2_1652 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__2_1656 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__2_1660 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__2_1664 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25])
    , .CIN (C[25]));
FA__2_1668 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__2_1672 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__2_1676 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__2_1680 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__2_1684 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__2_1688 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__2_1692 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__2_1696 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]), .CIN (C[17]));
FA__2_1700 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16])
    , .CIN (C[16]));
FA__2_1704 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]), .CIN (C[15]));
FA__2_1708 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]), .CIN (C[14]));
FA__2_1712 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]), .CIN (C[13]));
FA__2_1716 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12])
    , .CIN (C[12]));
FA__2_1720 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]), .CIN (C[11]));
FA__2_1724 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10]), .CIN (C[10]));
FA__2_1728 genblk1_9_fa (.COUT (carry[10]), .SUM (result[9]), .A (A[9]), .B (B[9]), .CIN (C[9]));
FA__2_1732 genblk1_8_fa (.COUT (carry[9]), .SUM (result[8]), .A (A[8]), .B (B[8]), .CIN (C[8]));
FA__2_1736 genblk1_7_fa (.COUT (carry[8]), .SUM (result[7]), .A (A[7]), .B (B[7]));
FA__2_1740 genblk1_6_fa (.COUT (carry[7]), .SUM (result[6]), .A (A[6]), .B (B[6]));

endmodule //CSAlike__2_1765

module FA__2_1347 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1347

module FA__2_1351 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1351

module FA__2_1355 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1355

module FA__2_1359 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n27;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X2 CLOCK_slo__sro_c14 (.ZN (CLOCK_slo__sro_n27), .A (B));
XNOR2_X2 CLOCK_slo__sro_c15 (.ZN (temp), .A (CLOCK_slo__sro_n27), .B (A));

endmodule //FA__2_1359

module FA__2_1363 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1363

module FA__2_1367 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__2_1367

module FA__2_1371 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__mro_n23;
wire temp;
wire n_0_0;
wire slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
INV_X1 CLOCK_slo__mro_c9 (.ZN (CLOCK_slo__mro_n23), .A (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n7), .A (CIN));
XNOR2_X1 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n7));
XNOR2_X2 CLOCK_slo__mro_c10 (.ZN (temp), .A (CLOCK_slo__mro_n23), .B (A));

endmodule //FA__2_1371

module FA__2_1375 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1375

module FA__2_1379 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1379

module FA__2_1383 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__2_1383

module FA__2_1387 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1387

module FA__2_1391 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1391

module FA__2_1395 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1395

module FA__2_1399 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1399

module FA__2_1403 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1403

module FA__2_1407 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1407

module FA__2_1411 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1411

module FA__2_1415 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1415

module FA__2_1419 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n7), .A (CIN));
XNOR2_X1 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n7));

endmodule //FA__2_1419

module FA__2_1423 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1423

module FA__2_1427 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1427

module FA__2_1431 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1431

module FA__2_1435 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1435

module FA__2_1439 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1439

module FA__2_1443 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1443

module FA__2_1447 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1447

module FA__2_1451 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1451

module FA__2_1455 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1455

module FA__2_1459 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_11 (.ZN (n_0_8), .A (B));
INV_X1 i_0_10 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_9 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_5), .A1 (A), .A2 (B));
AOI21_X1 i_0_7 (.ZN (n_0_4), .A (CIN), .B1 (n_0_6), .B2 (n_0_5));
NAND3_X1 i_0_6 (.ZN (n_0_3), .A1 (n_0_6), .A2 (CIN), .A3 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_2), .A (n_0_3));
NOR2_X1 i_0_4 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_0 (.ZN (temp), .A (n_0_1));
INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));

endmodule //FA__2_1459

module FA__2_1463 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_11 (.ZN (n_0_8), .A (B));
INV_X1 i_0_10 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_9 (.ZN (n_0_6), .A1 (n_0_7), .A2 (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_5), .A1 (A), .A2 (B));
AOI21_X1 i_0_7 (.ZN (n_0_4), .A (CIN), .B1 (n_0_6), .B2 (n_0_5));
NAND3_X1 i_0_6 (.ZN (n_0_3), .A1 (n_0_6), .A2 (CIN), .A3 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_2), .A (n_0_3));
NOR2_X1 i_0_4 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_0 (.ZN (temp), .A (n_0_1));
INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));

endmodule //FA__2_1463

module FA__2_1467 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__2_1467

module CSAlike__2_1512 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__2_1347 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__2_1351 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__2_1355 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__2_1359 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38])
    , .CIN (C[38]));
FA__2_1363 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__2_1367 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__2_1371 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35])
    , .CIN (C[35]));
FA__2_1375 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34])
    , .CIN (C[34]));
FA__2_1379 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__2_1383 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__2_1387 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__2_1391 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__2_1395 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__2_1399 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__2_1403 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__2_1407 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26])
    , .CIN (C[26]));
FA__2_1411 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__2_1415 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__2_1419 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__2_1423 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__2_1427 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__2_1431 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__2_1435 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__2_1439 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__2_1443 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]), .CIN (C[17]));
FA__2_1447 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16]), .CIN (C[16]));
FA__2_1451 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]), .CIN (C[15]));
FA__2_1455 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]), .CIN (C[14]));
FA__2_1459 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]), .CIN (C[13]));
FA__2_1463 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12]), .CIN (C[12]));
FA__2_1467 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]));

endmodule //CSAlike__2_1512

module FA__2_1070 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__2_1070

module FA__2_1074 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__2_1074

module FA__2_1078 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__2_1078

module FA__2_1082 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1082

module FA__2_1086 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1086

module FA__2_1090 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1090

module FA__2_1094 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1094

module FA__2_1098 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1098

module FA__2_1102 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1102

module FA__2_1106 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1106

module FA__2_1110 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1110

module FA__2_1114 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1114

module FA__2_1118 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1118

module FA__2_1122 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1122

module FA__2_1126 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1126

module FA__2_1130 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__n4;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__n4), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
XOR2_X1 slo__c2 (.Z (slo__n4), .A (A), .B (B));

endmodule //FA__2_1130

module FA__2_1134 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1134

module FA__2_1138 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1138

module FA__2_1142 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1142

module FA__2_1146 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n3), .A (CIN));
XNOR2_X1 CLOCK_slo__mro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__mro_n3));

endmodule //FA__2_1146

module FA__2_1150 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1150

module FA__2_1154 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1154

module FA__2_1158 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n7), .A (CIN));
XNOR2_X1 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n7));

endmodule //FA__2_1158

module FA__2_1162 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1162

module FA__2_1166 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1166

module FA__2_1170 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1170

module FA__2_1174 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1174

module FA__2_1178 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1178

module FA__2_1182 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1182

module FA__2_1186 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_1186

module FA__2_1190 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n15;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X2 CLOCK_slo__sro_c9 (.ZN (CLOCK_slo__sro_n15), .A1 (A), .A2 (B));
AOI21_X1 CLOCK_slo__sro_c10 (.ZN (n_0_0), .A (CLOCK_slo__sro_n15), .B1 (temp), .B2 (CIN));

endmodule //FA__2_1190

module FA__2_1194 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__2_1194

module FA__2_1198 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__2_1198

module CSAlike__2_1259 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__2_1070 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .B (B[47]), .CIN (C[47]));
FA__2_1074 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .B (B[46]), .CIN (C[46]));
FA__2_1078 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .B (B[45]), .CIN (C[45]));
FA__2_1082 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__2_1086 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__2_1090 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__2_1094 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__2_1098 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__2_1102 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39])
    , .CIN (C[39]));
FA__2_1106 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__2_1110 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__2_1114 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__2_1118 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__2_1122 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__2_1126 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__2_1130 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__2_1134 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__2_1138 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__2_1142 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__2_1146 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__2_1150 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__2_1154 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__2_1158 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__2_1162 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__2_1166 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__2_1170 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__2_1174 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__2_1178 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__2_1182 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__2_1186 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__2_1190 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]), .CIN (C[17]));
FA__2_1194 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16]));
FA__2_1198 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]));

endmodule //CSAlike__2_1259

module FA__2_805 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_805

module FA__2_809 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_809

module FA__2_813 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_813

module FA__2_817 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_817

module FA__2_821 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_821

module FA__2_825 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_825

module FA__2_829 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_829

module FA__2_833 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_833

module FA__2_837 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__2_837

module FA__2_841 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n1), .A (B));
XNOR2_X1 slo__mro_c2 (.ZN (temp), .A (A), .B (slo__mro_n1));

endmodule //FA__2_841

module FA__2_845 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_845

module FA__2_849 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_849

module FA__2_853 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_853

module FA__2_857 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_857

module FA__2_861 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_861

module FA__2_865 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_865

module FA__2_869 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_869

module FA__2_873 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n14;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XNOR2_X1 CLOCK_slo__sro_c7 (.ZN (CLOCK_slo__sro_n14), .A (B), .B (A));
INV_X1 CLOCK_slo__sro_c8 (.ZN (temp), .A (CLOCK_slo__sro_n14));

endmodule //FA__2_873

module FA__2_877 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n3;
wire CLOCK_slo__sro_n4;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n3), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n3), .B (CIN));
INV_X1 CLOCK_slo__sro_c3 (.ZN (CLOCK_slo__sro_n4), .A (B));
XNOR2_X2 CLOCK_slo__sro_c4 (.ZN (CLOCK_slo__sro_n3), .A (CLOCK_slo__sro_n4), .B (A));

endmodule //FA__2_877

module FA__2_881 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__mro_n5;
wire CLOCK_slo__mro_n6;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__mro_n5), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (CLOCK_slo__mro_n5), .B (CIN));
INV_X2 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n6), .A (B));
XNOR2_X2 CLOCK_slo__mro_c2 (.ZN (CLOCK_slo__mro_n5), .A (A), .B (CLOCK_slo__mro_n6));

endmodule //FA__2_881

module FA__2_885 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;


AOI22_X2 i_0_2 (.ZN (COUT), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__2_885

module FA__2_889 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__sro_n1;
wire slo__sro_n2;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__sro_n1), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (slo__sro_n1), .B (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n2), .A (B));
XNOR2_X2 slo__sro_c2 (.ZN (slo__sro_n1), .A (slo__sro_n2), .B (A));

endmodule //FA__2_889

module FA__2_893 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__sro_n1;
wire slo__sro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__sro_n1), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (slo__sro_n1), .B (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n2), .A (A));
XNOR2_X1 slo__sro_c2 (.ZN (slo__sro_n1), .A (slo__sro_n2), .B (B));

endmodule //FA__2_893

module FA__2_897 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_897

module FA__2_901 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire sgo__sro_n7;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X1 sgo__sro_c3 (.ZN (sgo__sro_n7), .A1 (B), .A2 (A));
AOI21_X2 sgo__sro_c4 (.ZN (n_0_0), .A (sgo__sro_n7), .B1 (temp), .B2 (CIN));

endmodule //FA__2_901

module FA__2_905 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_spw_n34;
wire temp;
wire n_0_0;
wire CLOCK_slo__n22;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (CLOCK_spw_n34), .B1 (CLOCK_slo__n22), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (CLOCK_spw_n34));
XOR2_X1 CLOCK_slo__c8 (.Z (CLOCK_slo__n22), .A (A), .B (B));
CLKBUF_X1 CLOCK_spw__L1_c1_c13 (.Z (CLOCK_spw_n34), .A (B));

endmodule //FA__2_905

module FA__2_909 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_909

module FA__2_913 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_913

module FA__2_917 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_917

module FA__2_921 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_921

module FA__2_925 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__2_925

module CSAlike__2_1006 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__2_805 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .B (B[50]), .CIN (C[50]));
FA__2_809 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .B (B[49]), .CIN (C[49]));
FA__2_813 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__2_817 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__2_821 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__2_825 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__2_829 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__2_833 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__2_837 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__2_841 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__2_845 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__2_849 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__2_853 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__2_857 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__2_861 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__2_865 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__2_869 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__2_873 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33])
    , .CIN (C[33]));
FA__2_877 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__2_881 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__2_885 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__2_889 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__2_893 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__2_897 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__2_901 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__2_905 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__2_909 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__2_913 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__2_917 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__2_921 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__2_925 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]));

endmodule //CSAlike__2_1006

module FA__2_528 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__2_528

module FA__2_532 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__2_532

module FA__2_536 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__2_536

module FA__2_540 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_540

module FA__2_544 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_544

module FA__2_548 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_548

module FA__2_552 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_552

module FA__2_556 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n5;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n5), .A (CIN));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n5));

endmodule //FA__2_556

module FA__2_560 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_560

module FA__2_564 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__mro_n5;
wire CLOCK_slo__mro_n6;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__mro_n5), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__mro_n5), .B (CIN));
INV_X1 CLOCK_slo__mro_c5 (.ZN (CLOCK_slo__mro_n6), .A (B));
XNOR2_X2 CLOCK_slo__mro_c6 (.ZN (CLOCK_slo__mro_n5), .A (CLOCK_slo__mro_n6), .B (A));

endmodule //FA__2_564

module FA__2_568 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n3;
wire CLOCK_slo__sro_n4;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n3), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n3), .B (CIN));
INV_X1 CLOCK_slo__sro_c3 (.ZN (CLOCK_slo__sro_n4), .A (A));
XNOR2_X2 CLOCK_slo__sro_c4 (.ZN (CLOCK_slo__sro_n3), .A (CLOCK_slo__sro_n4), .B (B));

endmodule //FA__2_568

module FA__2_572 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_572

module FA__2_576 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_576

module FA__2_580 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_580

module FA__2_584 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n3), .A (CIN));
XNOR2_X1 slo__mro_c2 (.ZN (SUM), .A (temp), .B (slo__mro_n3));

endmodule //FA__2_584

module FA__2_588 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_588

module FA__2_592 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_592

module FA__2_596 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_596

module FA__2_600 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_600

module FA__2_604 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_604

module FA__2_608 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_608

module FA__2_612 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_612

module FA__2_616 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_616

module FA__2_620 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_620

module FA__2_624 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_624

module FA__2_628 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_628

module FA__2_632 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_632

module FA__2_636 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n3), .A (CIN));
XNOR2_X2 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n3));

endmodule //FA__2_636

module FA__2_640 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_640

module FA__2_644 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_644

module FA__2_648 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_648

module FA__2_652 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__2_652

module FA__2_656 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__2_656

module CSAlike__2_753 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__2_528 genblk1_56_fa (.COUT (carry[57]), .SUM (result[56]), .B (B[56]), .CIN (C[56]));
FA__2_532 genblk1_55_fa (.COUT (carry[56]), .SUM (result[55]), .B (B[55]), .CIN (C[55]));
FA__2_536 genblk1_54_fa (.COUT (carry[55]), .SUM (result[54]), .B (B[54]), .CIN (C[54]));
FA__2_540 genblk1_53_fa (.COUT (carry[54]), .SUM (result[53]), .A (A[53]), .B (B[53]), .CIN (C[53]));
FA__2_544 genblk1_52_fa (.COUT (carry[53]), .SUM (result[52]), .A (A[52]), .B (B[52]), .CIN (C[52]));
FA__2_548 genblk1_51_fa (.COUT (carry[52]), .SUM (result[51]), .A (A[51]), .B (B[51])
    , .CIN (C[51]));
FA__2_552 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .B (B[50]), .CIN (C[50]));
FA__2_556 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .B (B[49]), .CIN (C[49]));
FA__2_560 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__2_564 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__2_568 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__2_572 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__2_576 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__2_580 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__2_584 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__2_588 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__2_592 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__2_596 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__2_600 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__2_604 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__2_608 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__2_612 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__2_616 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__2_620 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__2_624 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__2_628 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__2_632 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__2_636 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__2_640 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__2_644 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27])
    , .CIN (C[27]));
FA__2_648 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__2_652 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]));
FA__2_656 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]));

endmodule //CSAlike__2_753

module FA__2_263 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_263

module FA__2_267 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_267

module FA__2_271 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_271

module FA__2_275 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_275

module FA__2_279 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_279

module FA__2_283 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_283

module FA__2_287 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_287

module FA__2_291 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_291

module FA__2_295 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_295

module FA__2_299 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_299

module FA__2_303 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_303

module FA__2_307 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_307

module FA__2_311 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X2 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n7), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n7));

endmodule //FA__2_311

module FA__2_315 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_315

module FA__2_319 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_319

module FA__2_323 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_323

module FA__2_327 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_327

module FA__2_331 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_331

module FA__2_335 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_335

module FA__2_339 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_339

module FA__2_343 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_343

module FA__2_347 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_347

module FA__2_351 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_351

module FA__2_355 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_355

module FA__2_359 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_359

module FA__2_363 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_363

module FA__2_367 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_367

module FA__2_371 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_371

module FA__2_375 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_375

module FA__2_379 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__2_379

module FA__2_383 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__2_383

module CSAlike__2_500 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__2_263 genblk1_59_fa (.COUT (carry[60]), .SUM (result[59]), .A (A[59]), .B (B[59]), .CIN (C[59]));
FA__2_267 genblk1_58_fa (.COUT (carry[59]), .SUM (result[58]), .A (A[58]), .B (B[58]), .CIN (C[58]));
FA__2_271 genblk1_57_fa (.COUT (carry[58]), .SUM (result[57]), .A (A[57]), .B (B[57]), .CIN (C[57]));
FA__2_275 genblk1_56_fa (.COUT (carry[57]), .SUM (result[56]), .A (A[56]), .B (B[56]), .CIN (C[56]));
FA__2_279 genblk1_55_fa (.COUT (carry[56]), .SUM (result[55]), .A (A[55]), .B (B[55]), .CIN (C[55]));
FA__2_283 genblk1_54_fa (.COUT (carry[55]), .SUM (result[54]), .A (A[54]), .B (B[54]), .CIN (C[54]));
FA__2_287 genblk1_53_fa (.COUT (carry[54]), .SUM (result[53]), .A (A[53]), .B (B[53]), .CIN (C[53]));
FA__2_291 genblk1_52_fa (.COUT (carry[53]), .SUM (result[52]), .A (A[52]), .B (B[52]), .CIN (C[52]));
FA__2_295 genblk1_51_fa (.COUT (carry[52]), .SUM (result[51]), .A (A[51]), .B (B[51]), .CIN (C[51]));
FA__2_299 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .B (B[50]), .CIN (C[50]));
FA__2_303 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .B (B[49]), .CIN (C[49]));
FA__2_307 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__2_311 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__2_315 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__2_319 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__2_323 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__2_327 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__2_331 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42])
    , .CIN (C[42]));
FA__2_335 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__2_339 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__2_343 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__2_347 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__2_351 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__2_355 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__2_359 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__2_363 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__2_367 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__2_371 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32])
    , .CIN (C[32]));
FA__2_375 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__2_379 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__2_383 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]));

endmodule //CSAlike__2_500

module FA__1_127 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__1_127

module FA__1_123 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X1 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (CIN), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__1_123

module FA__1_119 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;


INV_X1 i_0_14 (.ZN (n_0_12), .A (B));
INV_X1 i_0_13 (.ZN (n_0_11), .A (CIN));
NAND2_X1 i_0_12 (.ZN (n_0_10), .A1 (n_0_12), .A2 (n_0_11));
NAND2_X1 i_0_11 (.ZN (n_0_9), .A1 (B), .A2 (CIN));
NAND3_X1 i_0_10 (.ZN (n_0_8), .A1 (A), .A2 (n_0_10), .A3 (n_0_9));
INV_X1 i_0_9 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_10), .A2 (n_0_9));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (n_0_5), .A2 (n_0_8));
INV_X1 i_0_5 (.ZN (SUM), .A (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_3), .A1 (A), .A2 (B));
AOI21_X1 i_0_3 (.ZN (n_0_2), .A (n_0_11), .B1 (A), .B2 (B));
NAND2_X1 i_0_2 (.ZN (n_0_1), .A1 (n_0_7), .A2 (n_0_12));
NAND2_X1 i_0_1 (.ZN (n_0_0), .A1 (n_0_2), .A2 (n_0_1));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_0), .A2 (n_0_3));

endmodule //FA__1_119

module FA__1_115 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_115

module FA__1_111 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_111

module FA__1_107 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_107

module FA__1_103 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__1_103

module FA__1_99 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__sro_n1;
wire slo__sro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__sro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__sro_n1), .B (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n2), .A (B));
XNOR2_X2 slo__sro_c2 (.ZN (slo__sro_n1), .A (slo__sro_n2), .B (A));

endmodule //FA__1_99

module FA__1_95 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_95

module FA__1_91 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_8;
wire opt_ipo_n11;
wire opt_ipo_n12;


INV_X1 i_0_11 (.ZN (n_0_8), .A (B));
NAND2_X1 i_0_9 (.ZN (n_0_6), .A1 (opt_ipo_n12), .A2 (n_0_8));
NAND2_X1 i_0_8 (.ZN (n_0_5), .A1 (A), .A2 (B));
AOI21_X1 i_0_7 (.ZN (n_0_4), .A (CIN), .B1 (n_0_6), .B2 (n_0_5));
NAND3_X1 i_0_6 (.ZN (n_0_3), .A1 (n_0_6), .A2 (CIN), .A3 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_2), .A (n_0_3));
NOR2_X1 i_0_4 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_0 (.ZN (temp), .A (n_0_1));
INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (opt_ipo_n11), .A2 (B), .B1 (temp), .B2 (CIN));
INV_X1 opt_ipo_c7 (.ZN (opt_ipo_n11), .A (opt_ipo_n12));
INV_X1 opt_ipo_c8 (.ZN (opt_ipo_n12), .A (A));

endmodule //FA__1_91

module FA__1_87 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_87

module FA__1_83 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_83

module FA__1_79 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo__n45;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n38;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__n45), .B2 (CIN));
XOR2_X1 CLOCK_slo__c24 (.Z (CLOCK_slo__n45), .A (A), .B (B));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c18 (.ZN (CLOCK_slo__sro_n38), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c19 (.ZN (SUM), .A (CLOCK_slo__sro_n38), .B (temp));

endmodule //FA__1_79

module FA__1_75 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__1_75

module FA__1_71 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__n4;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__n4), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));
XOR2_X2 slo__c2 (.Z (slo__n4), .A (B), .B (A));

endmodule //FA__1_71

module FA__1_67 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__n1), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
XOR2_X2 slo__c1 (.Z (slo__n1), .A (A), .B (B));

endmodule //FA__1_67

module FA__1_63 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire CLOCK_sgo__sro_n45;
wire CLOCK_sgo__sro_n46;
wire CLOCK_slo__sro_n106;


INV_X1 i_0_12 (.ZN (n_0_9), .A (CIN));
INV_X1 i_0_11 (.ZN (n_0_8), .A (B));
INV_X1 i_0_10 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_9 (.ZN (n_0_6), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X2 i_0_7 (.ZN (n_0_4), .A1 (n_0_6), .A2 (CLOCK_slo__sro_n106));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_9));
NAND3_X1 i_0_5 (.ZN (n_0_2), .A1 (CIN), .A2 (n_0_6), .A3 (CLOCK_slo__sro_n106));
NAND2_X1 i_0_4 (.ZN (n_0_1), .A1 (n_0_3), .A2 (n_0_2));
INV_X2 i_0_1 (.ZN (SUM), .A (n_0_1));
INV_X1 i_0_0 (.ZN (temp), .A (n_0_4));
INV_X4 i_0_3 (.ZN (COUT), .A (n_0_0));
NAND2_X2 CLOCK_slo__sro_c75 (.ZN (CLOCK_slo__sro_n106), .A1 (B), .A2 (A));
NAND2_X1 CLOCK_sgo__sro_c21 (.ZN (CLOCK_sgo__sro_n46), .A1 (B), .A2 (A));
INV_X1 CLOCK_sgo__sro_c22 (.ZN (CLOCK_sgo__sro_n45), .A (CLOCK_sgo__sro_n46));
AOI21_X4 CLOCK_sgo__sro_c23 (.ZN (n_0_0), .A (CLOCK_sgo__sro_n45), .B1 (temp), .B2 (CIN));

endmodule //FA__1_63

module FA__1_59 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire slo__n7;
wire opt_ipo_n18;
wire CLOCK_slo__sro_n39;


INV_X2 i_0_3 (.ZN (COUT), .A (CLOCK_slo__sro_n39));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__n7), .B (CIN));
XNOR2_X2 slo__c9 (.ZN (slo__n7), .A (A), .B (B));
XNOR2_X2 slo__mro_c2 (.ZN (temp), .A (A), .B (B));
INV_X1 opt_ipo_c16 (.ZN (opt_ipo_n18), .A (A));
AOI22_X1 CLOCK_slo__sro_c34 (.ZN (CLOCK_slo__sro_n39), .A1 (CIN), .A2 (temp), .B1 (opt_ipo_n18), .B2 (B));

endmodule //FA__1_59

module FA__1_55 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


NAND2_X1 i_0_10 (.ZN (n_0_8), .A1 (n_0_1), .A2 (n_0_2));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (A), .A2 (B));
NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (CIN));
INV_X1 i_0_6 (.ZN (n_0_4), .A (CIN));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_8), .A2 (n_0_4), .A3 (n_0_7));
NAND2_X1 i_0_4 (.ZN (SUM), .A1 (n_0_5), .A2 (n_0_3));
INV_X1 i_0_3 (.ZN (n_0_2), .A (B));
INV_X1 i_0_2 (.ZN (n_0_1), .A (A));
AOI21_X2 i_0_1 (.ZN (n_0_0), .A (CIN), .B1 (A), .B2 (B));
AOI21_X4 i_0_0 (.ZN (COUT), .A (n_0_0), .B1 (n_0_2), .B2 (n_0_1));

endmodule //FA__1_55

module FA__1_51 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (B), .A2 (A));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__1_51

module FA__1_47 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X1 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (CIN), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (A), .A2 (B));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (A), .A2 (B));

endmodule //FA__1_47

module FA__1_43 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


INV_X1 i_0_11 (.ZN (n_0_9), .A (CIN));
INV_X1 i_0_10 (.ZN (n_0_8), .A (A));
NAND2_X1 i_0_9 (.ZN (n_0_7), .A1 (B), .A2 (n_0_8));
INV_X1 i_0_8 (.ZN (n_0_6), .A (B));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_6), .A2 (A));
AOI21_X1 i_0_6 (.ZN (n_0_4), .A (n_0_9), .B1 (n_0_5), .B2 (n_0_7));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (B), .A2 (A));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_6), .A2 (n_0_8));
AOI21_X1 i_0_3 (.ZN (n_0_1), .A (CIN), .B1 (n_0_2), .B2 (n_0_3));
NOR2_X1 i_0_2 (.ZN (SUM), .A1 (n_0_4), .A2 (n_0_1));
INV_X1 i_0_1 (.ZN (n_0_0), .A (n_0_4));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_0), .A2 (n_0_3));

endmodule //FA__1_43

module FA__1_39 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__1_39

module FA__1_35 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;


AOI22_X2 i_0_2 (.ZN (COUT), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__1_35

module FA__1_31 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_10 (.ZN (n_0_8), .A (B));
INV_X1 i_0_9 (.ZN (n_0_7), .A (A));
INV_X1 i_0_8 (.ZN (n_0_6), .A (CIN));
NAND2_X1 i_0_7 (.ZN (n_0_5), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_6 (.ZN (n_0_4), .A1 (A), .A2 (CIN));
NAND3_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_8), .A3 (n_0_4));
NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (B));
NAND2_X2 i_0_2 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_3));
INV_X1 i_0_1 (.ZN (n_0_0), .A (n_0_5));
OAI21_X1 i_0_0 (.ZN (COUT), .A (n_0_4), .B1 (n_0_0), .B2 (n_0_8));

endmodule //FA__1_31

module FA__1_27 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


NOR2_X1 i_0_10 (.ZN (n_0_8), .A1 (A), .A2 (B));
NAND2_X2 i_0_9 (.ZN (n_0_7), .A1 (A), .A2 (B));
INV_X1 i_0_8 (.ZN (n_0_6), .A (n_0_7));
OAI21_X2 i_0_7 (.ZN (n_0_5), .A (CIN), .B1 (n_0_6), .B2 (n_0_8));
INV_X1 i_0_6 (.ZN (n_0_4), .A (CIN));
INV_X1 i_0_5 (.ZN (n_0_3), .A (B));
INV_X1 i_0_4 (.ZN (n_0_2), .A (A));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (n_0_2), .A2 (n_0_3));
NAND3_X1 i_0_2 (.ZN (n_0_0), .A1 (n_0_1), .A2 (n_0_4), .A3 (n_0_7));
NAND2_X2 i_0_1 (.ZN (SUM), .A1 (n_0_5), .A2 (n_0_0));
OAI21_X1 i_0_0 (.ZN (COUT), .A (n_0_7), .B1 (n_0_8), .B2 (n_0_4));

endmodule //FA__1_27

module FA__1_23 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_23

module FA__1_19 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_19

module FA__1_15 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_15

module FA__1_11 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_11

module FA__1_7 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__1_7

module CSAlike__0_108 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__1_127 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .B (B[31]), .CIN (C[31]));
FA__1_123 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__1_119 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__1_115 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__1_111 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__1_107 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__1_103 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__1_99 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__1_95 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23])
    , .CIN (C[23]));
FA__1_91 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__1_87 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__1_83 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__1_79 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__1_75 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__1_71 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17])
    , .CIN (C[17]));
FA__1_67 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16])
    , .CIN (C[16]));
FA__1_63 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15])
    , .CIN (C[15]));
FA__1_59 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]), .CIN (C[14]));
FA__1_55 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]), .CIN (C[13]));
FA__1_51 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12]), .CIN (C[12]));
FA__1_47 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]), .CIN (C[11]));
FA__1_43 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10]), .CIN (C[10]));
FA__1_39 genblk1_9_fa (.COUT (carry[10]), .SUM (result[9]), .A (A[9]), .B (B[9]), .CIN (C[9]));
FA__1_35 genblk1_8_fa (.COUT (carry[9]), .SUM (result[8]), .A (A[8]), .B (B[8]), .CIN (C[8]));
FA__1_31 genblk1_7_fa (.COUT (carry[8]), .SUM (result[7]), .A (A[7]), .B (B[7]), .CIN (C[7]));
FA__1_27 genblk1_6_fa (.COUT (carry[7]), .SUM (result[6]), .A (A[6]), .B (B[6]), .CIN (C[6]));
FA__1_23 genblk1_5_fa (.COUT (carry[6]), .SUM (result[5]), .A (A[5]), .B (B[5]), .CIN (C[5]));
FA__1_19 genblk1_4_fa (.COUT (carry[5]), .SUM (result[4]), .A (A[4]), .B (B[4]), .CIN (C[4]));
FA__1_15 genblk1_3_fa (.COUT (carry[4]), .SUM (result[3]), .A (A[3]), .B (B[3]), .CIN (C[3]));
FA__1_11 genblk1_2_fa (.COUT (carry[3]), .SUM (result[2]), .A (A[2]), .B (B[2]), .CIN (C[2]));
FA__1_7 genblk1_1_fa (.COUT (carry[2]), .SUM (result[1]), .A (A[1]), .B (B[1]));

endmodule //CSAlike__0_108

module FA__1_2387 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__1_2387

module FA__1_2391 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__mro_n1;
wire slo__mro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__mro_n1), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (slo__mro_n1), .B (CIN));
INV_X1 slo__mro_c1 (.ZN (slo__mro_n2), .A (B));
XNOR2_X1 slo__mro_c2 (.ZN (slo__mro_n1), .A (A), .B (slo__mro_n2));

endmodule //FA__1_2391

module FA__1_2395 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2395

module FA__1_2399 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2399

module FA__1_2403 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2403

module FA__1_2407 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__1_2407

module FA__1_2411 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2411

module FA__1_2415 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2415

module FA__1_2419 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2419

module FA__1_2423 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2423

module FA__1_2427 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2427

module FA__1_2431 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2431

module FA__1_2435 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2435

module FA__1_2439 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;


AOI22_X1 i_0_2 (.ZN (COUT), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2439

module FA__1_2443 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2443

module FA__1_2447 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2447

module FA__1_2451 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2451

module FA__1_2455 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X2 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n1), .A (B));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (temp), .A (A), .B (CLOCK_slo__sro_n1));

endmodule //FA__1_2455

module FA__1_2459 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X2 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n1), .A (B));
XNOR2_X2 CLOCK_slo__sro_c2 (.ZN (temp), .A (CLOCK_slo__sro_n1), .B (A));

endmodule //FA__1_2459

module FA__1_2463 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n12;
wire CLOCK_slo__sro_n13;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n12), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n12), .B (CIN));
INV_X2 CLOCK_slo__sro_c4 (.ZN (CLOCK_slo__sro_n13), .A (A));
XNOR2_X2 CLOCK_slo__sro_c5 (.ZN (CLOCK_slo__sro_n12), .A (CLOCK_slo__sro_n13), .B (B));

endmodule //FA__1_2463

module FA__1_2467 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2467

module FA__1_2471 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__1_2471

module FA__1_2475 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n20;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 CLOCK_slo__mro_c5 (.ZN (CLOCK_slo__mro_n20), .A (A));
XNOR2_X1 CLOCK_slo__mro_c6 (.ZN (temp), .A (CLOCK_slo__mro_n20), .B (B));

endmodule //FA__1_2475

module FA__1_2479 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2479

module FA__1_2483 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (B), .A2 (A));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_5), .A2 (n_0_4));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__1_2483

module FA__1_2487 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;


NAND2_X1 i_0_8 (.ZN (n_0_6), .A1 (A), .A2 (B));
INV_X1 i_0_7 (.ZN (n_0_5), .A (B));
INV_X1 i_0_6 (.ZN (n_0_4), .A (A));
NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (n_0_4), .A2 (n_0_5));
NAND3_X1 i_0_4 (.ZN (n_0_2), .A1 (n_0_3), .A2 (CIN), .A3 (n_0_6));
INV_X1 i_0_3 (.ZN (n_0_1), .A (n_0_2));
AOI21_X1 i_0_2 (.ZN (n_0_0), .A (CIN), .B1 (n_0_3), .B2 (n_0_6));
NOR2_X1 i_0_1 (.ZN (SUM), .A1 (n_0_1), .A2 (n_0_0));
NAND2_X1 i_0_0 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_6));

endmodule //FA__1_2487

module FA__1_2491 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2491

module FA__1_2495 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2495

module FA__1_2499 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2499

module FA__1_2503 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2503

module FA__1_2507 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__1_2507

module CSAlike__1_2524 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__1_2387 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .B (B[34]), .CIN (C[34]));
FA__1_2391 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__1_2395 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__1_2399 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__1_2403 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__1_2407 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__1_2411 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__1_2415 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__1_2419 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__1_2423 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__1_2427 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__1_2431 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__1_2435 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__1_2439 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__1_2443 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__1_2447 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__1_2451 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__1_2455 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]), .CIN (C[17]));
FA__1_2459 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16]), .CIN (C[16]));
FA__1_2463 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]), .CIN (C[15]));
FA__1_2467 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]), .CIN (C[14]));
FA__1_2471 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]), .CIN (C[13]));
FA__1_2475 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12])
    , .CIN (C[12]));
FA__1_2479 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]), .CIN (C[11]));
FA__1_2483 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10]), .CIN (C[10]));
FA__1_2487 genblk1_9_fa (.COUT (carry[10]), .SUM (result[9]), .A (A[9]), .B (B[9]), .CIN (C[9]));
FA__1_2491 genblk1_8_fa (.COUT (carry[9]), .SUM (result[8]), .A (A[8]), .B (B[8]), .CIN (C[8]));
FA__1_2495 genblk1_7_fa (.COUT (carry[8]), .SUM (result[7]), .A (A[7]), .B (B[7]), .CIN (C[7]));
FA__1_2499 genblk1_6_fa (.COUT (carry[7]), .SUM (result[6]), .A (A[6]), .B (B[6]), .CIN (C[6]));
FA__1_2503 genblk1_5_fa (.COUT (carry[6]), .SUM (result[5]), .A (A[5]), .B (B[5]), .CIN (C[5]));
FA__1_2507 genblk1_4_fa (.COUT (carry[5]), .SUM (result[4]), .A (A[4]), .B (B[4]));

endmodule //CSAlike__1_2524

module FA__1_2122 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__1_2122

module FA__1_2126 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2126

module FA__1_2130 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n1;
wire CLOCK_slo__sro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n1), .B (CIN));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n2), .A (B));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (CLOCK_slo__sro_n1), .A (A), .B (CLOCK_slo__sro_n2));

endmodule //FA__1_2130

module FA__1_2134 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2134

module FA__1_2138 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2138

module FA__1_2142 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n7), .A (CIN));
XNOR2_X1 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n7));

endmodule //FA__1_2142

module FA__1_2146 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2146

module FA__1_2150 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2150

module FA__1_2154 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2154

module FA__1_2158 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2158

module FA__1_2162 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2162

module FA__1_2166 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2166

module FA__1_2170 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n7), .A (CIN));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n7));

endmodule //FA__1_2170

module FA__1_2174 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2174

module FA__1_2178 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2178

module FA__1_2182 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2182

module FA__1_2186 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2186

module FA__1_2190 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2190

module FA__1_2194 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2194

module FA__1_2198 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2198

module FA__1_2202 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2202

module FA__1_2206 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2206

module FA__1_2210 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2210

module FA__1_2214 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2214

module FA__1_2218 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2218

module FA__1_2222 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n9;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c3 (.ZN (CLOCK_slo__sro_n9), .A (CIN));
XNOR2_X1 CLOCK_slo__sro_c4 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n9));

endmodule //FA__1_2222

module FA__1_2226 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2226

module FA__1_2230 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__1_2230

module FA__1_2234 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));
INV_X4 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n3), .A (CIN));
XNOR2_X2 CLOCK_slo__mro_c2 (.ZN (SUM), .A (CLOCK_slo__mro_n3), .B (temp));

endmodule //FA__1_2234

module FA__1_2238 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_2238

module FA__1_2242 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__1_2242

module CSAlike__1_2271 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__1_2122 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .B (B[37]), .CIN (C[37]));
FA__1_2126 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__1_2130 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__1_2134 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__1_2138 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__1_2142 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__1_2146 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__1_2150 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__1_2154 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__1_2158 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__1_2162 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__1_2166 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__1_2170 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__1_2174 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__1_2178 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__1_2182 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__1_2186 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__1_2190 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__1_2194 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__1_2198 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__1_2202 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]), .CIN (C[17]));
FA__1_2206 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16]), .CIN (C[16]));
FA__1_2210 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]), .CIN (C[15]));
FA__1_2214 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]), .CIN (C[14]));
FA__1_2218 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]), .CIN (C[13]));
FA__1_2222 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12]), .CIN (C[12]));
FA__1_2226 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]), .CIN (C[11]));
FA__1_2230 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10]), .CIN (C[10]));
FA__1_2234 genblk1_9_fa (.COUT (carry[10]), .SUM (result[9]), .A (A[9]), .B (B[9]), .CIN (C[9]));
FA__1_2238 genblk1_8_fa (.COUT (carry[9]), .SUM (result[8]), .A (A[8]), .B (B[8]), .CIN (C[8]));
FA__1_2242 genblk1_7_fa (.COUT (carry[8]), .SUM (result[7]), .A (A[7]), .B (B[7]));

endmodule //CSAlike__1_2271

module FA__1_1857 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__1_1857

module FA__1_1861 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1861

module FA__1_1865 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_opt_ipo_n4;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (CLOCK_opt_ipo_n4), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
CLKBUF_X1 CLOCK_opt_ipo_c2 (.Z (CLOCK_opt_ipo_n4), .A (B));

endmodule //FA__1_1865

module FA__1_1869 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1869

module FA__1_1873 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire sgo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X1 sgo__sro_c3 (.ZN (sgo__sro_n7), .A1 (A), .A2 (B));
AOI21_X1 sgo__sro_c4 (.ZN (n_0_0), .A (sgo__sro_n7), .B1 (temp), .B2 (CIN));

endmodule //FA__1_1873

module FA__1_1877 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n5;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n5), .A (CIN));
XNOR2_X2 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n5));

endmodule //FA__1_1877

module FA__1_1881 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n13;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XNOR2_X2 CLOCK_slo__mro_c12 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n13));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c6 (.ZN (CLOCK_slo__sro_n13), .A (CIN));

endmodule //FA__1_1881

module FA__1_1885 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1885

module FA__1_1889 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1889

module FA__1_1893 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__1_1893

module FA__1_1897 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1897

module FA__1_1901 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1901

module FA__1_1905 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo_n8;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n9;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (CLOCK_slo_n8), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
CLKBUF_X1 CLOCK_slo___L1_c1_c1 (.Z (CLOCK_slo_n8), .A (B));
INV_X1 CLOCK_slo__sro_c4 (.ZN (CLOCK_slo__sro_n9), .A (B));
XNOR2_X2 CLOCK_slo__sro_c5 (.ZN (temp), .A (CLOCK_slo__sro_n9), .B (A));

endmodule //FA__1_1905

module FA__1_1909 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1909

module FA__1_1913 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n7), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n7));

endmodule //FA__1_1913

module FA__1_1917 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1917

module FA__1_1921 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1921

module FA__1_1925 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1925

module FA__1_1929 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n1), .A (B));
XNOR2_X1 slo__sro_c2 (.ZN (temp), .A (slo__sro_n1), .B (A));

endmodule //FA__1_1929

module FA__1_1933 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1933

module FA__1_1937 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1937

module FA__1_1941 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1941

module FA__1_1945 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1945

module FA__1_1949 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1949

module FA__1_1953 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1953

module FA__1_1957 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1957

module FA__1_1961 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1961

module FA__1_1965 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire temp;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;


INV_X1 i_0_11 (.ZN (n_0_8), .A (B));
INV_X1 i_0_10 (.ZN (n_0_7), .A (A));
NAND2_X1 i_0_9 (.ZN (n_0_6), .A1 (n_0_8), .A2 (n_0_7));
NAND2_X1 i_0_8 (.ZN (n_0_5), .A1 (B), .A2 (A));
AOI21_X1 i_0_7 (.ZN (n_0_4), .A (CIN), .B1 (n_0_6), .B2 (n_0_5));
NAND3_X1 i_0_6 (.ZN (n_0_3), .A1 (n_0_6), .A2 (CIN), .A3 (n_0_5));
INV_X1 i_0_5 (.ZN (n_0_2), .A (n_0_3));
NOR2_X1 i_0_4 (.ZN (SUM), .A1 (n_0_2), .A2 (n_0_4));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (n_0_6), .A2 (n_0_5));
INV_X1 i_0_0 (.ZN (temp), .A (n_0_1));
INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));

endmodule //FA__1_1965

module FA__1_1969 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;


NOR2_X1 i_0_6 (.ZN (SUM), .A1 (n_0_3), .A2 (n_0_4));
AOI21_X1 i_0_5 (.ZN (n_0_4), .A (CIN), .B1 (n_0_0), .B2 (n_0_1));
INV_X1 i_0_4 (.ZN (n_0_3), .A (n_0_2));
NAND2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_2), .A2 (n_0_1));
NAND3_X1 i_0_2 (.ZN (n_0_2), .A1 (n_0_0), .A2 (CIN), .A3 (n_0_1));
NAND2_X1 i_0_1 (.ZN (n_0_1), .A1 (B), .A2 (A));
OR2_X1 i_0_0 (.ZN (n_0_0), .A1 (B), .A2 (A));

endmodule //FA__1_1969

module FA__1_1973 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NOR2_X1 i_0_5 (.ZN (n_0_2), .A1 (B), .A2 (A));
AOI21_X1 i_0_4 (.ZN (n_0_1), .A (CIN), .B1 (B), .B2 (A));
NOR2_X1 i_0_3 (.ZN (COUT), .A1 (n_0_1), .A2 (n_0_2));
XNOR2_X1 i_0_2 (.ZN (n_0_0), .A (B), .B (A));
INV_X1 i_0_0 (.ZN (temp), .A (n_0_0));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));

endmodule //FA__1_1973

module FA__1_1977 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__1_1977

module CSAlike__1_2018 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__1_1857 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .B (B[40]), .CIN (C[40]));
FA__1_1861 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__1_1865 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__1_1869 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__1_1873 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__1_1877 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__1_1881 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__1_1885 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33])
    , .CIN (C[33]));
FA__1_1889 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__1_1893 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__1_1897 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__1_1901 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__1_1905 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__1_1909 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__1_1913 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__1_1917 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__1_1921 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__1_1925 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__1_1929 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__1_1933 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__1_1937 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__1_1941 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__1_1945 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__1_1949 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]), .CIN (C[17]));
FA__1_1953 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16]), .CIN (C[16]));
FA__1_1957 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]), .CIN (C[15]));
FA__1_1961 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]), .CIN (C[14]));
FA__1_1965 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]), .CIN (C[13]));
FA__1_1969 genblk1_12_fa (.COUT (carry[13]), .SUM (result[12]), .A (A[12]), .B (B[12]), .CIN (C[12]));
FA__1_1973 genblk1_11_fa (.COUT (carry[12]), .SUM (result[11]), .A (A[11]), .B (B[11]), .CIN (C[11]));
FA__1_1977 genblk1_10_fa (.COUT (carry[11]), .SUM (result[10]), .A (A[10]), .B (B[10]));

endmodule //CSAlike__1_2018

module FA__1_1592 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__1_1592

module FA__1_1596 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__n29;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__n29), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
XOR2_X1 CLOCK_slo__c12 (.Z (CLOCK_slo__n29), .A (A), .B (B));

endmodule //FA__1_1596

module FA__1_1600 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__1_1600

module FA__1_1604 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire CLOCK_slo__sro_n18;
wire CLOCK_slo__sro_n19;


INV_X1 i_0_3 (.ZN (COUT), .A (CLOCK_slo__sro_n18));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
AND2_X1 CLOCK_slo__sro_c9 (.ZN (CLOCK_slo__sro_n19), .A1 (B), .A2 (A));
AOI21_X1 CLOCK_slo__sro_c10 (.ZN (CLOCK_slo__sro_n18), .A (CLOCK_slo__sro_n19), .B1 (temp), .B2 (CIN));

endmodule //FA__1_1604

module FA__1_1608 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__1_1608

module FA__1_1612 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__n1), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));
XOR2_X1 CLOCK_slo__c1 (.Z (CLOCK_slo__n1), .A (B), .B (A));

endmodule //FA__1_1612

module FA__1_1616 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1616

module FA__1_1620 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__1_1620

module FA__1_1624 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1624

module FA__1_1628 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1628

module FA__1_1632 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1632

module FA__1_1636 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1636

module FA__1_1640 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1640

module FA__1_1644 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1644

module FA__1_1648 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1648

module FA__1_1652 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1652

module FA__1_1656 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1656

module FA__1_1660 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1660

module FA__1_1664 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1664

module FA__1_1668 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1668

module FA__1_1672 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1672

module FA__1_1676 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1676

module FA__1_1680 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1680

module FA__1_1684 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1684

module FA__1_1688 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1688

module FA__1_1692 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1692

module FA__1_1696 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1696

module FA__1_1700 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1700

module FA__1_1704 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1704

module FA__1_1708 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1708

module FA__1_1712 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__1_1712

module CSAlike__1_1765 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__1_1592 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .B (B[43]), .CIN (C[43]));
FA__1_1596 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42])
    , .CIN (C[42]));
FA__1_1600 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__1_1604 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__1_1608 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__1_1612 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__1_1616 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__1_1620 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36])
    , .CIN (C[36]));
FA__1_1624 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__1_1628 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__1_1632 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__1_1636 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__1_1640 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31])
    , .CIN (C[31]));
FA__1_1644 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30])
    , .CIN (C[30]));
FA__1_1648 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__1_1652 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__1_1656 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__1_1660 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__1_1664 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__1_1668 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__1_1672 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__1_1676 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__1_1680 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__1_1684 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__1_1688 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__1_1692 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__1_1696 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17]), .CIN (C[17]));
FA__1_1700 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16])
    , .CIN (C[16]));
FA__1_1704 genblk1_15_fa (.COUT (carry[16]), .SUM (result[15]), .A (A[15]), .B (B[15]), .CIN (C[15]));
FA__1_1708 genblk1_14_fa (.COUT (carry[15]), .SUM (result[14]), .A (A[14]), .B (B[14]), .CIN (C[14]));
FA__1_1712 genblk1_13_fa (.COUT (carry[14]), .SUM (result[13]), .A (A[13]), .B (B[13]));

endmodule //CSAlike__1_1765

module FA__1_1327 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__1_1327

module FA__1_1331 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1331

module FA__1_1335 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1335

module FA__1_1339 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire CLOCK_slo__sro_n1;
wire CLOCK_slo__sro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (CLOCK_slo__sro_n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (CLOCK_slo__sro_n1), .B (CIN));
INV_X2 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n2), .A (B));
XNOR2_X2 CLOCK_slo__sro_c2 (.ZN (CLOCK_slo__sro_n1), .A (CLOCK_slo__sro_n2), .B (A));

endmodule //FA__1_1339

module FA__1_1343 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire spw__n17;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (spw__n17), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
CLKBUF_X1 spw__L1_c17 (.Z (spw__n17), .A (temp));

endmodule //FA__1_1343

module FA__1_1347 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1347

module FA__1_1351 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__1_1351

module FA__1_1355 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n5;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n5), .A (CIN));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n5));

endmodule //FA__1_1355

module FA__1_1359 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1359

module FA__1_1363 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1363

module FA__1_1367 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire spw_n8;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (spw_n8), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
CLKBUF_X1 spw__L1_c1_c1 (.Z (spw_n8), .A (B));

endmodule //FA__1_1367

module FA__1_1371 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1371

module FA__1_1375 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1375

module FA__1_1379 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1379

module FA__1_1383 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1383

module FA__1_1387 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1387

module FA__1_1391 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1391

module FA__1_1395 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1395

module FA__1_1399 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n3), .A (CIN));
XNOR2_X1 CLOCK_slo__mro_c2 (.ZN (SUM), .A (temp), .B (CLOCK_slo__mro_n3));

endmodule //FA__1_1399

module FA__1_1403 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1403

module FA__1_1407 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1407

module FA__1_1411 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire CLOCK_slo_n10;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (CLOCK_slo_n10), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
CLKBUF_X1 CLOCK_slo___L1_c1_c3 (.Z (CLOCK_slo_n10), .A (A));

endmodule //FA__1_1411

module FA__1_1415 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1415

module FA__1_1419 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1419

module FA__1_1423 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1423

module FA__1_1427 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1427

module FA__1_1431 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1431

module FA__1_1435 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1435

module FA__1_1439 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1439

module FA__1_1443 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1443

module FA__1_1447 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__1_1447

module CSAlike__1_1512 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__1_1327 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .B (B[46]), .CIN (C[46]));
FA__1_1331 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__1_1335 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__1_1339 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43])
    , .CIN (C[43]));
FA__1_1343 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__1_1347 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__1_1351 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__1_1355 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__1_1359 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__1_1363 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__1_1367 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__1_1371 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__1_1375 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__1_1379 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__1_1383 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__1_1387 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__1_1391 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__1_1395 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__1_1399 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__1_1403 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__1_1407 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__1_1411 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__1_1415 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__1_1419 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__1_1423 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__1_1427 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__1_1431 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__1_1435 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]), .CIN (C[19]));
FA__1_1439 genblk1_18_fa (.COUT (carry[19]), .SUM (result[18]), .A (A[18]), .B (B[18]), .CIN (C[18]));
FA__1_1443 genblk1_17_fa (.COUT (carry[18]), .SUM (result[17]), .A (A[17]), .B (B[17])
    , .CIN (C[17]));
FA__1_1447 genblk1_16_fa (.COUT (carry[17]), .SUM (result[16]), .A (A[16]), .B (B[16]));

endmodule //CSAlike__1_1512

module FA__1_1062 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__1_1062

module FA__1_1066 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n3;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n3), .A (CIN));
XNOR2_X1 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n3));

endmodule //FA__1_1066

module FA__1_1070 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1070

module FA__1_1074 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1074

module FA__1_1078 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1078

module FA__1_1082 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1082

module FA__1_1086 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1086

module FA__1_1090 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1090

module FA__1_1094 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1094

module FA__1_1098 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));

endmodule //FA__1_1098

module FA__1_1102 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__mro_n9;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__mro_c3 (.ZN (slo__mro_n9), .A (CIN));
XNOR2_X1 slo__mro_c4 (.ZN (SUM), .A (temp), .B (slo__mro_n9));

endmodule //FA__1_1102

module FA__1_1106 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1106

module FA__1_1110 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__mro_n4;
wire slo__mro_n5;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__mro_n4), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (slo__mro_n4), .B (CIN));
INV_X1 slo__mro_c2 (.ZN (slo__mro_n5), .A (B));
XNOR2_X2 slo__mro_c3 (.ZN (slo__mro_n4), .A (slo__mro_n5), .B (A));

endmodule //FA__1_1110

module FA__1_1114 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1114

module FA__1_1118 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1118

module FA__1_1122 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1122

module FA__1_1126 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n12;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (B), .B (A));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n12), .A (CIN));
XNOR2_X1 slo__sro_c4 (.ZN (SUM), .A (temp), .B (slo__sro_n12));

endmodule //FA__1_1126

module FA__1_1130 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1130

module FA__1_1134 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n19;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c4 (.ZN (CLOCK_slo__sro_n19), .A (CIN));
XNOR2_X1 CLOCK_slo__sro_c5 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n19));

endmodule //FA__1_1134

module FA__1_1138 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__n1;
wire CLOCK_slo__sro_n6;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__n1), .B2 (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
XOR2_X1 slo__c1 (.Z (slo__n1), .A (A), .B (B));
INV_X2 CLOCK_slo__sro_c4 (.ZN (CLOCK_slo__sro_n6), .A (CIN));
XNOR2_X2 CLOCK_slo__sro_c5 (.ZN (SUM), .A (temp), .B (CLOCK_slo__sro_n6));

endmodule //FA__1_1138

module FA__1_1142 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1142

module FA__1_1146 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n12;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c3 (.ZN (slo__sro_n12), .A (CIN));
XNOR2_X1 slo__sro_c4 (.ZN (SUM), .A (temp), .B (slo__sro_n12));

endmodule //FA__1_1146

module FA__1_1150 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1150

module FA__1_1154 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1154

module FA__1_1158 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1158

module FA__1_1162 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1162

module FA__1_1166 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1166

module FA__1_1170 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1170

module FA__1_1174 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1174

module FA__1_1178 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_1178

module FA__1_1182 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__1_1182

module CSAlike__1_1259 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__1_1062 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .B (B[49]), .CIN (C[49]));
FA__1_1066 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__1_1070 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__1_1074 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__1_1078 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__1_1082 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__1_1086 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__1_1090 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__1_1094 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__1_1098 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__1_1102 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__1_1106 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__1_1110 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__1_1114 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__1_1118 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35])
    , .CIN (C[35]));
FA__1_1122 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__1_1126 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33])
    , .CIN (C[33]));
FA__1_1130 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32])
    , .CIN (C[32]));
FA__1_1134 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31])
    , .CIN (C[31]));
FA__1_1138 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__1_1142 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29])
    , .CIN (C[29]));
FA__1_1146 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28])
    , .CIN (C[28]));
FA__1_1150 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27])
    , .CIN (C[27]));
FA__1_1154 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26])
    , .CIN (C[26]));
FA__1_1158 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25])
    , .CIN (C[25]));
FA__1_1162 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24])
    , .CIN (C[24]));
FA__1_1166 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__1_1170 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]), .CIN (C[22]));
FA__1_1174 genblk1_21_fa (.COUT (carry[22]), .SUM (result[21]), .A (A[21]), .B (B[21]), .CIN (C[21]));
FA__1_1178 genblk1_20_fa (.COUT (carry[21]), .SUM (result[20]), .A (A[20]), .B (B[20]), .CIN (C[20]));
FA__1_1182 genblk1_19_fa (.COUT (carry[20]), .SUM (result[19]), .A (A[19]), .B (B[19]));

endmodule //CSAlike__1_1259

module FA__1_797 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__1_797

module FA__1_801 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_801

module FA__1_805 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_805

module FA__1_809 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_809

module FA__1_813 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n1), .A (A));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (temp), .A (B), .B (CLOCK_slo__sro_n1));

endmodule //FA__1_813

module FA__1_817 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_817

module FA__1_821 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X2 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_821

module FA__1_825 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_825

module FA__1_829 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_829

module FA__1_833 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_833

module FA__1_837 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_837

module FA__1_841 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire sgo__sro_n7;
wire sgo__sro_n8;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
NAND2_X1 sgo__sro_c3 (.ZN (sgo__sro_n8), .A1 (A), .A2 (B));
INV_X1 sgo__sro_c4 (.ZN (sgo__sro_n7), .A (sgo__sro_n8));
AOI21_X1 sgo__sro_c5 (.ZN (n_0_0), .A (sgo__sro_n7), .B1 (temp), .B2 (CIN));

endmodule //FA__1_841

module FA__1_845 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_845

module FA__1_849 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_849

module FA__1_853 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_853

module FA__1_857 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_857

module FA__1_861 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_861

module FA__1_865 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_865

module FA__1_869 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_869

module FA__1_873 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire n_0_0;
wire slo__sro_n1;
wire slo__sro_n2;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo__sro_n1), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (slo__sro_n1), .B (CIN));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n2), .A (B));
XNOR2_X1 slo__sro_c2 (.ZN (slo__sro_n1), .A (A), .B (slo__sro_n2));

endmodule //FA__1_873

module FA__1_877 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_877

module FA__1_881 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_881

module FA__1_885 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n17;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X1 CLOCK_slo__sro_c4 (.ZN (CLOCK_slo__sro_n17), .A (B));
XNOR2_X2 CLOCK_slo__sro_c5 (.ZN (temp), .A (A), .B (CLOCK_slo__sro_n17));

endmodule //FA__1_885

module FA__1_889 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_889

module FA__1_893 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_893

module FA__1_897 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_897

module FA__1_901 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X2 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_901

module FA__1_905 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_905

module FA__1_909 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_909

module FA__1_913 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_913

module FA__1_917 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__1_917

module CSAlike__1_1006 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__1_797 genblk1_52_fa (.COUT (carry[53]), .SUM (result[52]), .B (B[52]), .CIN (C[52]));
FA__1_801 genblk1_51_fa (.COUT (carry[52]), .SUM (result[51]), .A (A[51]), .B (B[51]), .CIN (C[51]));
FA__1_805 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .B (B[50]), .CIN (C[50]));
FA__1_809 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .B (B[49]), .CIN (C[49]));
FA__1_813 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__1_817 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__1_821 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__1_825 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__1_829 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__1_833 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__1_837 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__1_841 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__1_845 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__1_849 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__1_853 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__1_857 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__1_861 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__1_865 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__1_869 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__1_873 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__1_877 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__1_881 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__1_885 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30])
    , .CIN (C[30]));
FA__1_889 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__1_893 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__1_897 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__1_901 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__1_905 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]), .CIN (C[25]));
FA__1_909 genblk1_24_fa (.COUT (carry[25]), .SUM (result[24]), .A (A[24]), .B (B[24]), .CIN (C[24]));
FA__1_913 genblk1_23_fa (.COUT (carry[24]), .SUM (result[23]), .A (A[23]), .B (B[23]), .CIN (C[23]));
FA__1_917 genblk1_22_fa (.COUT (carry[23]), .SUM (result[22]), .A (A[22]), .B (B[22]));

endmodule //CSAlike__1_1006

module FA__1_532 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__1_532

module FA__1_536 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_536

module FA__1_540 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_540

module FA__1_544 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_544

module FA__1_548 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_548

module FA__1_552 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_552

module FA__1_556 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_556

module FA__1_560 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_560

module FA__1_564 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo___n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (slo___n1), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));
CLKBUF_X1 slo___L1_c1 (.Z (slo___n1), .A (temp));

endmodule //FA__1_564

module FA__1_568 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_568

module FA__1_572 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_572

module FA__1_576 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_576

module FA__1_580 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_580

module FA__1_584 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_584

module FA__1_588 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_588

module FA__1_592 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_592

module FA__1_596 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_596

module FA__1_600 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_600

module FA__1_604 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_604

module FA__1_608 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_608

module FA__1_612 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_612

module FA__1_616 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_616

module FA__1_620 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_620

module FA__1_624 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_624

module FA__1_628 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_628

module FA__1_632 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__mro_n1;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
INV_X2 CLOCK_slo__mro_c1 (.ZN (CLOCK_slo__mro_n1), .A (B));
XNOR2_X2 CLOCK_slo__mro_c2 (.ZN (temp), .A (A), .B (CLOCK_slo__mro_n1));

endmodule //FA__1_632

module FA__1_636 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_636

module FA__1_640 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_640

module FA__1_644 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n7), .A (CIN));
XNOR2_X1 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n7));

endmodule //FA__1_644

module FA__1_648 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_648

module FA__1_652 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__1_652

module CSAlike__1_753 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__1_532 genblk1_55_fa (.COUT (carry[56]), .SUM (result[55]), .B (B[55]), .CIN (C[55]));
FA__1_536 genblk1_54_fa (.COUT (carry[55]), .SUM (result[54]), .A (A[54]), .B (B[54]), .CIN (C[54]));
FA__1_540 genblk1_53_fa (.COUT (carry[54]), .SUM (result[53]), .A (A[53]), .B (B[53]), .CIN (C[53]));
FA__1_544 genblk1_52_fa (.COUT (carry[53]), .SUM (result[52]), .A (A[52]), .B (B[52]), .CIN (C[52]));
FA__1_548 genblk1_51_fa (.COUT (carry[52]), .SUM (result[51]), .A (A[51]), .B (B[51]), .CIN (C[51]));
FA__1_552 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .B (B[50]), .CIN (C[50]));
FA__1_556 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .B (B[49]), .CIN (C[49]));
FA__1_560 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__1_564 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__1_568 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__1_572 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__1_576 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__1_580 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__1_584 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__1_588 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__1_592 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40])
    , .CIN (C[40]));
FA__1_596 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__1_600 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38])
    , .CIN (C[38]));
FA__1_604 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__1_608 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__1_612 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__1_616 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__1_620 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__1_624 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__1_628 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__1_632 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__1_636 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__1_640 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]), .CIN (C[28]));
FA__1_644 genblk1_27_fa (.COUT (carry[28]), .SUM (result[27]), .A (A[27]), .B (B[27]), .CIN (C[27]));
FA__1_648 genblk1_26_fa (.COUT (carry[27]), .SUM (result[26]), .A (A[26]), .B (B[26]), .CIN (C[26]));
FA__1_652 genblk1_25_fa (.COUT (carry[26]), .SUM (result[25]), .A (A[25]), .B (B[25]));

endmodule //CSAlike__1_753

module FA__1_267 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (CIN), .A2 (B));
XOR2_X1 i_0_0 (.Z (SUM), .A (B), .B (CIN));

endmodule //FA__1_267

module FA__1_271 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_271

module FA__1_275 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_275

module FA__1_279 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_279

module FA__1_283 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_283

module FA__1_287 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_287

module FA__1_291 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_291

module FA__1_295 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_295

module FA__1_299 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_299

module FA__1_303 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_303

module FA__1_307 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_307

module FA__1_311 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_311

module FA__1_315 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_315

module FA__1_319 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_319

module FA__1_323 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_323

module FA__1_327 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_327

module FA__1_331 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire slo__sro_n7;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n7), .A (CIN));
XNOR2_X1 slo__sro_c2 (.ZN (SUM), .A (temp), .B (slo__sro_n7));

endmodule //FA__1_331

module FA__1_335 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_335

module FA__1_339 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_339

module FA__1_343 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_343

module FA__1_347 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_347

module FA__1_351 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_351

module FA__1_355 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_355

module FA__1_359 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_359

module FA__1_363 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_363

module FA__1_367 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_367

module FA__1_371 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;
wire CLOCK_slo__sro_n5;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));
INV_X1 CLOCK_slo__sro_c1 (.ZN (CLOCK_slo__sro_n5), .A (temp));
XNOR2_X1 CLOCK_slo__sro_c2 (.ZN (SUM), .A (CIN), .B (CLOCK_slo__sro_n5));

endmodule //FA__1_371

module FA__1_375 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X2 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X2 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_375

module FA__1_379 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_379

module FA__1_383 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;
wire temp;
wire n_0_0;


INV_X1 i_0_3 (.ZN (COUT), .A (n_0_0));
AOI22_X1 i_0_2 (.ZN (n_0_0), .A1 (A), .A2 (B), .B1 (temp), .B2 (CIN));
XOR2_X1 i_0_1 (.Z (SUM), .A (temp), .B (CIN));
XOR2_X1 i_0_0 (.Z (temp), .A (A), .B (B));

endmodule //FA__1_383

module FA__1_387 (A, B, CIN, SUM, COUT);

output COUT;
output SUM;
input A;
input B;
input CIN;


AND2_X1 i_0_1 (.ZN (COUT), .A1 (B), .A2 (A));
XOR2_X1 i_0_0 (.Z (SUM), .A (A), .B (B));

endmodule //FA__1_387

module CSAlike__1_500 (result, carry, A, B, C);

output [63:0] carry;
output [63:0] result;
input [63:0] A;
input [63:0] B;
input [63:0] C;


FA__1_267 genblk1_58_fa (.COUT (carry[59]), .SUM (result[58]), .B (B[58]), .CIN (C[58]));
FA__1_271 genblk1_57_fa (.COUT (carry[58]), .SUM (result[57]), .A (A[57]), .B (B[57]), .CIN (C[57]));
FA__1_275 genblk1_56_fa (.COUT (carry[57]), .SUM (result[56]), .A (A[56]), .B (B[56]), .CIN (C[56]));
FA__1_279 genblk1_55_fa (.COUT (carry[56]), .SUM (result[55]), .A (A[55]), .B (B[55]), .CIN (C[55]));
FA__1_283 genblk1_54_fa (.COUT (carry[55]), .SUM (result[54]), .A (A[54]), .B (B[54]), .CIN (C[54]));
FA__1_287 genblk1_53_fa (.COUT (carry[54]), .SUM (result[53]), .A (A[53]), .B (B[53]), .CIN (C[53]));
FA__1_291 genblk1_52_fa (.COUT (carry[53]), .SUM (result[52]), .A (A[52]), .B (B[52]), .CIN (C[52]));
FA__1_295 genblk1_51_fa (.COUT (carry[52]), .SUM (result[51]), .A (A[51]), .B (B[51]), .CIN (C[51]));
FA__1_299 genblk1_50_fa (.COUT (carry[51]), .SUM (result[50]), .A (A[50]), .B (B[50]), .CIN (C[50]));
FA__1_303 genblk1_49_fa (.COUT (carry[50]), .SUM (result[49]), .A (A[49]), .B (B[49]), .CIN (C[49]));
FA__1_307 genblk1_48_fa (.COUT (carry[49]), .SUM (result[48]), .A (A[48]), .B (B[48]), .CIN (C[48]));
FA__1_311 genblk1_47_fa (.COUT (carry[48]), .SUM (result[47]), .A (A[47]), .B (B[47]), .CIN (C[47]));
FA__1_315 genblk1_46_fa (.COUT (carry[47]), .SUM (result[46]), .A (A[46]), .B (B[46]), .CIN (C[46]));
FA__1_319 genblk1_45_fa (.COUT (carry[46]), .SUM (result[45]), .A (A[45]), .B (B[45]), .CIN (C[45]));
FA__1_323 genblk1_44_fa (.COUT (carry[45]), .SUM (result[44]), .A (A[44]), .B (B[44]), .CIN (C[44]));
FA__1_327 genblk1_43_fa (.COUT (carry[44]), .SUM (result[43]), .A (A[43]), .B (B[43]), .CIN (C[43]));
FA__1_331 genblk1_42_fa (.COUT (carry[43]), .SUM (result[42]), .A (A[42]), .B (B[42]), .CIN (C[42]));
FA__1_335 genblk1_41_fa (.COUT (carry[42]), .SUM (result[41]), .A (A[41]), .B (B[41]), .CIN (C[41]));
FA__1_339 genblk1_40_fa (.COUT (carry[41]), .SUM (result[40]), .A (A[40]), .B (B[40]), .CIN (C[40]));
FA__1_343 genblk1_39_fa (.COUT (carry[40]), .SUM (result[39]), .A (A[39]), .B (B[39]), .CIN (C[39]));
FA__1_347 genblk1_38_fa (.COUT (carry[39]), .SUM (result[38]), .A (A[38]), .B (B[38]), .CIN (C[38]));
FA__1_351 genblk1_37_fa (.COUT (carry[38]), .SUM (result[37]), .A (A[37]), .B (B[37]), .CIN (C[37]));
FA__1_355 genblk1_36_fa (.COUT (carry[37]), .SUM (result[36]), .A (A[36]), .B (B[36]), .CIN (C[36]));
FA__1_359 genblk1_35_fa (.COUT (carry[36]), .SUM (result[35]), .A (A[35]), .B (B[35]), .CIN (C[35]));
FA__1_363 genblk1_34_fa (.COUT (carry[35]), .SUM (result[34]), .A (A[34]), .B (B[34]), .CIN (C[34]));
FA__1_367 genblk1_33_fa (.COUT (carry[34]), .SUM (result[33]), .A (A[33]), .B (B[33]), .CIN (C[33]));
FA__1_371 genblk1_32_fa (.COUT (carry[33]), .SUM (result[32]), .A (A[32]), .B (B[32]), .CIN (C[32]));
FA__1_375 genblk1_31_fa (.COUT (carry[32]), .SUM (result[31]), .A (A[31]), .B (B[31]), .CIN (C[31]));
FA__1_379 genblk1_30_fa (.COUT (carry[31]), .SUM (result[30]), .A (A[30]), .B (B[30]), .CIN (C[30]));
FA__1_383 genblk1_29_fa (.COUT (carry[30]), .SUM (result[29]), .A (A[29]), .B (B[29]), .CIN (C[29]));
FA__1_387 genblk1_28_fa (.COUT (carry[29]), .SUM (result[28]), .A (A[28]), .B (B[28]));

endmodule //CSAlike__1_500

module addIntermedaiteWires (Res, carry, normalizedWires);

output [63:0] Res;
output [63:0] carry;
input [2047:0] normalizedWires;
wire \intermediateWiresStage1[19][59] ;
wire \intermediateWiresStage1[19][58] ;
wire \intermediateWiresStage1[19][57] ;
wire \intermediateWiresStage1[19][56] ;
wire \intermediateWiresStage1[19][55] ;
wire \intermediateWiresStage1[19][54] ;
wire \intermediateWiresStage1[19][53] ;
wire \intermediateWiresStage1[19][52] ;
wire \intermediateWiresStage1[19][51] ;
wire \intermediateWiresStage1[19][50] ;
wire \intermediateWiresStage1[19][49] ;
wire \intermediateWiresStage1[19][48] ;
wire \intermediateWiresStage1[19][47] ;
wire \intermediateWiresStage1[19][46] ;
wire \intermediateWiresStage1[19][45] ;
wire \intermediateWiresStage1[19][44] ;
wire \intermediateWiresStage1[19][43] ;
wire \intermediateWiresStage1[19][42] ;
wire \intermediateWiresStage1[19][41] ;
wire \intermediateWiresStage1[19][40] ;
wire \intermediateWiresStage1[19][39] ;
wire \intermediateWiresStage1[19][38] ;
wire \intermediateWiresStage1[19][37] ;
wire \intermediateWiresStage1[19][36] ;
wire \intermediateWiresStage1[19][35] ;
wire \intermediateWiresStage1[19][34] ;
wire \intermediateWiresStage1[19][33] ;
wire \intermediateWiresStage1[19][32] ;
wire \intermediateWiresStage1[19][31] ;
wire \intermediateWiresStage1[19][30] ;
wire \intermediateWiresStage1[19][29] ;
wire \intermediateWiresStage1[18][58] ;
wire \intermediateWiresStage1[18][57] ;
wire \intermediateWiresStage1[18][56] ;
wire \intermediateWiresStage1[18][55] ;
wire \intermediateWiresStage1[18][54] ;
wire \intermediateWiresStage1[18][53] ;
wire \intermediateWiresStage1[18][52] ;
wire \intermediateWiresStage1[18][51] ;
wire \intermediateWiresStage1[18][50] ;
wire \intermediateWiresStage1[18][49] ;
wire \intermediateWiresStage1[18][48] ;
wire \intermediateWiresStage1[18][47] ;
wire \intermediateWiresStage1[18][46] ;
wire \intermediateWiresStage1[18][45] ;
wire \intermediateWiresStage1[18][44] ;
wire \intermediateWiresStage1[18][43] ;
wire \intermediateWiresStage1[18][42] ;
wire \intermediateWiresStage1[18][41] ;
wire \intermediateWiresStage1[18][40] ;
wire \intermediateWiresStage1[18][39] ;
wire \intermediateWiresStage1[18][38] ;
wire \intermediateWiresStage1[18][37] ;
wire \intermediateWiresStage1[18][36] ;
wire \intermediateWiresStage1[18][35] ;
wire \intermediateWiresStage1[18][34] ;
wire \intermediateWiresStage1[18][33] ;
wire \intermediateWiresStage1[18][32] ;
wire \intermediateWiresStage1[18][31] ;
wire \intermediateWiresStage1[18][30] ;
wire \intermediateWiresStage1[18][29] ;
wire \intermediateWiresStage1[18][28] ;
wire \intermediateWiresStage1[17][56] ;
wire \intermediateWiresStage1[17][55] ;
wire \intermediateWiresStage1[17][54] ;
wire \intermediateWiresStage1[17][53] ;
wire \intermediateWiresStage1[17][52] ;
wire \intermediateWiresStage1[17][51] ;
wire \intermediateWiresStage1[17][50] ;
wire \intermediateWiresStage1[17][49] ;
wire \intermediateWiresStage1[17][48] ;
wire \intermediateWiresStage1[17][47] ;
wire \intermediateWiresStage1[17][46] ;
wire \intermediateWiresStage1[17][45] ;
wire \intermediateWiresStage1[17][44] ;
wire \intermediateWiresStage1[17][43] ;
wire \intermediateWiresStage1[17][42] ;
wire \intermediateWiresStage1[17][41] ;
wire \intermediateWiresStage1[17][40] ;
wire \intermediateWiresStage1[17][39] ;
wire \intermediateWiresStage1[17][38] ;
wire \intermediateWiresStage1[17][37] ;
wire \intermediateWiresStage1[17][36] ;
wire \intermediateWiresStage1[17][35] ;
wire \intermediateWiresStage1[17][34] ;
wire \intermediateWiresStage1[17][33] ;
wire \intermediateWiresStage1[17][32] ;
wire \intermediateWiresStage1[17][31] ;
wire \intermediateWiresStage1[17][30] ;
wire \intermediateWiresStage1[17][29] ;
wire \intermediateWiresStage1[17][28] ;
wire \intermediateWiresStage1[17][27] ;
wire \intermediateWiresStage1[17][26] ;
wire \intermediateWiresStage1[16][55] ;
wire \intermediateWiresStage1[16][54] ;
wire \intermediateWiresStage1[16][53] ;
wire \intermediateWiresStage1[16][52] ;
wire \intermediateWiresStage1[16][51] ;
wire \intermediateWiresStage1[16][50] ;
wire \intermediateWiresStage1[16][49] ;
wire \intermediateWiresStage1[16][48] ;
wire \intermediateWiresStage1[16][47] ;
wire \intermediateWiresStage1[16][46] ;
wire \intermediateWiresStage1[16][45] ;
wire \intermediateWiresStage1[16][44] ;
wire \intermediateWiresStage1[16][43] ;
wire \intermediateWiresStage1[16][42] ;
wire \intermediateWiresStage1[16][41] ;
wire \intermediateWiresStage1[16][40] ;
wire \intermediateWiresStage1[16][39] ;
wire \intermediateWiresStage1[16][38] ;
wire \intermediateWiresStage1[16][37] ;
wire \intermediateWiresStage1[16][36] ;
wire \intermediateWiresStage1[16][35] ;
wire \intermediateWiresStage1[16][34] ;
wire \intermediateWiresStage1[16][33] ;
wire \intermediateWiresStage1[16][32] ;
wire \intermediateWiresStage1[16][31] ;
wire \intermediateWiresStage1[16][30] ;
wire \intermediateWiresStage1[16][29] ;
wire \intermediateWiresStage1[16][28] ;
wire \intermediateWiresStage1[16][27] ;
wire \intermediateWiresStage1[16][26] ;
wire \intermediateWiresStage1[16][25] ;
wire \intermediateWiresStage1[15][53] ;
wire \intermediateWiresStage1[15][52] ;
wire \intermediateWiresStage1[15][51] ;
wire \intermediateWiresStage1[15][50] ;
wire \intermediateWiresStage1[15][49] ;
wire \intermediateWiresStage1[15][48] ;
wire \intermediateWiresStage1[15][47] ;
wire \intermediateWiresStage1[15][46] ;
wire \intermediateWiresStage1[15][45] ;
wire \intermediateWiresStage1[15][44] ;
wire \intermediateWiresStage1[15][43] ;
wire \intermediateWiresStage1[15][42] ;
wire \intermediateWiresStage1[15][41] ;
wire \intermediateWiresStage1[15][40] ;
wire \intermediateWiresStage1[15][39] ;
wire \intermediateWiresStage1[15][38] ;
wire \intermediateWiresStage1[15][37] ;
wire \intermediateWiresStage1[15][36] ;
wire \intermediateWiresStage1[15][35] ;
wire \intermediateWiresStage1[15][34] ;
wire \intermediateWiresStage1[15][33] ;
wire \intermediateWiresStage1[15][32] ;
wire \intermediateWiresStage1[15][31] ;
wire \intermediateWiresStage1[15][30] ;
wire \intermediateWiresStage1[15][29] ;
wire \intermediateWiresStage1[15][28] ;
wire \intermediateWiresStage1[15][27] ;
wire \intermediateWiresStage1[15][26] ;
wire \intermediateWiresStage1[15][25] ;
wire \intermediateWiresStage1[15][24] ;
wire \intermediateWiresStage1[15][23] ;
wire \intermediateWiresStage1[14][52] ;
wire \intermediateWiresStage1[14][51] ;
wire \intermediateWiresStage1[14][50] ;
wire \intermediateWiresStage1[14][49] ;
wire \intermediateWiresStage1[14][48] ;
wire \intermediateWiresStage1[14][47] ;
wire \intermediateWiresStage1[14][46] ;
wire \intermediateWiresStage1[14][45] ;
wire \intermediateWiresStage1[14][44] ;
wire \intermediateWiresStage1[14][43] ;
wire \intermediateWiresStage1[14][42] ;
wire \intermediateWiresStage1[14][41] ;
wire \intermediateWiresStage1[14][40] ;
wire \intermediateWiresStage1[14][39] ;
wire \intermediateWiresStage1[14][38] ;
wire \intermediateWiresStage1[14][37] ;
wire \intermediateWiresStage1[14][36] ;
wire \intermediateWiresStage1[14][35] ;
wire \intermediateWiresStage1[14][34] ;
wire \intermediateWiresStage1[14][33] ;
wire \intermediateWiresStage1[14][32] ;
wire \intermediateWiresStage1[14][31] ;
wire \intermediateWiresStage1[14][30] ;
wire \intermediateWiresStage1[14][29] ;
wire \intermediateWiresStage1[14][28] ;
wire \intermediateWiresStage1[14][27] ;
wire \intermediateWiresStage1[14][26] ;
wire \intermediateWiresStage1[14][25] ;
wire \intermediateWiresStage1[14][24] ;
wire \intermediateWiresStage1[14][23] ;
wire \intermediateWiresStage1[14][22] ;
wire \intermediateWiresStage1[13][50] ;
wire \intermediateWiresStage1[13][49] ;
wire \intermediateWiresStage1[13][48] ;
wire \intermediateWiresStage1[13][47] ;
wire \intermediateWiresStage1[13][46] ;
wire \intermediateWiresStage1[13][45] ;
wire \intermediateWiresStage1[13][44] ;
wire \intermediateWiresStage1[13][43] ;
wire \intermediateWiresStage1[13][42] ;
wire \intermediateWiresStage1[13][41] ;
wire \intermediateWiresStage1[13][40] ;
wire \intermediateWiresStage1[13][39] ;
wire \intermediateWiresStage1[13][38] ;
wire \intermediateWiresStage1[13][37] ;
wire \intermediateWiresStage1[13][36] ;
wire \intermediateWiresStage1[13][35] ;
wire \intermediateWiresStage1[13][34] ;
wire \intermediateWiresStage1[13][33] ;
wire \intermediateWiresStage1[13][32] ;
wire \intermediateWiresStage1[13][31] ;
wire \intermediateWiresStage1[13][30] ;
wire \intermediateWiresStage1[13][29] ;
wire \intermediateWiresStage1[13][28] ;
wire \intermediateWiresStage1[13][27] ;
wire \intermediateWiresStage1[13][26] ;
wire \intermediateWiresStage1[13][25] ;
wire \intermediateWiresStage1[13][24] ;
wire \intermediateWiresStage1[13][23] ;
wire \intermediateWiresStage1[13][22] ;
wire \intermediateWiresStage1[13][21] ;
wire \intermediateWiresStage1[13][20] ;
wire \intermediateWiresStage1[12][49] ;
wire \intermediateWiresStage1[12][48] ;
wire \intermediateWiresStage1[12][47] ;
wire \intermediateWiresStage1[12][46] ;
wire \intermediateWiresStage1[12][45] ;
wire \intermediateWiresStage1[12][44] ;
wire \intermediateWiresStage1[12][43] ;
wire \intermediateWiresStage1[12][42] ;
wire \intermediateWiresStage1[12][41] ;
wire \intermediateWiresStage1[12][40] ;
wire \intermediateWiresStage1[12][39] ;
wire \intermediateWiresStage1[12][38] ;
wire \intermediateWiresStage1[12][37] ;
wire \intermediateWiresStage1[12][36] ;
wire \intermediateWiresStage1[12][35] ;
wire \intermediateWiresStage1[12][34] ;
wire \intermediateWiresStage1[12][33] ;
wire \intermediateWiresStage1[12][32] ;
wire \intermediateWiresStage1[12][31] ;
wire \intermediateWiresStage1[12][30] ;
wire \intermediateWiresStage1[12][29] ;
wire \intermediateWiresStage1[12][28] ;
wire \intermediateWiresStage1[12][27] ;
wire \intermediateWiresStage1[12][26] ;
wire \intermediateWiresStage1[12][25] ;
wire \intermediateWiresStage1[12][24] ;
wire \intermediateWiresStage1[12][23] ;
wire \intermediateWiresStage1[12][22] ;
wire \intermediateWiresStage1[12][21] ;
wire \intermediateWiresStage1[12][20] ;
wire \intermediateWiresStage1[12][19] ;
wire \intermediateWiresStage1[11][47] ;
wire \intermediateWiresStage1[11][46] ;
wire \intermediateWiresStage1[11][45] ;
wire \intermediateWiresStage1[11][44] ;
wire \intermediateWiresStage1[11][43] ;
wire \intermediateWiresStage1[11][42] ;
wire \intermediateWiresStage1[11][41] ;
wire \intermediateWiresStage1[11][40] ;
wire \intermediateWiresStage1[11][39] ;
wire \intermediateWiresStage1[11][38] ;
wire \intermediateWiresStage1[11][37] ;
wire \intermediateWiresStage1[11][36] ;
wire \intermediateWiresStage1[11][35] ;
wire \intermediateWiresStage1[11][34] ;
wire \intermediateWiresStage1[11][33] ;
wire \intermediateWiresStage1[11][32] ;
wire \intermediateWiresStage1[11][31] ;
wire \intermediateWiresStage1[11][30] ;
wire \intermediateWiresStage1[11][29] ;
wire \intermediateWiresStage1[11][28] ;
wire \intermediateWiresStage1[11][27] ;
wire \intermediateWiresStage1[11][26] ;
wire \intermediateWiresStage1[11][25] ;
wire \intermediateWiresStage1[11][24] ;
wire \intermediateWiresStage1[11][23] ;
wire \intermediateWiresStage1[11][22] ;
wire \intermediateWiresStage1[11][21] ;
wire \intermediateWiresStage1[11][20] ;
wire \intermediateWiresStage1[11][19] ;
wire \intermediateWiresStage1[11][18] ;
wire \intermediateWiresStage1[11][17] ;
wire \intermediateWiresStage1[10][46] ;
wire \intermediateWiresStage1[10][45] ;
wire \intermediateWiresStage1[10][44] ;
wire \intermediateWiresStage1[10][43] ;
wire \intermediateWiresStage1[10][42] ;
wire \intermediateWiresStage1[10][41] ;
wire \intermediateWiresStage1[10][40] ;
wire \intermediateWiresStage1[10][39] ;
wire \intermediateWiresStage1[10][38] ;
wire \intermediateWiresStage1[10][37] ;
wire \intermediateWiresStage1[10][36] ;
wire \intermediateWiresStage1[10][35] ;
wire \intermediateWiresStage1[10][34] ;
wire \intermediateWiresStage1[10][33] ;
wire \intermediateWiresStage1[10][32] ;
wire \intermediateWiresStage1[10][31] ;
wire \intermediateWiresStage1[10][30] ;
wire \intermediateWiresStage1[10][29] ;
wire \intermediateWiresStage1[10][28] ;
wire \intermediateWiresStage1[10][27] ;
wire \intermediateWiresStage1[10][26] ;
wire \intermediateWiresStage1[10][25] ;
wire \intermediateWiresStage1[10][24] ;
wire \intermediateWiresStage1[10][23] ;
wire \intermediateWiresStage1[10][22] ;
wire \intermediateWiresStage1[10][21] ;
wire \intermediateWiresStage1[10][20] ;
wire \intermediateWiresStage1[10][19] ;
wire \intermediateWiresStage1[10][18] ;
wire \intermediateWiresStage1[10][17] ;
wire \intermediateWiresStage1[10][16] ;
wire \intermediateWiresStage1[9][44] ;
wire \intermediateWiresStage1[9][43] ;
wire \intermediateWiresStage1[9][42] ;
wire \intermediateWiresStage1[9][41] ;
wire \intermediateWiresStage1[9][40] ;
wire \intermediateWiresStage1[9][39] ;
wire \intermediateWiresStage1[9][38] ;
wire \intermediateWiresStage1[9][37] ;
wire \intermediateWiresStage1[9][36] ;
wire \intermediateWiresStage1[9][35] ;
wire \intermediateWiresStage1[9][34] ;
wire \intermediateWiresStage1[9][33] ;
wire \intermediateWiresStage1[9][32] ;
wire \intermediateWiresStage1[9][31] ;
wire \intermediateWiresStage1[9][30] ;
wire \intermediateWiresStage1[9][29] ;
wire \intermediateWiresStage1[9][28] ;
wire \intermediateWiresStage1[9][27] ;
wire \intermediateWiresStage1[9][26] ;
wire \intermediateWiresStage1[9][25] ;
wire \intermediateWiresStage1[9][24] ;
wire \intermediateWiresStage1[9][23] ;
wire \intermediateWiresStage1[9][22] ;
wire \intermediateWiresStage1[9][21] ;
wire \intermediateWiresStage1[9][20] ;
wire \intermediateWiresStage1[9][19] ;
wire \intermediateWiresStage1[9][18] ;
wire \intermediateWiresStage1[9][17] ;
wire \intermediateWiresStage1[9][16] ;
wire \intermediateWiresStage1[9][15] ;
wire \intermediateWiresStage1[9][14] ;
wire \intermediateWiresStage1[8][43] ;
wire \intermediateWiresStage1[8][42] ;
wire \intermediateWiresStage1[8][41] ;
wire \intermediateWiresStage1[8][40] ;
wire \intermediateWiresStage1[8][39] ;
wire \intermediateWiresStage1[8][38] ;
wire \intermediateWiresStage1[8][37] ;
wire \intermediateWiresStage1[8][36] ;
wire \intermediateWiresStage1[8][35] ;
wire \intermediateWiresStage1[8][34] ;
wire \intermediateWiresStage1[8][33] ;
wire \intermediateWiresStage1[8][32] ;
wire \intermediateWiresStage1[8][31] ;
wire \intermediateWiresStage1[8][30] ;
wire \intermediateWiresStage1[8][29] ;
wire \intermediateWiresStage1[8][28] ;
wire \intermediateWiresStage1[8][27] ;
wire \intermediateWiresStage1[8][26] ;
wire \intermediateWiresStage1[8][25] ;
wire \intermediateWiresStage1[8][24] ;
wire \intermediateWiresStage1[8][23] ;
wire \intermediateWiresStage1[8][22] ;
wire \intermediateWiresStage1[8][21] ;
wire \intermediateWiresStage1[8][20] ;
wire \intermediateWiresStage1[8][19] ;
wire \intermediateWiresStage1[8][18] ;
wire \intermediateWiresStage1[8][17] ;
wire \intermediateWiresStage1[8][16] ;
wire \intermediateWiresStage1[8][15] ;
wire \intermediateWiresStage1[8][14] ;
wire \intermediateWiresStage1[8][13] ;
wire \intermediateWiresStage1[7][41] ;
wire \intermediateWiresStage1[7][40] ;
wire \intermediateWiresStage1[7][39] ;
wire \intermediateWiresStage1[7][38] ;
wire \intermediateWiresStage1[7][37] ;
wire \intermediateWiresStage1[7][36] ;
wire \intermediateWiresStage1[7][35] ;
wire \intermediateWiresStage1[7][34] ;
wire \intermediateWiresStage1[7][33] ;
wire \intermediateWiresStage1[7][32] ;
wire \intermediateWiresStage1[7][31] ;
wire \intermediateWiresStage1[7][30] ;
wire \intermediateWiresStage1[7][29] ;
wire \intermediateWiresStage1[7][28] ;
wire \intermediateWiresStage1[7][27] ;
wire \intermediateWiresStage1[7][26] ;
wire \intermediateWiresStage1[7][25] ;
wire \intermediateWiresStage1[7][24] ;
wire \intermediateWiresStage1[7][23] ;
wire \intermediateWiresStage1[7][22] ;
wire \intermediateWiresStage1[7][21] ;
wire \intermediateWiresStage1[7][20] ;
wire \intermediateWiresStage1[7][19] ;
wire \intermediateWiresStage1[7][18] ;
wire \intermediateWiresStage1[7][17] ;
wire \intermediateWiresStage1[7][16] ;
wire \intermediateWiresStage1[7][15] ;
wire \intermediateWiresStage1[7][14] ;
wire \intermediateWiresStage1[7][13] ;
wire \intermediateWiresStage1[7][12] ;
wire \intermediateWiresStage1[7][11] ;
wire \intermediateWiresStage1[6][40] ;
wire \intermediateWiresStage1[6][39] ;
wire \intermediateWiresStage1[6][38] ;
wire \intermediateWiresStage1[6][37] ;
wire \intermediateWiresStage1[6][36] ;
wire \intermediateWiresStage1[6][35] ;
wire \intermediateWiresStage1[6][34] ;
wire \intermediateWiresStage1[6][33] ;
wire \intermediateWiresStage1[6][32] ;
wire \intermediateWiresStage1[6][31] ;
wire \intermediateWiresStage1[6][30] ;
wire \intermediateWiresStage1[6][29] ;
wire \intermediateWiresStage1[6][28] ;
wire \intermediateWiresStage1[6][27] ;
wire \intermediateWiresStage1[6][26] ;
wire \intermediateWiresStage1[6][25] ;
wire \intermediateWiresStage1[6][24] ;
wire \intermediateWiresStage1[6][23] ;
wire \intermediateWiresStage1[6][22] ;
wire \intermediateWiresStage1[6][21] ;
wire \intermediateWiresStage1[6][20] ;
wire \intermediateWiresStage1[6][19] ;
wire \intermediateWiresStage1[6][18] ;
wire \intermediateWiresStage1[6][17] ;
wire \intermediateWiresStage1[6][16] ;
wire \intermediateWiresStage1[6][15] ;
wire \intermediateWiresStage1[6][14] ;
wire \intermediateWiresStage1[6][13] ;
wire \intermediateWiresStage1[6][12] ;
wire \intermediateWiresStage1[6][11] ;
wire \intermediateWiresStage1[6][10] ;
wire \intermediateWiresStage1[5][38] ;
wire \intermediateWiresStage1[5][37] ;
wire \intermediateWiresStage1[5][36] ;
wire \intermediateWiresStage1[5][35] ;
wire \intermediateWiresStage1[5][34] ;
wire \intermediateWiresStage1[5][33] ;
wire \intermediateWiresStage1[5][32] ;
wire \intermediateWiresStage1[5][31] ;
wire \intermediateWiresStage1[5][30] ;
wire \intermediateWiresStage1[5][29] ;
wire \intermediateWiresStage1[5][28] ;
wire \intermediateWiresStage1[5][27] ;
wire \intermediateWiresStage1[5][26] ;
wire \intermediateWiresStage1[5][25] ;
wire \intermediateWiresStage1[5][24] ;
wire \intermediateWiresStage1[5][23] ;
wire \intermediateWiresStage1[5][22] ;
wire \intermediateWiresStage1[5][21] ;
wire \intermediateWiresStage1[5][20] ;
wire \intermediateWiresStage1[5][19] ;
wire \intermediateWiresStage1[5][18] ;
wire \intermediateWiresStage1[5][17] ;
wire \intermediateWiresStage1[5][16] ;
wire \intermediateWiresStage1[5][15] ;
wire \intermediateWiresStage1[5][14] ;
wire \intermediateWiresStage1[5][13] ;
wire \intermediateWiresStage1[5][12] ;
wire \intermediateWiresStage1[5][11] ;
wire \intermediateWiresStage1[5][10] ;
wire \intermediateWiresStage1[5][9] ;
wire \intermediateWiresStage1[5][8] ;
wire \intermediateWiresStage1[4][37] ;
wire \intermediateWiresStage1[4][36] ;
wire \intermediateWiresStage1[4][35] ;
wire \intermediateWiresStage1[4][34] ;
wire \intermediateWiresStage1[4][33] ;
wire \intermediateWiresStage1[4][32] ;
wire \intermediateWiresStage1[4][31] ;
wire \intermediateWiresStage1[4][30] ;
wire \intermediateWiresStage1[4][29] ;
wire \intermediateWiresStage1[4][28] ;
wire \intermediateWiresStage1[4][27] ;
wire \intermediateWiresStage1[4][26] ;
wire \intermediateWiresStage1[4][25] ;
wire \intermediateWiresStage1[4][24] ;
wire \intermediateWiresStage1[4][23] ;
wire \intermediateWiresStage1[4][22] ;
wire \intermediateWiresStage1[4][21] ;
wire \intermediateWiresStage1[4][20] ;
wire \intermediateWiresStage1[4][19] ;
wire \intermediateWiresStage1[4][18] ;
wire \intermediateWiresStage1[4][17] ;
wire \intermediateWiresStage1[4][16] ;
wire \intermediateWiresStage1[4][15] ;
wire \intermediateWiresStage1[4][14] ;
wire \intermediateWiresStage1[4][13] ;
wire \intermediateWiresStage1[4][12] ;
wire \intermediateWiresStage1[4][11] ;
wire \intermediateWiresStage1[4][10] ;
wire \intermediateWiresStage1[4][9] ;
wire \intermediateWiresStage1[4][8] ;
wire \intermediateWiresStage1[4][7] ;
wire \intermediateWiresStage1[3][35] ;
wire \intermediateWiresStage1[3][34] ;
wire \intermediateWiresStage1[3][33] ;
wire \intermediateWiresStage1[3][32] ;
wire \intermediateWiresStage1[3][31] ;
wire \intermediateWiresStage1[3][30] ;
wire \intermediateWiresStage1[3][29] ;
wire \intermediateWiresStage1[3][28] ;
wire \intermediateWiresStage1[3][27] ;
wire \intermediateWiresStage1[3][26] ;
wire \intermediateWiresStage1[3][25] ;
wire \intermediateWiresStage1[3][24] ;
wire \intermediateWiresStage1[3][23] ;
wire \intermediateWiresStage1[3][22] ;
wire \intermediateWiresStage1[3][21] ;
wire \intermediateWiresStage1[3][20] ;
wire \intermediateWiresStage1[3][19] ;
wire \intermediateWiresStage1[3][18] ;
wire \intermediateWiresStage1[3][17] ;
wire \intermediateWiresStage1[3][16] ;
wire \intermediateWiresStage1[3][15] ;
wire \intermediateWiresStage1[3][14] ;
wire \intermediateWiresStage1[3][13] ;
wire \intermediateWiresStage1[3][12] ;
wire \intermediateWiresStage1[3][11] ;
wire \intermediateWiresStage1[3][10] ;
wire \intermediateWiresStage1[3][9] ;
wire \intermediateWiresStage1[3][8] ;
wire \intermediateWiresStage1[3][7] ;
wire \intermediateWiresStage1[3][6] ;
wire \intermediateWiresStage1[3][5] ;
wire \intermediateWiresStage1[2][34] ;
wire \intermediateWiresStage1[2][33] ;
wire \intermediateWiresStage1[2][32] ;
wire \intermediateWiresStage1[2][31] ;
wire \intermediateWiresStage1[2][30] ;
wire \intermediateWiresStage1[2][29] ;
wire \intermediateWiresStage1[2][28] ;
wire \intermediateWiresStage1[2][27] ;
wire \intermediateWiresStage1[2][26] ;
wire \intermediateWiresStage1[2][25] ;
wire \intermediateWiresStage1[2][24] ;
wire \intermediateWiresStage1[2][23] ;
wire \intermediateWiresStage1[2][22] ;
wire \intermediateWiresStage1[2][21] ;
wire \intermediateWiresStage1[2][20] ;
wire \intermediateWiresStage1[2][19] ;
wire \intermediateWiresStage1[2][18] ;
wire \intermediateWiresStage1[2][17] ;
wire \intermediateWiresStage1[2][16] ;
wire \intermediateWiresStage1[2][15] ;
wire \intermediateWiresStage1[2][14] ;
wire \intermediateWiresStage1[2][13] ;
wire \intermediateWiresStage1[2][12] ;
wire \intermediateWiresStage1[2][11] ;
wire \intermediateWiresStage1[2][10] ;
wire \intermediateWiresStage1[2][9] ;
wire \intermediateWiresStage1[2][8] ;
wire \intermediateWiresStage1[2][7] ;
wire \intermediateWiresStage1[2][6] ;
wire \intermediateWiresStage1[2][5] ;
wire \intermediateWiresStage1[2][4] ;
wire \intermediateWiresStage1[1][32] ;
wire \intermediateWiresStage1[1][31] ;
wire \intermediateWiresStage1[1][30] ;
wire \intermediateWiresStage1[1][29] ;
wire \intermediateWiresStage1[1][28] ;
wire \intermediateWiresStage1[1][27] ;
wire \intermediateWiresStage1[1][26] ;
wire \intermediateWiresStage1[1][25] ;
wire \intermediateWiresStage1[1][24] ;
wire \intermediateWiresStage1[1][23] ;
wire \intermediateWiresStage1[1][22] ;
wire \intermediateWiresStage1[1][21] ;
wire \intermediateWiresStage1[1][20] ;
wire \intermediateWiresStage1[1][19] ;
wire \intermediateWiresStage1[1][18] ;
wire \intermediateWiresStage1[1][17] ;
wire \intermediateWiresStage1[1][16] ;
wire \intermediateWiresStage1[1][15] ;
wire \intermediateWiresStage1[1][14] ;
wire \intermediateWiresStage1[1][13] ;
wire \intermediateWiresStage1[1][12] ;
wire \intermediateWiresStage1[1][11] ;
wire \intermediateWiresStage1[1][10] ;
wire \intermediateWiresStage1[1][9] ;
wire \intermediateWiresStage1[1][8] ;
wire \intermediateWiresStage1[1][7] ;
wire \intermediateWiresStage1[1][6] ;
wire \intermediateWiresStage1[1][5] ;
wire \intermediateWiresStage1[1][4] ;
wire \intermediateWiresStage1[1][3] ;
wire \intermediateWiresStage1[1][2] ;
wire \intermediateWiresStage1[0][31] ;
wire \intermediateWiresStage1[0][30] ;
wire \intermediateWiresStage1[0][29] ;
wire \intermediateWiresStage1[0][28] ;
wire \intermediateWiresStage1[0][27] ;
wire \intermediateWiresStage1[0][26] ;
wire \intermediateWiresStage1[0][25] ;
wire \intermediateWiresStage1[0][24] ;
wire \intermediateWiresStage1[0][23] ;
wire \intermediateWiresStage1[0][22] ;
wire \intermediateWiresStage1[0][21] ;
wire \intermediateWiresStage1[0][20] ;
wire \intermediateWiresStage1[0][19] ;
wire \intermediateWiresStage1[0][18] ;
wire \intermediateWiresStage1[0][17] ;
wire \intermediateWiresStage1[0][16] ;
wire \intermediateWiresStage1[0][15] ;
wire \intermediateWiresStage1[0][14] ;
wire \intermediateWiresStage1[0][13] ;
wire \intermediateWiresStage1[0][12] ;
wire \intermediateWiresStage1[0][11] ;
wire \intermediateWiresStage1[0][10] ;
wire \intermediateWiresStage1[0][9] ;
wire \intermediateWiresStage1[0][8] ;
wire \intermediateWiresStage1[0][7] ;
wire \intermediateWiresStage1[0][6] ;
wire \intermediateWiresStage1[0][5] ;
wire \intermediateWiresStage1[0][4] ;
wire \intermediateWiresStage1[0][3] ;
wire \intermediateWiresStage1[0][2] ;
wire \intermediateWiresStage2[13][60] ;
wire \intermediateWiresStage2[13][59] ;
wire \intermediateWiresStage2[13][58] ;
wire \intermediateWiresStage2[13][57] ;
wire \intermediateWiresStage2[13][56] ;
wire \intermediateWiresStage2[13][55] ;
wire \intermediateWiresStage2[13][54] ;
wire \intermediateWiresStage2[13][53] ;
wire \intermediateWiresStage2[13][52] ;
wire \intermediateWiresStage2[13][51] ;
wire \intermediateWiresStage2[13][50] ;
wire \intermediateWiresStage2[13][49] ;
wire \intermediateWiresStage2[13][48] ;
wire \intermediateWiresStage2[13][47] ;
wire \intermediateWiresStage2[13][46] ;
wire \intermediateWiresStage2[13][45] ;
wire \intermediateWiresStage2[13][44] ;
wire \intermediateWiresStage2[13][43] ;
wire \intermediateWiresStage2[13][42] ;
wire \intermediateWiresStage2[13][41] ;
wire \intermediateWiresStage2[13][40] ;
wire \intermediateWiresStage2[13][39] ;
wire \intermediateWiresStage2[13][38] ;
wire \intermediateWiresStage2[13][37] ;
wire \intermediateWiresStage2[13][36] ;
wire \intermediateWiresStage2[13][35] ;
wire \intermediateWiresStage2[13][34] ;
wire \intermediateWiresStage2[13][33] ;
wire \intermediateWiresStage2[13][32] ;
wire \intermediateWiresStage2[13][31] ;
wire \intermediateWiresStage2[13][30] ;
wire \intermediateWiresStage2[12][59] ;
wire \intermediateWiresStage2[12][58] ;
wire \intermediateWiresStage2[12][57] ;
wire \intermediateWiresStage2[12][56] ;
wire \intermediateWiresStage2[12][55] ;
wire \intermediateWiresStage2[12][54] ;
wire \intermediateWiresStage2[12][53] ;
wire \intermediateWiresStage2[12][52] ;
wire \intermediateWiresStage2[12][51] ;
wire \intermediateWiresStage2[12][50] ;
wire \intermediateWiresStage2[12][49] ;
wire \intermediateWiresStage2[12][48] ;
wire \intermediateWiresStage2[12][47] ;
wire \intermediateWiresStage2[12][46] ;
wire \intermediateWiresStage2[12][45] ;
wire \intermediateWiresStage2[12][44] ;
wire \intermediateWiresStage2[12][43] ;
wire \intermediateWiresStage2[12][42] ;
wire \intermediateWiresStage2[12][41] ;
wire \intermediateWiresStage2[12][40] ;
wire \intermediateWiresStage2[12][39] ;
wire \intermediateWiresStage2[12][38] ;
wire \intermediateWiresStage2[12][37] ;
wire \intermediateWiresStage2[12][36] ;
wire \intermediateWiresStage2[12][35] ;
wire \intermediateWiresStage2[12][34] ;
wire \intermediateWiresStage2[12][33] ;
wire \intermediateWiresStage2[12][32] ;
wire \intermediateWiresStage2[12][31] ;
wire \intermediateWiresStage2[12][30] ;
wire \intermediateWiresStage2[12][29] ;
wire \intermediateWiresStage2[11][57] ;
wire \intermediateWiresStage2[11][56] ;
wire \intermediateWiresStage2[11][55] ;
wire \intermediateWiresStage2[11][54] ;
wire \intermediateWiresStage2[11][53] ;
wire \intermediateWiresStage2[11][52] ;
wire \intermediateWiresStage2[11][51] ;
wire \intermediateWiresStage2[11][50] ;
wire \intermediateWiresStage2[11][49] ;
wire \intermediateWiresStage2[11][48] ;
wire \intermediateWiresStage2[11][47] ;
wire \intermediateWiresStage2[11][46] ;
wire \intermediateWiresStage2[11][45] ;
wire \intermediateWiresStage2[11][44] ;
wire \intermediateWiresStage2[11][43] ;
wire \intermediateWiresStage2[11][42] ;
wire \intermediateWiresStage2[11][41] ;
wire \intermediateWiresStage2[11][40] ;
wire \intermediateWiresStage2[11][39] ;
wire \intermediateWiresStage2[11][38] ;
wire \intermediateWiresStage2[11][37] ;
wire \intermediateWiresStage2[11][36] ;
wire \intermediateWiresStage2[11][35] ;
wire \intermediateWiresStage2[11][34] ;
wire \intermediateWiresStage2[11][33] ;
wire \intermediateWiresStage2[11][32] ;
wire \intermediateWiresStage2[11][31] ;
wire \intermediateWiresStage2[11][30] ;
wire \intermediateWiresStage2[11][29] ;
wire \intermediateWiresStage2[11][28] ;
wire \intermediateWiresStage2[11][27] ;
wire \intermediateWiresStage2[11][26] ;
wire \intermediateWiresStage2[11][25] ;
wire \intermediateWiresStage2[10][56] ;
wire \intermediateWiresStage2[10][55] ;
wire \intermediateWiresStage2[10][54] ;
wire \intermediateWiresStage2[10][53] ;
wire \intermediateWiresStage2[10][52] ;
wire \intermediateWiresStage2[10][51] ;
wire \intermediateWiresStage2[10][50] ;
wire \intermediateWiresStage2[10][49] ;
wire \intermediateWiresStage2[10][48] ;
wire \intermediateWiresStage2[10][47] ;
wire \intermediateWiresStage2[10][46] ;
wire \intermediateWiresStage2[10][45] ;
wire \intermediateWiresStage2[10][44] ;
wire \intermediateWiresStage2[10][43] ;
wire \intermediateWiresStage2[10][42] ;
wire \intermediateWiresStage2[10][41] ;
wire \intermediateWiresStage2[10][40] ;
wire \intermediateWiresStage2[10][39] ;
wire \intermediateWiresStage2[10][38] ;
wire \intermediateWiresStage2[10][37] ;
wire \intermediateWiresStage2[10][36] ;
wire \intermediateWiresStage2[10][35] ;
wire \intermediateWiresStage2[10][34] ;
wire \intermediateWiresStage2[10][33] ;
wire \intermediateWiresStage2[10][32] ;
wire \intermediateWiresStage2[10][31] ;
wire \intermediateWiresStage2[10][30] ;
wire \intermediateWiresStage2[10][29] ;
wire \intermediateWiresStage2[10][28] ;
wire \intermediateWiresStage2[10][27] ;
wire \intermediateWiresStage2[10][26] ;
wire \intermediateWiresStage2[10][25] ;
wire \intermediateWiresStage2[10][24] ;
wire \intermediateWiresStage2[9][51] ;
wire \intermediateWiresStage2[9][50] ;
wire \intermediateWiresStage2[9][49] ;
wire \intermediateWiresStage2[9][48] ;
wire \intermediateWiresStage2[9][47] ;
wire \intermediateWiresStage2[9][46] ;
wire \intermediateWiresStage2[9][45] ;
wire \intermediateWiresStage2[9][44] ;
wire \intermediateWiresStage2[9][43] ;
wire \intermediateWiresStage2[9][42] ;
wire \intermediateWiresStage2[9][41] ;
wire \intermediateWiresStage2[9][40] ;
wire \intermediateWiresStage2[9][39] ;
wire \intermediateWiresStage2[9][38] ;
wire \intermediateWiresStage2[9][37] ;
wire \intermediateWiresStage2[9][36] ;
wire \intermediateWiresStage2[9][35] ;
wire \intermediateWiresStage2[9][34] ;
wire \intermediateWiresStage2[9][33] ;
wire \intermediateWiresStage2[9][32] ;
wire \intermediateWiresStage2[9][31] ;
wire \intermediateWiresStage2[9][30] ;
wire \intermediateWiresStage2[9][29] ;
wire \intermediateWiresStage2[9][28] ;
wire \intermediateWiresStage2[9][27] ;
wire \intermediateWiresStage2[9][26] ;
wire \intermediateWiresStage2[9][25] ;
wire \intermediateWiresStage2[9][24] ;
wire \intermediateWiresStage2[9][23] ;
wire \intermediateWiresStage2[9][22] ;
wire \intermediateWiresStage2[9][21] ;
wire \intermediateWiresStage2[8][50] ;
wire \intermediateWiresStage2[8][49] ;
wire \intermediateWiresStage2[8][48] ;
wire \intermediateWiresStage2[8][47] ;
wire \intermediateWiresStage2[8][46] ;
wire \intermediateWiresStage2[8][45] ;
wire \intermediateWiresStage2[8][44] ;
wire \intermediateWiresStage2[8][43] ;
wire \intermediateWiresStage2[8][42] ;
wire \intermediateWiresStage2[8][41] ;
wire \intermediateWiresStage2[8][40] ;
wire \intermediateWiresStage2[8][39] ;
wire \intermediateWiresStage2[8][38] ;
wire \intermediateWiresStage2[8][37] ;
wire \intermediateWiresStage2[8][36] ;
wire \intermediateWiresStage2[8][35] ;
wire \intermediateWiresStage2[8][34] ;
wire \intermediateWiresStage2[8][33] ;
wire \intermediateWiresStage2[8][32] ;
wire \intermediateWiresStage2[8][31] ;
wire \intermediateWiresStage2[8][30] ;
wire \intermediateWiresStage2[8][29] ;
wire \intermediateWiresStage2[8][28] ;
wire \intermediateWiresStage2[8][27] ;
wire \intermediateWiresStage2[8][26] ;
wire \intermediateWiresStage2[8][25] ;
wire \intermediateWiresStage2[8][24] ;
wire \intermediateWiresStage2[8][23] ;
wire \intermediateWiresStage2[8][22] ;
wire \intermediateWiresStage2[8][21] ;
wire \intermediateWiresStage2[8][20] ;
wire \intermediateWiresStage2[7][48] ;
wire \intermediateWiresStage2[7][47] ;
wire \intermediateWiresStage2[7][46] ;
wire \intermediateWiresStage2[7][45] ;
wire \intermediateWiresStage2[7][44] ;
wire \intermediateWiresStage2[7][43] ;
wire \intermediateWiresStage2[7][42] ;
wire \intermediateWiresStage2[7][41] ;
wire \intermediateWiresStage2[7][40] ;
wire \intermediateWiresStage2[7][39] ;
wire \intermediateWiresStage2[7][38] ;
wire \intermediateWiresStage2[7][37] ;
wire \intermediateWiresStage2[7][36] ;
wire \intermediateWiresStage2[7][35] ;
wire \intermediateWiresStage2[7][34] ;
wire \intermediateWiresStage2[7][33] ;
wire \intermediateWiresStage2[7][32] ;
wire \intermediateWiresStage2[7][31] ;
wire \intermediateWiresStage2[7][30] ;
wire \intermediateWiresStage2[7][29] ;
wire \intermediateWiresStage2[7][28] ;
wire \intermediateWiresStage2[7][27] ;
wire \intermediateWiresStage2[7][26] ;
wire \intermediateWiresStage2[7][25] ;
wire \intermediateWiresStage2[7][24] ;
wire \intermediateWiresStage2[7][23] ;
wire \intermediateWiresStage2[7][22] ;
wire \intermediateWiresStage2[7][21] ;
wire \intermediateWiresStage2[7][20] ;
wire \intermediateWiresStage2[7][19] ;
wire \intermediateWiresStage2[7][18] ;
wire \intermediateWiresStage2[7][17] ;
wire \intermediateWiresStage2[7][16] ;
wire \intermediateWiresStage2[6][47] ;
wire \intermediateWiresStage2[6][46] ;
wire \intermediateWiresStage2[6][45] ;
wire \intermediateWiresStage2[6][44] ;
wire \intermediateWiresStage2[6][43] ;
wire \intermediateWiresStage2[6][42] ;
wire \intermediateWiresStage2[6][41] ;
wire \intermediateWiresStage2[6][40] ;
wire \intermediateWiresStage2[6][39] ;
wire \intermediateWiresStage2[6][38] ;
wire \intermediateWiresStage2[6][37] ;
wire \intermediateWiresStage2[6][36] ;
wire \intermediateWiresStage2[6][35] ;
wire \intermediateWiresStage2[6][34] ;
wire \intermediateWiresStage2[6][33] ;
wire \intermediateWiresStage2[6][32] ;
wire \intermediateWiresStage2[6][31] ;
wire \intermediateWiresStage2[6][30] ;
wire \intermediateWiresStage2[6][29] ;
wire \intermediateWiresStage2[6][28] ;
wire \intermediateWiresStage2[6][27] ;
wire \intermediateWiresStage2[6][26] ;
wire \intermediateWiresStage2[6][25] ;
wire \intermediateWiresStage2[6][24] ;
wire \intermediateWiresStage2[6][23] ;
wire \intermediateWiresStage2[6][22] ;
wire \intermediateWiresStage2[6][21] ;
wire \intermediateWiresStage2[6][20] ;
wire \intermediateWiresStage2[6][19] ;
wire \intermediateWiresStage2[6][18] ;
wire \intermediateWiresStage2[6][17] ;
wire \intermediateWiresStage2[6][16] ;
wire \intermediateWiresStage2[6][15] ;
wire \intermediateWiresStage2[5][42] ;
wire \intermediateWiresStage2[5][41] ;
wire \intermediateWiresStage2[5][40] ;
wire \intermediateWiresStage2[5][39] ;
wire \intermediateWiresStage2[5][38] ;
wire \intermediateWiresStage2[5][37] ;
wire \intermediateWiresStage2[5][36] ;
wire \intermediateWiresStage2[5][35] ;
wire \intermediateWiresStage2[5][34] ;
wire \intermediateWiresStage2[5][33] ;
wire \intermediateWiresStage2[5][32] ;
wire \intermediateWiresStage2[5][31] ;
wire \intermediateWiresStage2[5][30] ;
wire \intermediateWiresStage2[5][29] ;
wire \intermediateWiresStage2[5][28] ;
wire \intermediateWiresStage2[5][27] ;
wire \intermediateWiresStage2[5][26] ;
wire \intermediateWiresStage2[5][25] ;
wire \intermediateWiresStage2[5][24] ;
wire \intermediateWiresStage2[5][23] ;
wire \intermediateWiresStage2[5][22] ;
wire \intermediateWiresStage2[5][21] ;
wire \intermediateWiresStage2[5][20] ;
wire \intermediateWiresStage2[5][19] ;
wire \intermediateWiresStage2[5][18] ;
wire \intermediateWiresStage2[5][17] ;
wire \intermediateWiresStage2[5][16] ;
wire \intermediateWiresStage2[5][15] ;
wire \intermediateWiresStage2[5][14] ;
wire \intermediateWiresStage2[5][13] ;
wire \intermediateWiresStage2[5][12] ;
wire \intermediateWiresStage2[4][41] ;
wire \intermediateWiresStage2[4][40] ;
wire \intermediateWiresStage2[4][39] ;
wire \intermediateWiresStage2[4][38] ;
wire \intermediateWiresStage2[4][37] ;
wire \intermediateWiresStage2[4][36] ;
wire \intermediateWiresStage2[4][35] ;
wire \intermediateWiresStage2[4][34] ;
wire \intermediateWiresStage2[4][33] ;
wire \intermediateWiresStage2[4][32] ;
wire \intermediateWiresStage2[4][31] ;
wire \intermediateWiresStage2[4][30] ;
wire \intermediateWiresStage2[4][29] ;
wire \intermediateWiresStage2[4][28] ;
wire \intermediateWiresStage2[4][27] ;
wire \intermediateWiresStage2[4][26] ;
wire \intermediateWiresStage2[4][25] ;
wire \intermediateWiresStage2[4][24] ;
wire \intermediateWiresStage2[4][23] ;
wire \intermediateWiresStage2[4][22] ;
wire \intermediateWiresStage2[4][21] ;
wire \intermediateWiresStage2[4][20] ;
wire \intermediateWiresStage2[4][19] ;
wire \intermediateWiresStage2[4][18] ;
wire \intermediateWiresStage2[4][17] ;
wire \intermediateWiresStage2[4][16] ;
wire \intermediateWiresStage2[4][15] ;
wire \intermediateWiresStage2[4][14] ;
wire \intermediateWiresStage2[4][13] ;
wire \intermediateWiresStage2[4][12] ;
wire \intermediateWiresStage2[4][11] ;
wire \intermediateWiresStage2[3][39] ;
wire \intermediateWiresStage2[3][38] ;
wire \intermediateWiresStage2[3][37] ;
wire \intermediateWiresStage2[3][36] ;
wire \intermediateWiresStage2[3][35] ;
wire \intermediateWiresStage2[3][34] ;
wire \intermediateWiresStage2[3][33] ;
wire \intermediateWiresStage2[3][32] ;
wire \intermediateWiresStage2[3][31] ;
wire \intermediateWiresStage2[3][30] ;
wire \intermediateWiresStage2[3][29] ;
wire \intermediateWiresStage2[3][28] ;
wire \intermediateWiresStage2[3][27] ;
wire \intermediateWiresStage2[3][26] ;
wire \intermediateWiresStage2[3][25] ;
wire \intermediateWiresStage2[3][24] ;
wire \intermediateWiresStage2[3][23] ;
wire \intermediateWiresStage2[3][22] ;
wire \intermediateWiresStage2[3][21] ;
wire \intermediateWiresStage2[3][20] ;
wire \intermediateWiresStage2[3][19] ;
wire \intermediateWiresStage2[3][18] ;
wire \intermediateWiresStage2[3][17] ;
wire \intermediateWiresStage2[3][16] ;
wire \intermediateWiresStage2[3][15] ;
wire \intermediateWiresStage2[3][14] ;
wire \intermediateWiresStage2[3][13] ;
wire \intermediateWiresStage2[3][12] ;
wire \intermediateWiresStage2[3][11] ;
wire \intermediateWiresStage2[3][10] ;
wire \intermediateWiresStage2[3][9] ;
wire \intermediateWiresStage2[3][8] ;
wire \intermediateWiresStage2[3][7] ;
wire \intermediateWiresStage2[2][38] ;
wire \intermediateWiresStage2[2][37] ;
wire \intermediateWiresStage2[2][36] ;
wire \intermediateWiresStage2[2][35] ;
wire \intermediateWiresStage2[2][34] ;
wire \intermediateWiresStage2[2][33] ;
wire \intermediateWiresStage2[2][32] ;
wire \intermediateWiresStage2[2][31] ;
wire \intermediateWiresStage2[2][30] ;
wire \intermediateWiresStage2[2][29] ;
wire \intermediateWiresStage2[2][28] ;
wire \intermediateWiresStage2[2][27] ;
wire \intermediateWiresStage2[2][26] ;
wire \intermediateWiresStage2[2][25] ;
wire \intermediateWiresStage2[2][24] ;
wire \intermediateWiresStage2[2][23] ;
wire \intermediateWiresStage2[2][22] ;
wire \intermediateWiresStage2[2][21] ;
wire \intermediateWiresStage2[2][20] ;
wire \intermediateWiresStage2[2][19] ;
wire \intermediateWiresStage2[2][18] ;
wire \intermediateWiresStage2[2][17] ;
wire \intermediateWiresStage2[2][16] ;
wire \intermediateWiresStage2[2][15] ;
wire \intermediateWiresStage2[2][14] ;
wire \intermediateWiresStage2[2][13] ;
wire \intermediateWiresStage2[2][12] ;
wire \intermediateWiresStage2[2][11] ;
wire \intermediateWiresStage2[2][10] ;
wire \intermediateWiresStage2[2][9] ;
wire \intermediateWiresStage2[2][8] ;
wire \intermediateWiresStage2[2][7] ;
wire \intermediateWiresStage2[2][6] ;
wire \intermediateWiresStage2[1][33] ;
wire \intermediateWiresStage2[1][32] ;
wire \intermediateWiresStage2[1][31] ;
wire \intermediateWiresStage2[1][30] ;
wire \intermediateWiresStage2[1][29] ;
wire \intermediateWiresStage2[1][28] ;
wire \intermediateWiresStage2[1][27] ;
wire \intermediateWiresStage2[1][26] ;
wire \intermediateWiresStage2[1][25] ;
wire \intermediateWiresStage2[1][24] ;
wire \intermediateWiresStage2[1][23] ;
wire \intermediateWiresStage2[1][22] ;
wire \intermediateWiresStage2[1][21] ;
wire \intermediateWiresStage2[1][20] ;
wire \intermediateWiresStage2[1][19] ;
wire \intermediateWiresStage2[1][18] ;
wire \intermediateWiresStage2[1][17] ;
wire \intermediateWiresStage2[1][16] ;
wire \intermediateWiresStage2[1][15] ;
wire \intermediateWiresStage2[1][14] ;
wire \intermediateWiresStage2[1][13] ;
wire \intermediateWiresStage2[1][12] ;
wire \intermediateWiresStage2[1][11] ;
wire \intermediateWiresStage2[1][10] ;
wire \intermediateWiresStage2[1][9] ;
wire \intermediateWiresStage2[1][8] ;
wire \intermediateWiresStage2[1][7] ;
wire \intermediateWiresStage2[1][6] ;
wire \intermediateWiresStage2[1][5] ;
wire \intermediateWiresStage2[1][4] ;
wire \intermediateWiresStage2[1][3] ;
wire \intermediateWiresStage2[0][32] ;
wire \intermediateWiresStage2[0][31] ;
wire \intermediateWiresStage2[0][30] ;
wire \intermediateWiresStage2[0][29] ;
wire \intermediateWiresStage2[0][28] ;
wire \intermediateWiresStage2[0][27] ;
wire \intermediateWiresStage2[0][26] ;
wire \intermediateWiresStage2[0][25] ;
wire \intermediateWiresStage2[0][24] ;
wire \intermediateWiresStage2[0][23] ;
wire \intermediateWiresStage2[0][22] ;
wire \intermediateWiresStage2[0][21] ;
wire \intermediateWiresStage2[0][20] ;
wire \intermediateWiresStage2[0][19] ;
wire \intermediateWiresStage2[0][18] ;
wire \intermediateWiresStage2[0][17] ;
wire \intermediateWiresStage2[0][16] ;
wire \intermediateWiresStage2[0][15] ;
wire \intermediateWiresStage2[0][14] ;
wire \intermediateWiresStage2[0][13] ;
wire \intermediateWiresStage2[0][12] ;
wire \intermediateWiresStage2[0][11] ;
wire \intermediateWiresStage2[0][10] ;
wire \intermediateWiresStage2[0][9] ;
wire \intermediateWiresStage2[0][8] ;
wire \intermediateWiresStage2[0][7] ;
wire \intermediateWiresStage2[0][6] ;
wire \intermediateWiresStage2[0][5] ;
wire \intermediateWiresStage2[0][4] ;
wire \intermediateWiresStage2[0][3] ;
wire \intermediateWiresStage3[9][61] ;
wire \intermediateWiresStage3[9][60] ;
wire \intermediateWiresStage3[9][59] ;
wire \intermediateWiresStage3[9][58] ;
wire \intermediateWiresStage3[9][57] ;
wire \intermediateWiresStage3[9][56] ;
wire \intermediateWiresStage3[9][55] ;
wire \intermediateWiresStage3[9][54] ;
wire \intermediateWiresStage3[9][53] ;
wire \intermediateWiresStage3[9][52] ;
wire \intermediateWiresStage3[9][51] ;
wire \intermediateWiresStage3[9][50] ;
wire \intermediateWiresStage3[9][49] ;
wire \intermediateWiresStage3[9][48] ;
wire \intermediateWiresStage3[9][47] ;
wire \intermediateWiresStage3[9][46] ;
wire \intermediateWiresStage3[9][45] ;
wire \intermediateWiresStage3[9][44] ;
wire \intermediateWiresStage3[9][43] ;
wire \intermediateWiresStage3[9][42] ;
wire \intermediateWiresStage3[9][41] ;
wire \intermediateWiresStage3[9][40] ;
wire \intermediateWiresStage3[9][39] ;
wire \intermediateWiresStage3[9][38] ;
wire \intermediateWiresStage3[9][37] ;
wire \intermediateWiresStage3[9][36] ;
wire \intermediateWiresStage3[9][35] ;
wire \intermediateWiresStage3[9][34] ;
wire \intermediateWiresStage3[9][33] ;
wire \intermediateWiresStage3[9][32] ;
wire \intermediateWiresStage3[9][31] ;
wire \intermediateWiresStage3[8][60] ;
wire \intermediateWiresStage3[8][59] ;
wire \intermediateWiresStage3[8][58] ;
wire \intermediateWiresStage3[8][57] ;
wire \intermediateWiresStage3[8][56] ;
wire \intermediateWiresStage3[8][55] ;
wire \intermediateWiresStage3[8][54] ;
wire \intermediateWiresStage3[8][53] ;
wire \intermediateWiresStage3[8][52] ;
wire \intermediateWiresStage3[8][51] ;
wire \intermediateWiresStage3[8][50] ;
wire \intermediateWiresStage3[8][49] ;
wire \intermediateWiresStage3[8][48] ;
wire \intermediateWiresStage3[8][47] ;
wire \intermediateWiresStage3[8][46] ;
wire \intermediateWiresStage3[8][45] ;
wire \intermediateWiresStage3[8][44] ;
wire \intermediateWiresStage3[8][43] ;
wire \intermediateWiresStage3[8][42] ;
wire \intermediateWiresStage3[8][41] ;
wire \intermediateWiresStage3[8][40] ;
wire \intermediateWiresStage3[8][39] ;
wire \intermediateWiresStage3[8][38] ;
wire \intermediateWiresStage3[8][37] ;
wire \intermediateWiresStage3[8][36] ;
wire \intermediateWiresStage3[8][35] ;
wire \intermediateWiresStage3[8][34] ;
wire \intermediateWiresStage3[8][33] ;
wire \intermediateWiresStage3[8][32] ;
wire \intermediateWiresStage3[8][31] ;
wire \intermediateWiresStage3[8][30] ;
wire \intermediateWiresStage3[7][57] ;
wire \intermediateWiresStage3[7][56] ;
wire \intermediateWiresStage3[7][55] ;
wire \intermediateWiresStage3[7][54] ;
wire \intermediateWiresStage3[7][53] ;
wire \intermediateWiresStage3[7][52] ;
wire \intermediateWiresStage3[7][51] ;
wire \intermediateWiresStage3[7][50] ;
wire \intermediateWiresStage3[7][49] ;
wire \intermediateWiresStage3[7][48] ;
wire \intermediateWiresStage3[7][47] ;
wire \intermediateWiresStage3[7][46] ;
wire \intermediateWiresStage3[7][45] ;
wire \intermediateWiresStage3[7][44] ;
wire \intermediateWiresStage3[7][43] ;
wire \intermediateWiresStage3[7][42] ;
wire \intermediateWiresStage3[7][41] ;
wire \intermediateWiresStage3[7][40] ;
wire \intermediateWiresStage3[7][39] ;
wire \intermediateWiresStage3[7][38] ;
wire \intermediateWiresStage3[7][37] ;
wire \intermediateWiresStage3[7][36] ;
wire \intermediateWiresStage3[7][35] ;
wire \intermediateWiresStage3[7][34] ;
wire \intermediateWiresStage3[7][33] ;
wire \intermediateWiresStage3[7][32] ;
wire \intermediateWiresStage3[7][31] ;
wire \intermediateWiresStage3[7][30] ;
wire \intermediateWiresStage3[7][29] ;
wire \intermediateWiresStage3[7][28] ;
wire \intermediateWiresStage3[7][27] ;
wire \intermediateWiresStage3[7][26] ;
wire \intermediateWiresStage3[7][25] ;
wire \intermediateWiresStage3[7][24] ;
wire \intermediateWiresStage3[6][56] ;
wire \intermediateWiresStage3[6][55] ;
wire \intermediateWiresStage3[6][54] ;
wire \intermediateWiresStage3[6][53] ;
wire \intermediateWiresStage3[6][52] ;
wire \intermediateWiresStage3[6][51] ;
wire \intermediateWiresStage3[6][50] ;
wire \intermediateWiresStage3[6][49] ;
wire \intermediateWiresStage3[6][48] ;
wire \intermediateWiresStage3[6][47] ;
wire \intermediateWiresStage3[6][46] ;
wire \intermediateWiresStage3[6][45] ;
wire \intermediateWiresStage3[6][44] ;
wire \intermediateWiresStage3[6][43] ;
wire \intermediateWiresStage3[6][42] ;
wire \intermediateWiresStage3[6][41] ;
wire \intermediateWiresStage3[6][40] ;
wire \intermediateWiresStage3[6][39] ;
wire \intermediateWiresStage3[6][38] ;
wire \intermediateWiresStage3[6][37] ;
wire \intermediateWiresStage3[6][36] ;
wire \intermediateWiresStage3[6][35] ;
wire \intermediateWiresStage3[6][34] ;
wire \intermediateWiresStage3[6][33] ;
wire \intermediateWiresStage3[6][32] ;
wire \intermediateWiresStage3[6][31] ;
wire \intermediateWiresStage3[6][30] ;
wire \intermediateWiresStage3[6][29] ;
wire \intermediateWiresStage3[6][28] ;
wire \intermediateWiresStage3[6][27] ;
wire \intermediateWiresStage3[6][26] ;
wire \intermediateWiresStage3[6][25] ;
wire \intermediateWiresStage3[6][24] ;
wire \intermediateWiresStage3[6][23] ;
wire \intermediateWiresStage3[5][49] ;
wire \intermediateWiresStage3[5][48] ;
wire \intermediateWiresStage3[5][47] ;
wire \intermediateWiresStage3[5][46] ;
wire \intermediateWiresStage3[5][45] ;
wire \intermediateWiresStage3[5][44] ;
wire \intermediateWiresStage3[5][43] ;
wire \intermediateWiresStage3[5][42] ;
wire \intermediateWiresStage3[5][41] ;
wire \intermediateWiresStage3[5][40] ;
wire \intermediateWiresStage3[5][39] ;
wire \intermediateWiresStage3[5][38] ;
wire \intermediateWiresStage3[5][37] ;
wire \intermediateWiresStage3[5][36] ;
wire \intermediateWiresStage3[5][35] ;
wire \intermediateWiresStage3[5][34] ;
wire \intermediateWiresStage3[5][33] ;
wire \intermediateWiresStage3[5][32] ;
wire \intermediateWiresStage3[5][31] ;
wire \intermediateWiresStage3[5][30] ;
wire \intermediateWiresStage3[5][29] ;
wire \intermediateWiresStage3[5][28] ;
wire \intermediateWiresStage3[5][27] ;
wire \intermediateWiresStage3[5][26] ;
wire \intermediateWiresStage3[5][25] ;
wire \intermediateWiresStage3[5][24] ;
wire \intermediateWiresStage3[5][23] ;
wire \intermediateWiresStage3[5][22] ;
wire \intermediateWiresStage3[5][21] ;
wire \intermediateWiresStage3[5][20] ;
wire \intermediateWiresStage3[5][19] ;
wire \intermediateWiresStage3[5][18] ;
wire \intermediateWiresStage3[5][17] ;
wire \intermediateWiresStage3[4][48] ;
wire \intermediateWiresStage3[4][47] ;
wire \intermediateWiresStage3[4][46] ;
wire \intermediateWiresStage3[4][45] ;
wire \intermediateWiresStage3[4][44] ;
wire \intermediateWiresStage3[4][43] ;
wire \intermediateWiresStage3[4][42] ;
wire \intermediateWiresStage3[4][41] ;
wire \intermediateWiresStage3[4][40] ;
wire \intermediateWiresStage3[4][39] ;
wire \intermediateWiresStage3[4][38] ;
wire \intermediateWiresStage3[4][37] ;
wire \intermediateWiresStage3[4][36] ;
wire \intermediateWiresStage3[4][35] ;
wire \intermediateWiresStage3[4][34] ;
wire \intermediateWiresStage3[4][33] ;
wire \intermediateWiresStage3[4][32] ;
wire \intermediateWiresStage3[4][31] ;
wire \intermediateWiresStage3[4][30] ;
wire \intermediateWiresStage3[4][29] ;
wire \intermediateWiresStage3[4][28] ;
wire \intermediateWiresStage3[4][27] ;
wire \intermediateWiresStage3[4][26] ;
wire \intermediateWiresStage3[4][25] ;
wire \intermediateWiresStage3[4][24] ;
wire \intermediateWiresStage3[4][23] ;
wire \intermediateWiresStage3[4][22] ;
wire \intermediateWiresStage3[4][21] ;
wire \intermediateWiresStage3[4][20] ;
wire \intermediateWiresStage3[4][19] ;
wire \intermediateWiresStage3[4][18] ;
wire \intermediateWiresStage3[4][17] ;
wire \intermediateWiresStage3[4][16] ;
wire \intermediateWiresStage3[3][43] ;
wire \intermediateWiresStage3[3][42] ;
wire \intermediateWiresStage3[3][41] ;
wire \intermediateWiresStage3[3][40] ;
wire \intermediateWiresStage3[3][39] ;
wire \intermediateWiresStage3[3][38] ;
wire \intermediateWiresStage3[3][37] ;
wire \intermediateWiresStage3[3][36] ;
wire \intermediateWiresStage3[3][35] ;
wire \intermediateWiresStage3[3][34] ;
wire \intermediateWiresStage3[3][33] ;
wire \intermediateWiresStage3[3][32] ;
wire \intermediateWiresStage3[3][31] ;
wire \intermediateWiresStage3[3][30] ;
wire \intermediateWiresStage3[3][29] ;
wire \intermediateWiresStage3[3][28] ;
wire \intermediateWiresStage3[3][27] ;
wire \intermediateWiresStage3[3][26] ;
wire \intermediateWiresStage3[3][25] ;
wire \intermediateWiresStage3[3][24] ;
wire \intermediateWiresStage3[3][23] ;
wire \intermediateWiresStage3[3][22] ;
wire \intermediateWiresStage3[3][21] ;
wire \intermediateWiresStage3[3][20] ;
wire \intermediateWiresStage3[3][19] ;
wire \intermediateWiresStage3[3][18] ;
wire \intermediateWiresStage3[3][17] ;
wire \intermediateWiresStage3[3][16] ;
wire \intermediateWiresStage3[3][15] ;
wire \intermediateWiresStage3[3][14] ;
wire \intermediateWiresStage3[3][13] ;
wire \intermediateWiresStage3[3][12] ;
wire \intermediateWiresStage3[3][11] ;
wire \intermediateWiresStage3[3][10] ;
wire \intermediateWiresStage3[2][42] ;
wire \intermediateWiresStage3[2][41] ;
wire \intermediateWiresStage3[2][40] ;
wire \intermediateWiresStage3[2][39] ;
wire \intermediateWiresStage3[2][38] ;
wire \intermediateWiresStage3[2][37] ;
wire \intermediateWiresStage3[2][36] ;
wire \intermediateWiresStage3[2][35] ;
wire \intermediateWiresStage3[2][34] ;
wire \intermediateWiresStage3[2][33] ;
wire \intermediateWiresStage3[2][32] ;
wire \intermediateWiresStage3[2][31] ;
wire \intermediateWiresStage3[2][30] ;
wire \intermediateWiresStage3[2][29] ;
wire \intermediateWiresStage3[2][28] ;
wire \intermediateWiresStage3[2][27] ;
wire \intermediateWiresStage3[2][26] ;
wire \intermediateWiresStage3[2][25] ;
wire \intermediateWiresStage3[2][24] ;
wire \intermediateWiresStage3[2][23] ;
wire \intermediateWiresStage3[2][22] ;
wire \intermediateWiresStage3[2][21] ;
wire \intermediateWiresStage3[2][20] ;
wire \intermediateWiresStage3[2][19] ;
wire \intermediateWiresStage3[2][18] ;
wire \intermediateWiresStage3[2][17] ;
wire \intermediateWiresStage3[2][16] ;
wire \intermediateWiresStage3[2][15] ;
wire \intermediateWiresStage3[2][14] ;
wire \intermediateWiresStage3[2][13] ;
wire \intermediateWiresStage3[2][12] ;
wire \intermediateWiresStage3[2][11] ;
wire \intermediateWiresStage3[2][10] ;
wire \intermediateWiresStage3[2][9] ;
wire \intermediateWiresStage3[1][36] ;
wire \intermediateWiresStage3[1][35] ;
wire \intermediateWiresStage3[1][34] ;
wire \intermediateWiresStage3[1][33] ;
wire \intermediateWiresStage3[1][32] ;
wire \intermediateWiresStage3[1][31] ;
wire \intermediateWiresStage3[1][30] ;
wire \intermediateWiresStage3[1][29] ;
wire \intermediateWiresStage3[1][28] ;
wire \intermediateWiresStage3[1][27] ;
wire \intermediateWiresStage3[1][26] ;
wire \intermediateWiresStage3[1][25] ;
wire \intermediateWiresStage3[1][24] ;
wire \intermediateWiresStage3[1][23] ;
wire \intermediateWiresStage3[1][22] ;
wire \intermediateWiresStage3[1][21] ;
wire \intermediateWiresStage3[1][20] ;
wire \intermediateWiresStage3[1][19] ;
wire \intermediateWiresStage3[1][18] ;
wire \intermediateWiresStage3[1][17] ;
wire \intermediateWiresStage3[1][16] ;
wire \intermediateWiresStage3[1][15] ;
wire \intermediateWiresStage3[1][14] ;
wire \intermediateWiresStage3[1][13] ;
wire \intermediateWiresStage3[1][12] ;
wire \intermediateWiresStage3[1][11] ;
wire \intermediateWiresStage3[1][10] ;
wire \intermediateWiresStage3[1][9] ;
wire \intermediateWiresStage3[1][8] ;
wire \intermediateWiresStage3[1][7] ;
wire \intermediateWiresStage3[1][6] ;
wire \intermediateWiresStage3[1][5] ;
wire \intermediateWiresStage3[1][4] ;
wire \intermediateWiresStage3[0][35] ;
wire \intermediateWiresStage3[0][34] ;
wire \intermediateWiresStage3[0][33] ;
wire \intermediateWiresStage3[0][32] ;
wire \intermediateWiresStage3[0][31] ;
wire \intermediateWiresStage3[0][30] ;
wire \intermediateWiresStage3[0][29] ;
wire \intermediateWiresStage3[0][28] ;
wire \intermediateWiresStage3[0][27] ;
wire \intermediateWiresStage3[0][26] ;
wire \intermediateWiresStage3[0][25] ;
wire \intermediateWiresStage3[0][24] ;
wire \intermediateWiresStage3[0][23] ;
wire \intermediateWiresStage3[0][22] ;
wire \intermediateWiresStage3[0][21] ;
wire \intermediateWiresStage3[0][20] ;
wire \intermediateWiresStage3[0][19] ;
wire \intermediateWiresStage3[0][18] ;
wire \intermediateWiresStage3[0][17] ;
wire \intermediateWiresStage3[0][16] ;
wire \intermediateWiresStage3[0][15] ;
wire \intermediateWiresStage3[0][14] ;
wire \intermediateWiresStage3[0][13] ;
wire \intermediateWiresStage3[0][12] ;
wire \intermediateWiresStage3[0][11] ;
wire \intermediateWiresStage3[0][10] ;
wire \intermediateWiresStage3[0][9] ;
wire \intermediateWiresStage3[0][8] ;
wire \intermediateWiresStage3[0][7] ;
wire \intermediateWiresStage3[0][6] ;
wire \intermediateWiresStage3[0][5] ;
wire \intermediateWiresStage3[0][4] ;
wire \intermediateWiresStage4[5][58] ;
wire \intermediateWiresStage4[5][57] ;
wire \intermediateWiresStage4[5][56] ;
wire \intermediateWiresStage4[5][55] ;
wire \intermediateWiresStage4[5][54] ;
wire \intermediateWiresStage4[5][53] ;
wire \intermediateWiresStage4[5][52] ;
wire \intermediateWiresStage4[5][51] ;
wire \intermediateWiresStage4[5][50] ;
wire \intermediateWiresStage4[5][49] ;
wire \intermediateWiresStage4[5][48] ;
wire \intermediateWiresStage4[5][47] ;
wire \intermediateWiresStage4[5][46] ;
wire \intermediateWiresStage4[5][45] ;
wire \intermediateWiresStage4[5][44] ;
wire \intermediateWiresStage4[5][43] ;
wire \intermediateWiresStage4[5][42] ;
wire \intermediateWiresStage4[5][41] ;
wire \intermediateWiresStage4[5][40] ;
wire \intermediateWiresStage4[5][39] ;
wire \intermediateWiresStage4[5][38] ;
wire \intermediateWiresStage4[5][37] ;
wire \intermediateWiresStage4[5][36] ;
wire \intermediateWiresStage4[5][35] ;
wire \intermediateWiresStage4[5][34] ;
wire \intermediateWiresStage4[5][33] ;
wire \intermediateWiresStage4[5][32] ;
wire \intermediateWiresStage4[5][31] ;
wire \intermediateWiresStage4[5][30] ;
wire \intermediateWiresStage4[5][29] ;
wire \intermediateWiresStage4[5][28] ;
wire \intermediateWiresStage4[5][27] ;
wire \intermediateWiresStage4[5][26] ;
wire \intermediateWiresStage4[5][25] ;
wire \intermediateWiresStage4[4][57] ;
wire \intermediateWiresStage4[4][56] ;
wire \intermediateWiresStage4[4][55] ;
wire \intermediateWiresStage4[4][54] ;
wire \intermediateWiresStage4[4][53] ;
wire \intermediateWiresStage4[4][52] ;
wire \intermediateWiresStage4[4][51] ;
wire \intermediateWiresStage4[4][50] ;
wire \intermediateWiresStage4[4][49] ;
wire \intermediateWiresStage4[4][48] ;
wire \intermediateWiresStage4[4][47] ;
wire \intermediateWiresStage4[4][46] ;
wire \intermediateWiresStage4[4][45] ;
wire \intermediateWiresStage4[4][44] ;
wire \intermediateWiresStage4[4][43] ;
wire \intermediateWiresStage4[4][42] ;
wire \intermediateWiresStage4[4][41] ;
wire \intermediateWiresStage4[4][40] ;
wire \intermediateWiresStage4[4][39] ;
wire \intermediateWiresStage4[4][38] ;
wire \intermediateWiresStage4[4][37] ;
wire \intermediateWiresStage4[4][36] ;
wire \intermediateWiresStage4[4][35] ;
wire \intermediateWiresStage4[4][34] ;
wire \intermediateWiresStage4[4][33] ;
wire \intermediateWiresStage4[4][32] ;
wire \intermediateWiresStage4[4][31] ;
wire \intermediateWiresStage4[4][30] ;
wire \intermediateWiresStage4[4][29] ;
wire \intermediateWiresStage4[4][28] ;
wire \intermediateWiresStage4[4][27] ;
wire \intermediateWiresStage4[4][26] ;
wire \intermediateWiresStage4[4][25] ;
wire \intermediateWiresStage4[4][24] ;
wire \intermediateWiresStage4[3][50] ;
wire \intermediateWiresStage4[3][49] ;
wire \intermediateWiresStage4[3][48] ;
wire \intermediateWiresStage4[3][47] ;
wire \intermediateWiresStage4[3][46] ;
wire \intermediateWiresStage4[3][45] ;
wire \intermediateWiresStage4[3][44] ;
wire \intermediateWiresStage4[3][43] ;
wire \intermediateWiresStage4[3][42] ;
wire \intermediateWiresStage4[3][41] ;
wire \intermediateWiresStage4[3][40] ;
wire \intermediateWiresStage4[3][39] ;
wire \intermediateWiresStage4[3][38] ;
wire \intermediateWiresStage4[3][37] ;
wire \intermediateWiresStage4[3][36] ;
wire \intermediateWiresStage4[3][35] ;
wire \intermediateWiresStage4[3][34] ;
wire \intermediateWiresStage4[3][33] ;
wire \intermediateWiresStage4[3][32] ;
wire \intermediateWiresStage4[3][31] ;
wire \intermediateWiresStage4[3][30] ;
wire \intermediateWiresStage4[3][29] ;
wire \intermediateWiresStage4[3][28] ;
wire \intermediateWiresStage4[3][27] ;
wire \intermediateWiresStage4[3][26] ;
wire \intermediateWiresStage4[3][25] ;
wire \intermediateWiresStage4[3][24] ;
wire \intermediateWiresStage4[3][23] ;
wire \intermediateWiresStage4[3][22] ;
wire \intermediateWiresStage4[3][21] ;
wire \intermediateWiresStage4[3][20] ;
wire \intermediateWiresStage4[3][19] ;
wire \intermediateWiresStage4[3][18] ;
wire \intermediateWiresStage4[3][17] ;
wire \intermediateWiresStage4[3][16] ;
wire \intermediateWiresStage4[3][15] ;
wire \intermediateWiresStage4[2][49] ;
wire \intermediateWiresStage4[2][48] ;
wire \intermediateWiresStage4[2][47] ;
wire \intermediateWiresStage4[2][46] ;
wire \intermediateWiresStage4[2][45] ;
wire \intermediateWiresStage4[2][44] ;
wire \intermediateWiresStage4[2][43] ;
wire \intermediateWiresStage4[2][42] ;
wire \intermediateWiresStage4[2][41] ;
wire \intermediateWiresStage4[2][40] ;
wire \intermediateWiresStage4[2][39] ;
wire \intermediateWiresStage4[2][38] ;
wire \intermediateWiresStage4[2][37] ;
wire \intermediateWiresStage4[2][36] ;
wire \intermediateWiresStage4[2][35] ;
wire \intermediateWiresStage4[2][34] ;
wire \intermediateWiresStage4[2][33] ;
wire \intermediateWiresStage4[2][32] ;
wire \intermediateWiresStage4[2][31] ;
wire \intermediateWiresStage4[2][30] ;
wire \intermediateWiresStage4[2][29] ;
wire \intermediateWiresStage4[2][28] ;
wire \intermediateWiresStage4[2][27] ;
wire \intermediateWiresStage4[2][26] ;
wire \intermediateWiresStage4[2][25] ;
wire \intermediateWiresStage4[2][24] ;
wire \intermediateWiresStage4[2][23] ;
wire \intermediateWiresStage4[2][22] ;
wire \intermediateWiresStage4[2][21] ;
wire \intermediateWiresStage4[2][20] ;
wire \intermediateWiresStage4[2][19] ;
wire \intermediateWiresStage4[2][18] ;
wire \intermediateWiresStage4[2][17] ;
wire \intermediateWiresStage4[2][16] ;
wire \intermediateWiresStage4[2][15] ;
wire \intermediateWiresStage4[2][14] ;
wire \intermediateWiresStage4[1][39] ;
wire \intermediateWiresStage4[1][38] ;
wire \intermediateWiresStage4[1][37] ;
wire \intermediateWiresStage4[1][36] ;
wire \intermediateWiresStage4[1][35] ;
wire \intermediateWiresStage4[1][34] ;
wire \intermediateWiresStage4[1][33] ;
wire \intermediateWiresStage4[1][32] ;
wire \intermediateWiresStage4[1][31] ;
wire \intermediateWiresStage4[1][30] ;
wire \intermediateWiresStage4[1][29] ;
wire \intermediateWiresStage4[1][28] ;
wire \intermediateWiresStage4[1][27] ;
wire \intermediateWiresStage4[1][26] ;
wire \intermediateWiresStage4[1][25] ;
wire \intermediateWiresStage4[1][24] ;
wire \intermediateWiresStage4[1][23] ;
wire \intermediateWiresStage4[1][22] ;
wire \intermediateWiresStage4[1][21] ;
wire \intermediateWiresStage4[1][20] ;
wire \intermediateWiresStage4[1][19] ;
wire \intermediateWiresStage4[1][18] ;
wire \intermediateWiresStage4[1][17] ;
wire \intermediateWiresStage4[1][16] ;
wire \intermediateWiresStage4[1][15] ;
wire \intermediateWiresStage4[1][14] ;
wire \intermediateWiresStage4[1][13] ;
wire \intermediateWiresStage4[1][12] ;
wire \intermediateWiresStage4[1][11] ;
wire \intermediateWiresStage4[1][10] ;
wire \intermediateWiresStage4[1][9] ;
wire \intermediateWiresStage4[1][8] ;
wire \intermediateWiresStage4[1][7] ;
wire \intermediateWiresStage4[1][6] ;
wire \intermediateWiresStage4[1][5] ;
wire \intermediateWiresStage4[0][38] ;
wire \intermediateWiresStage4[0][37] ;
wire \intermediateWiresStage4[0][36] ;
wire \intermediateWiresStage4[0][35] ;
wire \intermediateWiresStage4[0][34] ;
wire \intermediateWiresStage4[0][33] ;
wire \intermediateWiresStage4[0][32] ;
wire \intermediateWiresStage4[0][31] ;
wire \intermediateWiresStage4[0][30] ;
wire \intermediateWiresStage4[0][29] ;
wire \intermediateWiresStage4[0][28] ;
wire \intermediateWiresStage4[0][27] ;
wire \intermediateWiresStage4[0][26] ;
wire \intermediateWiresStage4[0][25] ;
wire \intermediateWiresStage4[0][24] ;
wire \intermediateWiresStage4[0][23] ;
wire \intermediateWiresStage4[0][22] ;
wire \intermediateWiresStage4[0][21] ;
wire \intermediateWiresStage4[0][20] ;
wire \intermediateWiresStage4[0][19] ;
wire \intermediateWiresStage4[0][18] ;
wire \intermediateWiresStage4[0][17] ;
wire \intermediateWiresStage4[0][16] ;
wire \intermediateWiresStage4[0][15] ;
wire \intermediateWiresStage4[0][14] ;
wire \intermediateWiresStage4[0][13] ;
wire \intermediateWiresStage4[0][12] ;
wire \intermediateWiresStage4[0][11] ;
wire \intermediateWiresStage4[0][10] ;
wire \intermediateWiresStage4[0][9] ;
wire \intermediateWiresStage4[0][8] ;
wire \intermediateWiresStage4[0][7] ;
wire \intermediateWiresStage4[0][6] ;
wire \intermediateWiresStage4[0][5] ;
wire \intermediateWiresStage5[3][59] ;
wire \intermediateWiresStage5[3][58] ;
wire \intermediateWiresStage5[3][57] ;
wire \intermediateWiresStage5[3][56] ;
wire \intermediateWiresStage5[3][55] ;
wire \intermediateWiresStage5[3][54] ;
wire \intermediateWiresStage5[3][53] ;
wire \intermediateWiresStage5[3][52] ;
wire \intermediateWiresStage5[3][51] ;
wire \intermediateWiresStage5[3][50] ;
wire \intermediateWiresStage5[3][49] ;
wire \intermediateWiresStage5[3][48] ;
wire \intermediateWiresStage5[3][47] ;
wire \intermediateWiresStage5[3][46] ;
wire \intermediateWiresStage5[3][45] ;
wire \intermediateWiresStage5[3][44] ;
wire \intermediateWiresStage5[3][43] ;
wire \intermediateWiresStage5[3][42] ;
wire \intermediateWiresStage5[3][41] ;
wire \intermediateWiresStage5[3][40] ;
wire \intermediateWiresStage5[3][39] ;
wire \intermediateWiresStage5[3][38] ;
wire \intermediateWiresStage5[3][37] ;
wire \intermediateWiresStage5[3][36] ;
wire \intermediateWiresStage5[3][35] ;
wire \intermediateWiresStage5[3][34] ;
wire \intermediateWiresStage5[3][33] ;
wire \intermediateWiresStage5[3][32] ;
wire \intermediateWiresStage5[3][31] ;
wire \intermediateWiresStage5[3][30] ;
wire \intermediateWiresStage5[3][29] ;
wire \intermediateWiresStage5[3][28] ;
wire \intermediateWiresStage5[3][27] ;
wire \intermediateWiresStage5[3][26] ;
wire \intermediateWiresStage5[3][25] ;
wire \intermediateWiresStage5[3][24] ;
wire \intermediateWiresStage5[3][23] ;
wire \intermediateWiresStage5[3][22] ;
wire \intermediateWiresStage5[2][58] ;
wire \intermediateWiresStage5[2][57] ;
wire \intermediateWiresStage5[2][56] ;
wire \intermediateWiresStage5[2][55] ;
wire \intermediateWiresStage5[2][54] ;
wire \intermediateWiresStage5[2][53] ;
wire \intermediateWiresStage5[2][52] ;
wire \intermediateWiresStage5[2][51] ;
wire \intermediateWiresStage5[2][50] ;
wire \intermediateWiresStage5[2][49] ;
wire \intermediateWiresStage5[2][48] ;
wire \intermediateWiresStage5[2][47] ;
wire \intermediateWiresStage5[2][46] ;
wire \intermediateWiresStage5[2][45] ;
wire \intermediateWiresStage5[2][44] ;
wire \intermediateWiresStage5[2][43] ;
wire \intermediateWiresStage5[2][42] ;
wire \intermediateWiresStage5[2][41] ;
wire \intermediateWiresStage5[2][40] ;
wire \intermediateWiresStage5[2][39] ;
wire \intermediateWiresStage5[2][38] ;
wire \intermediateWiresStage5[2][37] ;
wire \intermediateWiresStage5[2][36] ;
wire \intermediateWiresStage5[2][35] ;
wire \intermediateWiresStage5[2][34] ;
wire \intermediateWiresStage5[2][33] ;
wire \intermediateWiresStage5[2][32] ;
wire \intermediateWiresStage5[2][31] ;
wire \intermediateWiresStage5[2][30] ;
wire \intermediateWiresStage5[2][29] ;
wire \intermediateWiresStage5[2][28] ;
wire \intermediateWiresStage5[2][27] ;
wire \intermediateWiresStage5[2][26] ;
wire \intermediateWiresStage5[2][25] ;
wire \intermediateWiresStage5[2][24] ;
wire \intermediateWiresStage5[2][23] ;
wire \intermediateWiresStage5[2][22] ;
wire \intermediateWiresStage5[2][21] ;
wire \intermediateWiresStage5[1][45] ;
wire \intermediateWiresStage5[1][44] ;
wire \intermediateWiresStage5[1][43] ;
wire \intermediateWiresStage5[1][42] ;
wire \intermediateWiresStage5[1][41] ;
wire \intermediateWiresStage5[1][40] ;
wire \intermediateWiresStage5[1][39] ;
wire \intermediateWiresStage5[1][38] ;
wire \intermediateWiresStage5[1][37] ;
wire \intermediateWiresStage5[1][36] ;
wire \intermediateWiresStage5[1][35] ;
wire \intermediateWiresStage5[1][34] ;
wire \intermediateWiresStage5[1][33] ;
wire \intermediateWiresStage5[1][32] ;
wire \intermediateWiresStage5[1][31] ;
wire \intermediateWiresStage5[1][30] ;
wire \intermediateWiresStage5[1][29] ;
wire \intermediateWiresStage5[1][28] ;
wire \intermediateWiresStage5[1][27] ;
wire \intermediateWiresStage5[1][26] ;
wire \intermediateWiresStage5[1][25] ;
wire \intermediateWiresStage5[1][24] ;
wire \intermediateWiresStage5[1][23] ;
wire \intermediateWiresStage5[1][22] ;
wire \intermediateWiresStage5[1][21] ;
wire \intermediateWiresStage5[1][20] ;
wire \intermediateWiresStage5[1][19] ;
wire \intermediateWiresStage5[1][18] ;
wire \intermediateWiresStage5[1][17] ;
wire \intermediateWiresStage5[1][16] ;
wire \intermediateWiresStage5[1][15] ;
wire \intermediateWiresStage5[1][14] ;
wire \intermediateWiresStage5[1][13] ;
wire \intermediateWiresStage5[1][12] ;
wire \intermediateWiresStage5[1][11] ;
wire \intermediateWiresStage5[1][10] ;
wire \intermediateWiresStage5[1][9] ;
wire \intermediateWiresStage5[1][8] ;
wire \intermediateWiresStage5[1][7] ;
wire \intermediateWiresStage5[1][6] ;
wire \intermediateWiresStage5[0][44] ;
wire \intermediateWiresStage5[0][43] ;
wire \intermediateWiresStage5[0][42] ;
wire \intermediateWiresStage5[0][41] ;
wire \intermediateWiresStage5[0][40] ;
wire \intermediateWiresStage5[0][39] ;
wire \intermediateWiresStage5[0][38] ;
wire \intermediateWiresStage5[0][37] ;
wire \intermediateWiresStage5[0][36] ;
wire \intermediateWiresStage5[0][35] ;
wire \intermediateWiresStage5[0][34] ;
wire \intermediateWiresStage5[0][33] ;
wire \intermediateWiresStage5[0][32] ;
wire \intermediateWiresStage5[0][31] ;
wire \intermediateWiresStage5[0][30] ;
wire \intermediateWiresStage5[0][29] ;
wire \intermediateWiresStage5[0][28] ;
wire \intermediateWiresStage5[0][27] ;
wire \intermediateWiresStage5[0][26] ;
wire \intermediateWiresStage5[0][25] ;
wire \intermediateWiresStage5[0][24] ;
wire \intermediateWiresStage5[0][23] ;
wire \intermediateWiresStage5[0][22] ;
wire \intermediateWiresStage5[0][21] ;
wire \intermediateWiresStage5[0][20] ;
wire \intermediateWiresStage5[0][19] ;
wire \intermediateWiresStage5[0][18] ;
wire \intermediateWiresStage5[0][17] ;
wire \intermediateWiresStage5[0][16] ;
wire \intermediateWiresStage5[0][15] ;
wire \intermediateWiresStage5[0][14] ;
wire \intermediateWiresStage5[0][13] ;
wire \intermediateWiresStage5[0][12] ;
wire \intermediateWiresStage5[0][11] ;
wire \intermediateWiresStage5[0][10] ;
wire \intermediateWiresStage5[0][9] ;
wire \intermediateWiresStage5[0][8] ;
wire \intermediateWiresStage5[0][7] ;
wire \intermediateWiresStage5[0][6] ;
wire \intermediateWiresStage6[1][54] ;
wire \intermediateWiresStage6[1][53] ;
wire \intermediateWiresStage6[1][52] ;
wire \intermediateWiresStage6[1][51] ;
wire \intermediateWiresStage6[1][50] ;
wire \intermediateWiresStage6[1][49] ;
wire \intermediateWiresStage6[1][48] ;
wire \intermediateWiresStage6[1][47] ;
wire \intermediateWiresStage6[1][46] ;
wire \intermediateWiresStage6[1][45] ;
wire \intermediateWiresStage6[1][44] ;
wire \intermediateWiresStage6[1][43] ;
wire \intermediateWiresStage6[1][42] ;
wire \intermediateWiresStage6[1][41] ;
wire \intermediateWiresStage6[1][40] ;
wire \intermediateWiresStage6[1][39] ;
wire \intermediateWiresStage6[1][38] ;
wire \intermediateWiresStage6[1][37] ;
wire \intermediateWiresStage6[1][36] ;
wire \intermediateWiresStage6[1][35] ;
wire \intermediateWiresStage6[1][34] ;
wire \intermediateWiresStage6[1][33] ;
wire \intermediateWiresStage6[1][32] ;
wire \intermediateWiresStage6[1][31] ;
wire \intermediateWiresStage6[1][30] ;
wire \intermediateWiresStage6[1][29] ;
wire \intermediateWiresStage6[1][28] ;
wire \intermediateWiresStage6[1][27] ;
wire \intermediateWiresStage6[1][26] ;
wire \intermediateWiresStage6[1][25] ;
wire \intermediateWiresStage6[1][24] ;
wire \intermediateWiresStage6[1][23] ;
wire \intermediateWiresStage6[1][22] ;
wire \intermediateWiresStage6[1][21] ;
wire \intermediateWiresStage6[1][20] ;
wire \intermediateWiresStage6[1][19] ;
wire \intermediateWiresStage6[1][18] ;
wire \intermediateWiresStage6[1][17] ;
wire \intermediateWiresStage6[1][16] ;
wire \intermediateWiresStage6[1][15] ;
wire \intermediateWiresStage6[1][14] ;
wire \intermediateWiresStage6[1][13] ;
wire \intermediateWiresStage6[1][12] ;
wire \intermediateWiresStage6[1][11] ;
wire \intermediateWiresStage6[1][10] ;
wire \intermediateWiresStage6[1][9] ;
wire \intermediateWiresStage6[1][8] ;
wire \intermediateWiresStage6[1][7] ;
wire \intermediateWiresStage6[0][53] ;
wire \intermediateWiresStage6[0][52] ;
wire \intermediateWiresStage6[0][51] ;
wire \intermediateWiresStage6[0][50] ;
wire \intermediateWiresStage6[0][49] ;
wire \intermediateWiresStage6[0][48] ;
wire \intermediateWiresStage6[0][47] ;
wire \intermediateWiresStage6[0][46] ;
wire \intermediateWiresStage6[0][45] ;
wire \intermediateWiresStage6[0][44] ;
wire \intermediateWiresStage6[0][43] ;
wire \intermediateWiresStage6[0][42] ;
wire \intermediateWiresStage6[0][41] ;
wire \intermediateWiresStage6[0][40] ;
wire \intermediateWiresStage6[0][39] ;
wire \intermediateWiresStage6[0][38] ;
wire \intermediateWiresStage6[0][37] ;
wire \intermediateWiresStage6[0][36] ;
wire \intermediateWiresStage6[0][35] ;
wire \intermediateWiresStage6[0][34] ;
wire \intermediateWiresStage6[0][33] ;
wire \intermediateWiresStage6[0][32] ;
wire \intermediateWiresStage6[0][31] ;
wire \intermediateWiresStage6[0][30] ;
wire \intermediateWiresStage6[0][29] ;
wire \intermediateWiresStage6[0][28] ;
wire \intermediateWiresStage6[0][27] ;
wire \intermediateWiresStage6[0][26] ;
wire \intermediateWiresStage6[0][25] ;
wire \intermediateWiresStage6[0][24] ;
wire \intermediateWiresStage6[0][23] ;
wire \intermediateWiresStage6[0][22] ;
wire \intermediateWiresStage6[0][21] ;
wire \intermediateWiresStage6[0][20] ;
wire \intermediateWiresStage6[0][19] ;
wire \intermediateWiresStage6[0][18] ;
wire \intermediateWiresStage6[0][17] ;
wire \intermediateWiresStage6[0][16] ;
wire \intermediateWiresStage6[0][15] ;
wire \intermediateWiresStage6[0][14] ;
wire \intermediateWiresStage6[0][13] ;
wire \intermediateWiresStage6[0][12] ;
wire \intermediateWiresStage6[0][11] ;
wire \intermediateWiresStage6[0][10] ;
wire \intermediateWiresStage6[0][9] ;
wire \intermediateWiresStage6[0][8] ;
wire \intermediateWiresStage6[0][7] ;
wire \intermediateWiresStage7[1][60] ;
wire \intermediateWiresStage7[1][59] ;
wire \intermediateWiresStage7[1][58] ;
wire \intermediateWiresStage7[1][57] ;
wire \intermediateWiresStage7[1][56] ;
wire \intermediateWiresStage7[1][55] ;
wire \intermediateWiresStage7[1][54] ;
wire \intermediateWiresStage7[1][53] ;
wire \intermediateWiresStage7[1][52] ;
wire \intermediateWiresStage7[1][51] ;
wire \intermediateWiresStage7[1][50] ;
wire \intermediateWiresStage7[1][49] ;
wire \intermediateWiresStage7[1][48] ;
wire \intermediateWiresStage7[1][47] ;
wire \intermediateWiresStage7[1][46] ;
wire \intermediateWiresStage7[1][45] ;
wire \intermediateWiresStage7[1][44] ;
wire \intermediateWiresStage7[1][43] ;
wire \intermediateWiresStage7[1][42] ;
wire \intermediateWiresStage7[1][41] ;
wire \intermediateWiresStage7[1][40] ;
wire \intermediateWiresStage7[1][39] ;
wire \intermediateWiresStage7[1][38] ;
wire \intermediateWiresStage7[1][37] ;
wire \intermediateWiresStage7[1][36] ;
wire \intermediateWiresStage7[1][35] ;
wire \intermediateWiresStage7[1][34] ;
wire \intermediateWiresStage7[1][33] ;
wire \intermediateWiresStage7[1][32] ;
wire \intermediateWiresStage7[1][31] ;
wire \intermediateWiresStage7[1][30] ;
wire \intermediateWiresStage7[1][29] ;
wire \intermediateWiresStage7[1][28] ;
wire \intermediateWiresStage7[1][27] ;
wire \intermediateWiresStage7[1][26] ;
wire \intermediateWiresStage7[1][25] ;
wire \intermediateWiresStage7[1][24] ;
wire \intermediateWiresStage7[1][23] ;
wire \intermediateWiresStage7[1][22] ;
wire \intermediateWiresStage7[1][21] ;
wire \intermediateWiresStage7[1][20] ;
wire \intermediateWiresStage7[1][19] ;
wire \intermediateWiresStage7[1][18] ;
wire \intermediateWiresStage7[1][17] ;
wire \intermediateWiresStage7[1][16] ;
wire \intermediateWiresStage7[1][15] ;
wire \intermediateWiresStage7[1][14] ;
wire \intermediateWiresStage7[1][13] ;
wire \intermediateWiresStage7[1][12] ;
wire \intermediateWiresStage7[1][11] ;
wire \intermediateWiresStage7[1][10] ;
wire \intermediateWiresStage7[1][9] ;
wire \intermediateWiresStage7[1][8] ;
wire \intermediateWiresStage7[0][59] ;
wire \intermediateWiresStage7[0][58] ;
wire \intermediateWiresStage7[0][57] ;
wire \intermediateWiresStage7[0][56] ;
wire \intermediateWiresStage7[0][55] ;
wire \intermediateWiresStage7[0][54] ;
wire \intermediateWiresStage7[0][53] ;
wire \intermediateWiresStage7[0][52] ;
wire \intermediateWiresStage7[0][51] ;
wire \intermediateWiresStage7[0][50] ;
wire \intermediateWiresStage7[0][49] ;
wire \intermediateWiresStage7[0][48] ;
wire \intermediateWiresStage7[0][47] ;
wire \intermediateWiresStage7[0][46] ;
wire \intermediateWiresStage7[0][45] ;
wire \intermediateWiresStage7[0][44] ;
wire \intermediateWiresStage7[0][43] ;
wire \intermediateWiresStage7[0][42] ;
wire \intermediateWiresStage7[0][41] ;
wire \intermediateWiresStage7[0][40] ;
wire \intermediateWiresStage7[0][39] ;
wire \intermediateWiresStage7[0][38] ;
wire \intermediateWiresStage7[0][37] ;
wire \intermediateWiresStage7[0][36] ;
wire \intermediateWiresStage7[0][35] ;
wire \intermediateWiresStage7[0][34] ;
wire \intermediateWiresStage7[0][33] ;
wire \intermediateWiresStage7[0][32] ;
wire \intermediateWiresStage7[0][31] ;
wire \intermediateWiresStage7[0][30] ;
wire \intermediateWiresStage7[0][29] ;
wire \intermediateWiresStage7[0][28] ;
wire \intermediateWiresStage7[0][27] ;
wire \intermediateWiresStage7[0][26] ;
wire \intermediateWiresStage7[0][25] ;
wire \intermediateWiresStage7[0][24] ;
wire \intermediateWiresStage7[0][23] ;
wire \intermediateWiresStage7[0][22] ;
wire \intermediateWiresStage7[0][21] ;
wire \intermediateWiresStage7[0][20] ;
wire \intermediateWiresStage7[0][19] ;
wire \intermediateWiresStage7[0][18] ;
wire \intermediateWiresStage7[0][17] ;
wire \intermediateWiresStage7[0][16] ;
wire \intermediateWiresStage7[0][15] ;
wire \intermediateWiresStage7[0][14] ;
wire \intermediateWiresStage7[0][13] ;
wire \intermediateWiresStage7[0][12] ;
wire \intermediateWiresStage7[0][11] ;
wire \intermediateWiresStage7[0][10] ;
wire \intermediateWiresStage7[0][9] ;
wire \intermediateWiresStage7[0][8] ;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire uc_28;
wire uc_29;
wire uc_30;
wire uc_31;
wire uc_32;
wire uc_33;
wire uc_34;
wire uc_35;
wire uc_36;
wire uc_37;
wire uc_38;
wire uc_39;
wire uc_40;
wire uc_41;
wire uc_42;
wire uc_43;
wire uc_44;
wire uc_45;
wire uc_46;
wire uc_47;
wire uc_48;
wire uc_49;
wire uc_50;
wire uc_51;
wire uc_52;
wire uc_53;
wire uc_54;
wire uc_55;
wire uc_56;
wire uc_57;
wire uc_58;
wire uc_59;
wire uc_60;
wire uc_61;
wire uc_62;
wire uc_63;
wire uc_64;
wire uc_65;
wire uc_66;
wire uc_67;
wire uc_68;
wire uc_69;
wire uc_70;
wire uc_71;
wire uc_72;
wire uc_73;
wire uc_74;
wire uc_75;
wire uc_76;
wire uc_77;
wire uc_78;
wire uc_79;
wire uc_80;
wire uc_81;
wire uc_82;
wire uc_83;
wire uc_84;
wire uc_85;
wire uc_86;
wire uc_87;
wire uc_88;
wire uc_89;
wire uc_90;
wire uc_91;
wire uc_92;
wire uc_93;
wire uc_94;
wire uc_95;
wire uc_96;
wire uc_97;
wire uc_98;
wire uc_99;
wire uc_100;
wire uc_101;
wire uc_102;
wire uc_103;
wire uc_104;
wire uc_105;
wire uc_106;
wire uc_107;
wire uc_108;
wire uc_109;
wire uc_110;
wire uc_111;
wire uc_112;
wire uc_113;
wire uc_114;
wire uc_115;
wire uc_116;
wire uc_117;
wire uc_118;
wire uc_119;
wire uc_120;
wire uc_121;
wire uc_122;
wire uc_123;
wire uc_124;
wire uc_125;
wire uc_126;
wire uc_127;
wire uc_128;
wire uc_129;
wire uc_130;
wire uc_131;
wire uc_132;
wire uc_133;
wire uc_134;
wire uc_135;
wire uc_136;
wire uc_137;
wire uc_138;
wire uc_139;
wire uc_140;
wire uc_141;
wire uc_142;
wire uc_143;
wire uc_144;
wire uc_145;
wire uc_146;
wire uc_147;
wire uc_148;
wire uc_149;
wire uc_150;
wire uc_151;
wire uc_152;
wire uc_153;
wire uc_154;
wire uc_155;
wire uc_156;
wire uc_157;
wire uc_158;
wire uc_159;
wire uc_160;
wire uc_161;
wire uc_162;
wire uc_163;
wire uc_164;
wire uc_165;
wire uc_166;
wire uc_167;
wire uc_168;
wire uc_169;
wire uc_170;
wire uc_171;
wire uc_172;
wire uc_173;
wire uc_174;
wire uc_175;
wire uc_176;
wire uc_177;
wire uc_178;
wire uc_179;
wire uc_180;
wire uc_181;
wire uc_182;
wire uc_183;
wire uc_184;
wire uc_185;
wire uc_186;
wire uc_187;
wire uc_188;
wire uc_189;
wire uc_190;
wire uc_191;
wire uc_192;
wire uc_193;
wire uc_194;
wire uc_195;
wire uc_196;
wire uc_197;
wire uc_198;
wire uc_199;
wire uc_200;
wire uc_201;
wire uc_202;
wire uc_203;
wire uc_204;
wire uc_205;
wire uc_206;
wire uc_207;
wire uc_208;
wire uc_209;
wire uc_210;
wire uc_211;
wire uc_212;
wire uc_213;
wire uc_214;
wire uc_215;
wire uc_216;
wire uc_217;
wire uc_218;
wire uc_219;
wire uc_220;
wire uc_221;
wire uc_222;
wire uc_223;
wire uc_224;
wire uc_225;
wire uc_226;
wire uc_227;
wire uc_228;
wire uc_229;
wire uc_230;
wire uc_231;
wire uc_232;
wire uc_233;
wire uc_234;
wire uc_235;
wire uc_236;
wire uc_237;
wire uc_238;
wire uc_239;
wire uc_240;
wire uc_241;
wire uc_242;
wire uc_243;
wire uc_244;
wire uc_245;
wire uc_246;
wire uc_247;
wire uc_248;
wire uc_249;
wire uc_250;
wire uc_251;
wire uc_252;
wire uc_253;
wire uc_254;
wire uc_255;
wire uc_256;
wire uc_257;
wire uc_258;
wire uc_259;
wire uc_260;
wire uc_261;
wire uc_262;
wire uc_263;
wire uc_264;
wire uc_265;
wire uc_266;
wire uc_267;
wire uc_268;
wire uc_269;
wire uc_270;
wire uc_271;
wire uc_272;
wire uc_273;
wire uc_274;
wire uc_275;
wire uc_276;
wire uc_277;
wire uc_278;
wire uc_279;
wire uc_280;
wire uc_281;
wire uc_282;
wire uc_283;
wire uc_284;
wire uc_285;
wire uc_286;
wire uc_287;
wire uc_288;
wire uc_289;
wire uc_290;
wire uc_291;
wire uc_292;
wire uc_293;
wire uc_294;
wire uc_295;
wire uc_296;
wire uc_297;
wire uc_298;
wire uc_299;
wire uc_300;
wire uc_301;
wire uc_302;
wire uc_303;
wire uc_304;
wire uc_305;
wire uc_306;
wire uc_307;
wire uc_308;
wire uc_309;
wire uc_310;
wire uc_311;
wire uc_312;
wire uc_313;
wire uc_314;
wire uc_315;
wire uc_316;
wire uc_317;
wire uc_318;
wire uc_319;
wire uc_320;
wire uc_321;
wire uc_322;
wire uc_323;
wire uc_324;
wire uc_325;
wire uc_326;
wire uc_327;
wire uc_328;
wire uc_329;
wire uc_330;
wire uc_331;
wire uc_332;
wire uc_333;
wire uc_334;
wire uc_335;
wire uc_336;
wire uc_337;
wire uc_338;
wire uc_339;
wire uc_340;
wire uc_341;
wire uc_342;
wire uc_343;
wire uc_344;
wire uc_345;
wire uc_346;
wire uc_347;
wire uc_348;
wire uc_349;
wire uc_350;
wire uc_351;
wire uc_352;
wire uc_353;
wire uc_354;
wire uc_355;
wire uc_356;
wire uc_357;
wire uc_358;
wire uc_359;
wire uc_360;
wire uc_361;
wire uc_362;
wire uc_363;
wire uc_364;
wire uc_365;
wire uc_366;
wire uc_367;
wire uc_368;
wire uc_369;
wire uc_370;
wire uc_371;
wire uc_372;
wire uc_373;
wire uc_374;
wire uc_375;
wire uc_376;
wire uc_377;
wire uc_378;
wire uc_379;
wire uc_380;
wire uc_381;
wire uc_382;
wire uc_383;
wire uc_384;
wire uc_385;
wire uc_386;
wire uc_387;
wire uc_388;
wire uc_389;
wire uc_390;
wire uc_391;
wire uc_392;
wire uc_393;
wire uc_394;
wire uc_395;
wire uc_396;
wire uc_397;
wire uc_398;
wire uc_399;
wire uc_400;
wire uc_401;
wire uc_402;
wire uc_403;
wire uc_404;
wire uc_405;
wire uc_406;
wire uc_407;
wire uc_408;
wire uc_409;
wire uc_410;
wire uc_411;
wire uc_412;
wire uc_413;
wire uc_414;
wire uc_415;
wire uc_416;
wire uc_417;
wire uc_418;
wire uc_419;
wire uc_420;
wire uc_421;
wire uc_422;
wire uc_423;
wire uc_424;
wire uc_425;
wire uc_426;
wire uc_427;
wire uc_428;
wire uc_429;
wire uc_430;
wire uc_431;
wire uc_432;
wire uc_433;
wire uc_434;
wire uc_435;
wire uc_436;
wire uc_437;
wire uc_438;
wire uc_439;
wire uc_440;
wire uc_441;
wire uc_442;
wire uc_443;
wire uc_444;
wire uc_445;
wire uc_446;
wire uc_447;
wire uc_448;
wire uc_449;
wire uc_450;
wire uc_451;
wire uc_452;
wire uc_453;
wire uc_454;
wire uc_455;
wire uc_456;
wire uc_457;
wire uc_458;
wire uc_459;
wire uc_460;
wire uc_461;
wire uc_462;
wire uc_463;
wire uc_464;
wire uc_465;
wire uc_466;
wire uc_467;
wire uc_468;
wire uc_469;
wire uc_470;
wire uc_471;
wire uc_472;
wire uc_473;
wire uc_474;
wire uc_475;
wire uc_476;
wire uc_477;
wire uc_478;
wire uc_479;
wire uc_480;
wire uc_481;
wire uc_482;
wire uc_483;
wire uc_484;
wire uc_485;
wire uc_486;
wire uc_487;
wire uc_488;
wire uc_489;
wire uc_490;
wire uc_491;
wire uc_492;
wire uc_493;
wire uc_494;
wire uc_495;
wire uc_496;
wire uc_497;
wire uc_498;
wire uc_499;
wire uc_500;
wire uc_501;
wire uc_502;
wire uc_503;
wire uc_504;
wire uc_505;
wire uc_506;
wire uc_507;
wire uc_508;
wire uc_509;
wire uc_510;
wire uc_511;
wire uc_512;
wire uc_513;
wire uc_514;
wire uc_515;
wire uc_516;
wire uc_517;
wire uc_518;
wire uc_519;
wire uc_520;
wire uc_521;
wire uc_522;
wire uc_523;
wire uc_524;
wire uc_525;
wire uc_526;
wire uc_527;
wire uc_528;
wire uc_529;
wire uc_530;
wire uc_531;
wire uc_532;
wire uc_533;
wire uc_534;
wire uc_535;
wire uc_536;
wire uc_537;
wire uc_538;
wire uc_539;
wire uc_540;
wire uc_541;
wire uc_542;
wire uc_543;
wire uc_544;
wire uc_545;
wire uc_546;
wire uc_547;
wire uc_548;
wire uc_549;
wire uc_550;
wire uc_551;
wire uc_552;
wire uc_553;
wire uc_554;
wire uc_555;
wire uc_556;
wire uc_557;
wire uc_558;
wire uc_559;
wire uc_560;
wire uc_561;
wire uc_562;
wire uc_563;
wire uc_564;
wire uc_565;
wire uc_566;
wire uc_567;
wire uc_568;
wire uc_569;
wire uc_570;
wire uc_571;
wire uc_572;
wire uc_573;
wire uc_574;
wire uc_575;
wire uc_576;
wire uc_577;
wire uc_578;
wire uc_579;
wire uc_580;
wire uc_581;
wire uc_582;
wire uc_583;
wire uc_584;
wire uc_585;
wire uc_586;
wire uc_587;
wire uc_588;
wire uc_589;
wire uc_590;
wire uc_591;
wire uc_592;
wire uc_593;
wire uc_594;
wire uc_595;
wire uc_596;
wire uc_597;
wire uc_598;
wire uc_599;
wire uc_600;
wire uc_601;
wire uc_602;
wire uc_603;
wire uc_604;
wire uc_605;
wire uc_606;
wire uc_607;
wire uc_608;
wire uc_609;
wire uc_610;
wire uc_611;
wire uc_612;
wire uc_613;
wire uc_614;
wire uc_615;
wire uc_616;
wire uc_617;
wire uc_618;
wire uc_619;
wire uc_620;
wire uc_621;
wire uc_622;
wire uc_623;
wire uc_624;
wire uc_625;
wire uc_626;
wire uc_627;
wire uc_628;
wire uc_629;
wire uc_630;
wire uc_631;
wire uc_632;
wire uc_633;
wire uc_634;
wire uc_635;
wire uc_636;
wire uc_637;
wire uc_638;
wire uc_639;
wire uc_640;
wire uc_641;
wire uc_642;
wire uc_643;
wire uc_644;
wire uc_645;
wire uc_646;
wire uc_647;
wire uc_648;
wire uc_649;
wire uc_650;
wire uc_651;
wire uc_652;
wire uc_653;
wire uc_654;
wire uc_655;
wire uc_656;
wire uc_657;
wire uc_658;
wire uc_659;
wire uc_660;
wire uc_661;
wire uc_662;
wire uc_663;
wire uc_664;
wire uc_665;
wire uc_666;
wire uc_667;
wire uc_668;
wire uc_669;
wire uc_670;
wire uc_671;
wire uc_672;
wire uc_673;
wire uc_674;
wire uc_675;
wire uc_676;
wire uc_677;
wire uc_678;
wire uc_679;
wire uc_680;
wire uc_681;
wire uc_682;
wire uc_683;
wire uc_684;
wire uc_685;
wire uc_686;
wire uc_687;
wire uc_688;
wire uc_689;
wire uc_690;
wire uc_691;
wire uc_692;
wire uc_693;
wire uc_694;
wire uc_695;
wire uc_696;
wire uc_697;
wire uc_698;
wire uc_699;
wire uc_700;
wire uc_701;
wire uc_702;
wire uc_703;
wire uc_704;
wire uc_705;
wire uc_706;
wire uc_707;
wire uc_708;
wire uc_709;
wire uc_710;
wire uc_711;
wire uc_712;
wire uc_713;
wire uc_714;
wire uc_715;
wire uc_716;
wire uc_717;
wire uc_718;
wire uc_719;
wire uc_720;
wire uc_721;
wire uc_722;
wire uc_723;
wire uc_724;
wire uc_725;
wire uc_726;
wire uc_727;
wire uc_728;
wire uc_729;
wire uc_730;
wire uc_731;
wire uc_732;
wire uc_733;
wire uc_734;
wire uc_735;
wire uc_736;
wire uc_737;
wire uc_738;
wire uc_739;
wire uc_740;
wire uc_741;
wire uc_742;
wire uc_743;
wire uc_744;
wire uc_745;
wire uc_746;
wire uc_747;
wire uc_748;
wire uc_749;
wire uc_750;
wire uc_751;
wire uc_752;
wire uc_753;
wire uc_754;
wire uc_755;
wire uc_756;
wire uc_757;
wire uc_758;
wire uc_759;
wire uc_760;
wire uc_761;
wire uc_762;
wire uc_763;
wire uc_764;
wire uc_765;
wire uc_766;
wire uc_767;
wire uc_768;
wire uc_769;
wire uc_770;
wire uc_771;
wire uc_772;
wire uc_773;
wire uc_774;
wire uc_775;
wire uc_776;
wire uc_777;
wire uc_778;
wire uc_779;
wire uc_780;
wire uc_781;
wire uc_782;
wire uc_783;
wire uc_784;
wire uc_785;
wire uc_786;
wire uc_787;
wire uc_788;
wire uc_789;
wire uc_790;
wire uc_791;
wire uc_792;
wire uc_793;
wire uc_794;
wire uc_795;
wire uc_796;
wire uc_797;
wire uc_798;
wire uc_799;
wire uc_800;
wire uc_801;
wire uc_802;
wire uc_803;
wire uc_804;
wire uc_805;
wire uc_806;
wire uc_807;
wire uc_808;
wire uc_809;
wire uc_810;
wire uc_811;
wire uc_812;
wire uc_813;
wire uc_814;
wire uc_815;
wire uc_816;
wire uc_817;
wire uc_818;
wire uc_819;
wire uc_820;
wire uc_821;
wire uc_822;
wire uc_823;
wire uc_824;
wire uc_825;
wire uc_826;
wire uc_827;
wire uc_828;
wire uc_829;
wire uc_830;
wire uc_831;
wire uc_832;
wire uc_833;
wire uc_834;
wire uc_835;
wire uc_836;
wire uc_837;
wire uc_838;
wire uc_839;
wire uc_840;
wire uc_841;
wire uc_842;
wire uc_843;
wire uc_844;
wire uc_845;
wire uc_846;
wire uc_847;
wire uc_848;
wire uc_849;
wire uc_850;
wire uc_851;
wire uc_852;
wire uc_853;
wire uc_854;
wire uc_855;
wire uc_856;
wire uc_857;
wire uc_858;
wire uc_859;
wire uc_860;
wire uc_861;
wire uc_862;
wire uc_863;
wire uc_864;
wire uc_865;
wire uc_866;
wire uc_867;
wire uc_868;
wire uc_869;
wire uc_870;
wire uc_871;
wire uc_872;
wire uc_873;
wire uc_874;
wire uc_875;
wire uc_876;
wire uc_877;
wire uc_878;
wire uc_879;
wire uc_880;
wire uc_881;
wire uc_882;
wire uc_883;
wire uc_884;
wire uc_885;
wire uc_886;
wire uc_887;
wire uc_888;
wire uc_889;
wire uc_890;
wire uc_891;
wire uc_892;
wire uc_893;
wire uc_894;
wire uc_895;
wire uc_896;
wire uc_897;
wire uc_898;
wire uc_899;
wire uc_900;
wire uc_901;
wire uc_902;
wire uc_903;
wire uc_904;
wire uc_905;
wire uc_906;
wire uc_907;
wire uc_908;
wire uc_909;
wire uc_910;
wire uc_911;
wire uc_912;
wire uc_913;
wire uc_914;
wire uc_915;
wire uc_916;
wire uc_917;
wire uc_918;
wire uc_919;
wire uc_920;
wire uc_921;
wire uc_922;
wire uc_923;
wire uc_924;
wire uc_925;
wire uc_926;
wire uc_927;
wire uc_928;
wire uc_929;
wire uc_930;
wire uc_931;
wire uc_932;
wire uc_933;
wire uc_934;
wire uc_935;
wire uc_936;
wire uc_937;
wire uc_938;
wire uc_939;
wire uc_940;
wire uc_941;
wire uc_942;
wire uc_943;
wire uc_944;
wire uc_945;
wire uc_946;
wire uc_947;
wire uc_948;
wire uc_949;
wire uc_950;
wire uc_951;
wire uc_952;
wire uc_953;
wire uc_954;
wire uc_955;
wire uc_956;
wire uc_957;
wire uc_958;
wire uc_959;
wire uc_960;
wire uc_961;
wire uc_962;
wire uc_963;
wire uc_964;
wire uc_965;
wire uc_966;
wire uc_967;
wire uc_968;
wire uc_969;
wire uc_970;
wire uc_971;
wire uc_972;
wire uc_973;
wire uc_974;
wire uc_975;
wire uc_976;
wire uc_977;
wire uc_978;
wire uc_979;
wire uc_980;
wire uc_981;
wire uc_982;
wire uc_983;
wire uc_984;
wire uc_985;
wire uc_986;
wire uc_987;
wire uc_988;
wire uc_989;
wire uc_990;
wire uc_991;
wire uc_992;
wire uc_993;
wire uc_994;
wire uc_995;
wire uc_996;
wire uc_997;
wire uc_998;
wire uc_999;
wire uc_1000;
wire uc_1001;
wire uc_1002;
wire uc_1003;
wire uc_1004;
wire uc_1005;
wire uc_1006;
wire uc_1007;
wire uc_1008;
wire uc_1009;
wire uc_1010;
wire uc_1011;
wire uc_1012;
wire uc_1013;
wire uc_1014;
wire uc_1015;
wire uc_1016;
wire uc_1017;
wire uc_1018;
wire uc_1019;
wire uc_1020;
wire uc_1021;
wire uc_1022;
wire uc_1023;
wire uc_1024;
wire uc_1025;
wire uc_1026;
wire uc_1027;
wire uc_1028;
wire uc_1029;
wire uc_1030;
wire uc_1031;
wire uc_1032;
wire uc_1033;
wire uc_1034;
wire uc_1035;
wire uc_1036;
wire uc_1037;
wire uc_1038;
wire uc_1039;
wire uc_1040;
wire uc_1041;
wire uc_1042;
wire uc_1043;
wire uc_1044;
wire uc_1045;
wire uc_1046;
wire uc_1047;
wire uc_1048;
wire uc_1049;
wire uc_1050;
wire uc_1051;
wire uc_1052;
wire uc_1053;
wire uc_1054;
wire uc_1055;
wire uc_1056;
wire uc_1057;
wire uc_1058;
wire uc_1059;
wire uc_1060;
wire uc_1061;
wire uc_1062;
wire uc_1063;
wire uc_1064;
wire uc_1065;
wire uc_1066;
wire uc_1067;
wire uc_1068;
wire uc_1069;
wire uc_1070;
wire uc_1071;
wire uc_1072;
wire uc_1073;
wire uc_1074;
wire uc_1075;
wire uc_1076;
wire uc_1077;
wire uc_1078;
wire uc_1079;
wire uc_1080;
wire uc_1081;
wire uc_1082;
wire uc_1083;
wire uc_1084;
wire uc_1085;
wire uc_1086;
wire uc_1087;
wire uc_1088;
wire uc_1089;
wire uc_1090;
wire uc_1091;
wire uc_1092;
wire uc_1093;
wire uc_1094;
wire uc_1095;
wire uc_1096;
wire uc_1097;
wire uc_1098;
wire uc_1099;
wire uc_1100;
wire uc_1101;
wire uc_1102;
wire uc_1103;
wire uc_1104;
wire uc_1105;
wire uc_1106;
wire uc_1107;
wire uc_1108;
wire uc_1109;
wire uc_1110;
wire uc_1111;
wire uc_1112;
wire uc_1113;
wire uc_1114;
wire uc_1115;
wire uc_1116;
wire uc_1117;
wire uc_1118;
wire uc_1119;
wire uc_1120;
wire uc_1121;
wire uc_1122;
wire uc_1123;
wire uc_1124;
wire uc_1125;
wire uc_1126;
wire uc_1127;
wire uc_1128;
wire uc_1129;
wire uc_1130;
wire uc_1131;
wire uc_1132;
wire uc_1133;
wire uc_1134;
wire uc_1135;
wire uc_1136;
wire uc_1137;
wire uc_1138;
wire uc_1139;
wire uc_1140;
wire uc_1141;
wire uc_1142;
wire uc_1143;
wire uc_1144;
wire uc_1145;
wire uc_1146;
wire uc_1147;
wire uc_1148;
wire uc_1149;
wire uc_1150;
wire uc_1151;
wire uc_1152;
wire uc_1153;
wire uc_1154;
wire uc_1155;
wire uc_1156;
wire uc_1157;
wire uc_1158;
wire uc_1159;
wire uc_1160;
wire uc_1161;
wire uc_1162;
wire uc_1163;
wire uc_1164;
wire uc_1165;
wire uc_1166;
wire uc_1167;
wire uc_1168;
wire uc_1169;
wire uc_1170;
wire uc_1171;
wire uc_1172;
wire uc_1173;
wire uc_1174;
wire uc_1175;
wire uc_1176;
wire uc_1177;
wire uc_1178;
wire uc_1179;
wire uc_1180;
wire uc_1181;
wire uc_1182;
wire uc_1183;
wire uc_1184;
wire uc_1185;
wire uc_1186;
wire uc_1187;
wire uc_1188;
wire uc_1189;
wire uc_1190;
wire uc_1191;
wire uc_1192;
wire uc_1193;
wire uc_1194;
wire uc_1195;
wire uc_1196;
wire uc_1197;
wire uc_1198;
wire uc_1199;
wire uc_1200;
wire uc_1201;
wire uc_1202;
wire uc_1203;
wire uc_1204;
wire uc_1205;
wire uc_1206;
wire uc_1207;
wire uc_1208;
wire uc_1209;
wire uc_1210;
wire uc_1211;
wire uc_1212;
wire uc_1213;
wire uc_1214;
wire uc_1215;
wire uc_1216;
wire uc_1217;
wire uc_1218;
wire uc_1219;
wire uc_1220;
wire uc_1221;
wire uc_1222;
wire uc_1223;
wire uc_1224;
wire uc_1225;
wire uc_1226;
wire uc_1227;
wire uc_1228;
wire uc_1229;
wire uc_1230;
wire uc_1231;
wire uc_1232;
wire uc_1233;
wire uc_1234;
wire uc_1235;
wire uc_1236;
wire uc_1237;
wire uc_1238;
wire uc_1239;
wire uc_1240;
wire uc_1241;
wire uc_1242;
wire uc_1243;
wire uc_1244;
wire uc_1245;
wire uc_1246;
wire uc_1247;
wire uc_1248;
wire uc_1249;
wire uc_1250;
wire uc_1251;
wire uc_1252;
wire uc_1253;
wire uc_1254;
wire uc_1255;
wire uc_1256;
wire uc_1257;
wire uc_1258;
wire uc_1259;
wire uc_1260;
wire uc_1261;
wire uc_1262;
wire uc_1263;
wire uc_1264;
wire uc_1265;
wire uc_1266;
wire uc_1267;
wire uc_1268;
wire uc_1269;
wire uc_1270;
wire uc_1271;
wire uc_1272;
wire uc_1273;
wire uc_1274;
wire uc_1275;
wire uc_1276;
wire uc_1277;
wire uc_1278;
wire uc_1279;
wire uc_1280;
wire uc_1281;
wire uc_1282;
wire uc_1283;
wire uc_1284;
wire uc_1285;
wire uc_1286;
wire uc_1287;
wire uc_1288;
wire uc_1289;
wire uc_1290;
wire uc_1291;
wire uc_1292;
wire uc_1293;
wire uc_1294;
wire uc_1295;
wire uc_1296;
wire uc_1297;
wire uc_1298;
wire uc_1299;
wire uc_1300;
wire uc_1301;
wire uc_1302;
wire uc_1303;
wire uc_1304;
wire uc_1305;
wire uc_1306;
wire uc_1307;
wire uc_1308;
wire uc_1309;
wire uc_1310;
wire uc_1311;
wire uc_1312;
wire uc_1313;
wire uc_1314;
wire uc_1315;
wire uc_1316;
wire uc_1317;
wire uc_1318;
wire uc_1319;
wire uc_1320;
wire uc_1321;
wire uc_1322;
wire uc_1323;
wire uc_1324;
wire uc_1325;
wire uc_1326;
wire uc_1327;
wire uc_1328;
wire uc_1329;
wire uc_1330;
wire uc_1331;
wire uc_1332;
wire uc_1333;
wire uc_1334;
wire uc_1335;
wire uc_1336;
wire uc_1337;
wire uc_1338;
wire uc_1339;
wire uc_1340;
wire uc_1341;
wire uc_1342;
wire uc_1343;
wire uc_1344;
wire uc_1345;
wire uc_1346;
wire uc_1347;
wire uc_1348;
wire uc_1349;
wire uc_1350;
wire uc_1351;
wire uc_1352;
wire uc_1353;
wire uc_1354;
wire uc_1355;
wire uc_1356;
wire uc_1357;
wire uc_1358;
wire uc_1359;
wire uc_1360;
wire uc_1361;
wire uc_1362;
wire uc_1363;
wire uc_1364;
wire uc_1365;
wire uc_1366;
wire uc_1367;
wire uc_1368;
wire uc_1369;
wire uc_1370;
wire uc_1371;
wire uc_1372;
wire uc_1373;
wire uc_1374;
wire uc_1375;
wire uc_1376;
wire uc_1377;
wire uc_1378;
wire uc_1379;
wire uc_1380;
wire uc_1381;
wire uc_1382;
wire uc_1383;
wire uc_1384;
wire uc_1385;
wire uc_1386;
wire uc_1387;
wire uc_1388;
wire uc_1389;
wire uc_1390;
wire uc_1391;
wire uc_1392;
wire uc_1393;
wire uc_1394;
wire uc_1395;
wire uc_1396;
wire uc_1397;
wire uc_1398;
wire uc_1399;
wire uc_1400;
wire uc_1401;
wire uc_1402;
wire uc_1403;
wire uc_1404;
wire uc_1405;
wire uc_1406;
wire uc_1407;
wire uc_1408;
wire uc_1409;
wire uc_1410;
wire uc_1411;
wire uc_1412;
wire uc_1413;
wire uc_1414;
wire uc_1415;
wire uc_1416;
wire uc_1417;
wire uc_1418;
wire uc_1419;
wire uc_1420;
wire uc_1421;
wire uc_1422;
wire uc_1423;
wire uc_1424;
wire uc_1425;
wire uc_1426;
wire uc_1427;
wire uc_1428;
wire uc_1429;
wire uc_1430;
wire uc_1431;
wire uc_1432;
wire uc_1433;
wire uc_1434;
wire uc_1435;
wire uc_1436;
wire uc_1437;
wire uc_1438;
wire uc_1439;
wire uc_1440;
wire uc_1441;
wire uc_1442;
wire uc_1443;
wire uc_1444;
wire uc_1445;
wire uc_1446;
wire uc_1447;
wire uc_1448;
wire uc_1449;
wire uc_1450;
wire uc_1451;
wire uc_1452;
wire uc_1453;
wire uc_1454;
wire uc_1455;
wire uc_1456;
wire uc_1457;
wire uc_1458;
wire uc_1459;
wire uc_1460;
wire uc_1461;
wire uc_1462;
wire uc_1463;
wire uc_1464;
wire uc_1465;
wire uc_1466;
wire uc_1467;
wire uc_1468;
wire uc_1469;
wire uc_1470;
wire uc_1471;
wire uc_1472;
wire uc_1473;
wire uc_1474;
wire uc_1475;
wire uc_1476;
wire uc_1477;
wire uc_1478;
wire uc_1479;
wire uc_1480;
wire uc_1481;
wire uc_1482;
wire uc_1483;
wire uc_1484;
wire uc_1485;
wire uc_1486;
wire uc_1487;
wire uc_1488;
wire uc_1489;
wire uc_1490;
wire uc_1491;
wire uc_1492;
wire uc_1493;
wire uc_1494;
wire uc_1495;
wire uc_1496;
wire uc_1497;
wire uc_1498;
wire uc_1499;
wire uc_1500;
wire uc_1501;
wire uc_1502;
wire uc_1503;
wire uc_1504;
wire uc_1505;
wire uc_1506;
wire uc_1507;
wire uc_1508;
wire uc_1509;
wire uc_1510;
wire uc_1511;
wire uc_1512;
wire uc_1513;
wire uc_1514;
wire uc_1515;
wire uc_1516;
wire uc_1517;
wire uc_1518;
wire uc_1519;
wire uc_1520;
wire uc_1521;
wire uc_1522;
wire uc_1523;
wire uc_1524;
wire uc_1525;
wire uc_1526;
wire uc_1527;
wire uc_1528;
wire uc_1529;
wire uc_1530;
wire uc_1531;
wire uc_1532;
wire uc_1533;
wire uc_1534;
wire uc_1535;
wire uc_1536;
wire uc_1537;
wire uc_1538;
wire uc_1539;
wire uc_1540;
wire uc_1541;
wire uc_1542;
wire uc_1543;
wire uc_1544;
wire uc_1545;
wire uc_1546;
wire uc_1547;
wire uc_1548;
wire uc_1549;
wire uc_1550;
wire uc_1551;
wire uc_1552;
wire uc_1553;
wire uc_1554;
wire uc_1555;
wire uc_1556;
wire uc_1557;
wire uc_1558;
wire uc_1559;
wire uc_1560;
wire uc_1561;
wire uc_1562;
wire uc_1563;
wire uc_1564;
wire uc_1565;
wire uc_1566;
wire uc_1567;
wire uc_1568;
wire uc_1569;
wire uc_1570;
wire uc_1571;
wire uc_1572;
wire uc_1573;
wire uc_1574;
wire uc_1575;
wire uc_1576;
wire uc_1577;
wire uc_1578;
wire uc_1579;
wire uc_1580;
wire uc_1581;
wire uc_1582;
wire uc_1583;
wire uc_1584;
wire uc_1585;
wire uc_1586;
wire uc_1587;
wire uc_1588;
wire uc_1589;
wire uc_1590;
wire uc_1591;
wire uc_1592;
wire uc_1593;
wire uc_1594;
wire uc_1595;
wire uc_1596;
wire uc_1597;
wire uc_1598;
wire uc_1599;
wire uc_1600;
wire uc_1601;
wire uc_1602;
wire uc_1603;
wire uc_1604;
wire uc_1605;
wire uc_1606;
wire uc_1607;
wire uc_1608;
wire uc_1609;
wire uc_1610;
wire uc_1611;
wire uc_1612;
wire uc_1613;
wire uc_1614;
wire uc_1615;
wire uc_1616;
wire uc_1617;
wire uc_1618;
wire uc_1619;
wire uc_1620;
wire uc_1621;
wire uc_1622;
wire uc_1623;
wire uc_1624;
wire uc_1625;
wire uc_1626;
wire uc_1627;
wire uc_1628;
wire uc_1629;
wire uc_1630;
wire uc_1631;
wire uc_1632;
wire uc_1633;
wire uc_1634;
wire uc_1635;
wire uc_1636;
wire uc_1637;
wire uc_1638;
wire uc_1639;
wire uc_1640;
wire uc_1641;
wire uc_1642;
wire uc_1643;
wire uc_1644;
wire uc_1645;
wire uc_1646;
wire uc_1647;
wire uc_1648;
wire uc_1649;
wire uc_1650;
wire uc_1651;
wire uc_1652;
wire uc_1653;
wire uc_1654;
wire uc_1655;
wire uc_1656;
wire uc_1657;
wire uc_1658;
wire uc_1659;
wire uc_1660;
wire uc_1661;
wire uc_1662;
wire uc_1663;
wire uc_1664;
wire uc_1665;
wire uc_1666;
wire uc_1667;
wire uc_1668;
wire uc_1669;
wire uc_1670;
wire uc_1671;
wire uc_1672;
wire uc_1673;
wire uc_1674;
wire uc_1675;
wire uc_1676;
wire uc_1677;
wire uc_1678;
wire uc_1679;
wire uc_1680;
wire uc_1681;
wire uc_1682;
wire uc_1683;
wire uc_1684;
wire uc_1685;
wire uc_1686;
wire uc_1687;
wire uc_1688;
wire uc_1689;
wire uc_1690;
wire uc_1691;
wire uc_1692;
wire uc_1693;
wire uc_1694;
wire uc_1695;
wire uc_1696;
wire uc_1697;
wire uc_1698;
wire uc_1699;
wire uc_1700;
wire uc_1701;
wire uc_1702;
wire uc_1703;
wire uc_1704;
wire uc_1705;
wire uc_1706;
wire uc_1707;
wire uc_1708;
wire uc_1709;
wire uc_1710;
wire uc_1711;
wire uc_1712;
wire uc_1713;
wire uc_1714;
wire uc_1715;
wire uc_1716;
wire uc_1717;
wire uc_1718;
wire uc_1719;
wire uc_1720;
wire uc_1721;
wire uc_1722;
wire uc_1723;
wire uc_1724;
wire uc_1725;
wire uc_1726;
wire uc_1727;
wire uc_1728;
wire uc_1729;
wire uc_1730;
wire uc_1731;
wire uc_1732;
wire uc_1733;
wire uc_1734;
wire uc_1735;
wire uc_1736;
wire uc_1737;
wire uc_1738;
wire uc_1739;
wire uc_1740;
wire uc_1741;
wire uc_1742;
wire uc_1743;
wire uc_1744;
wire uc_1745;
wire uc_1746;
wire uc_1747;
wire uc_1748;
wire uc_1749;
wire uc_1750;
wire uc_1751;
wire uc_1752;
wire uc_1753;
wire uc_1754;
wire uc_1755;
wire uc_1756;
wire uc_1757;
wire uc_1758;
wire uc_1759;
wire uc_1760;
wire uc_1761;
wire uc_1762;
wire uc_1763;
wire uc_1764;
wire uc_1765;
wire uc_1766;
wire uc_1767;
wire uc_1768;
wire uc_1769;
wire uc_1770;
wire uc_1771;
wire uc_1772;
wire uc_1773;
wire uc_1774;
wire uc_1775;
wire uc_1776;
wire uc_1777;
wire uc_1778;
wire uc_1779;
wire uc_1780;
wire uc_1781;
wire uc_1782;
wire uc_1783;
wire uc_1784;
wire uc_1785;
wire uc_1786;
wire uc_1787;
wire uc_1788;
wire uc_1789;
wire uc_1790;
wire uc_1791;
wire uc_1792;
wire uc_1793;
wire uc_1794;
wire uc_1795;
wire uc_1796;
wire uc_1797;
wire uc_1798;
wire uc_1799;
wire uc_1800;
wire uc_1801;
wire uc_1802;
wire uc_1803;
wire uc_1804;
wire uc_1805;
wire uc_1806;
wire uc_1807;
wire uc_1808;
wire uc_1809;
wire uc_1810;
wire uc_1811;
wire uc_1812;
wire uc_1813;
wire uc_1814;
wire uc_1815;
wire uc_1816;
wire uc_1817;
wire uc_1818;
wire uc_1819;
wire uc_1820;
wire uc_1821;
wire uc_1822;
wire uc_1823;
wire uc_1824;
wire uc_1825;
wire uc_1826;
wire uc_1827;
wire uc_1828;
wire uc_1829;
wire uc_1830;
wire uc_1831;
wire uc_1832;
wire uc_1833;
wire uc_1834;
wire uc_1835;
wire uc_1836;
wire uc_1837;
wire uc_1838;
wire uc_1839;
wire uc_1840;
wire uc_1841;
wire uc_1842;
wire uc_1843;
wire uc_1844;
wire uc_1845;
wire uc_1846;
wire uc_1847;
wire uc_1848;
wire uc_1849;
wire uc_1850;
wire uc_1851;
wire uc_1852;
wire uc_1853;
wire uc_1854;
wire uc_1855;
wire uc_1856;
wire uc_1857;
wire uc_1858;
wire uc_1859;
wire uc_1860;
wire uc_1861;
wire uc_1862;
wire uc_1863;
wire uc_1864;
wire uc_1865;
wire uc_1866;
wire uc_1867;
wire uc_1868;
wire uc_1869;
wire uc_1870;
wire uc_1871;
wire uc_1872;
wire uc_1873;
wire uc_1874;
wire uc_1875;
wire uc_1876;
wire uc_1877;
wire uc_1878;
wire uc_1879;
wire uc_1880;
wire uc_1881;
wire uc_1882;
wire uc_1883;
wire uc_1884;
wire uc_1885;
wire uc_1886;
wire uc_1887;
wire uc_1888;
wire uc_1889;
wire uc_1890;
wire uc_1891;
wire uc_1892;
wire uc_1893;
wire uc_1894;
wire uc_1895;
wire uc_1896;
wire uc_1897;
wire uc_1898;
wire uc_1899;
wire uc_1900;
wire uc_1901;
wire uc_1902;
wire uc_1903;
wire uc_1904;
wire uc_1905;
wire uc_1906;
wire uc_1907;
wire uc_1908;
wire uc_1909;
wire uc_1910;
wire uc_1911;
wire uc_1912;
wire uc_1913;
wire uc_1914;
wire uc_1915;
wire uc_1916;
wire uc_1917;
wire uc_1918;
wire uc_1919;
wire uc_1920;
wire uc_1921;
wire uc_1922;
wire uc_1923;
wire uc_1924;
wire uc_1925;
wire uc_1926;
wire uc_1927;
wire uc_1928;
wire uc_1929;
wire uc_1930;
wire uc_1931;
wire uc_1932;
wire uc_1933;
wire uc_1934;
wire uc_1935;
wire uc_1936;
wire uc_1937;
wire uc_1938;
wire uc_1939;
wire uc_1940;
wire uc_1941;
wire uc_1942;
wire uc_1943;
wire uc_1944;
wire uc_1945;
wire uc_1946;
wire uc_1947;
wire uc_1948;
wire uc_1949;
wire uc_1950;
wire uc_1951;
wire uc_1952;
wire uc_1953;
wire uc_1954;
wire uc_1955;
wire uc_1956;
wire uc_1957;
wire uc_1958;
wire uc_1959;
wire uc_1960;
wire uc_1961;
wire uc_1962;
wire uc_1963;
wire uc_1964;
wire uc_1965;
wire uc_1966;
wire uc_1967;
wire uc_1968;
wire uc_1969;
wire uc_1970;
wire uc_1971;
wire uc_1972;
wire uc_1973;
wire uc_1974;
wire uc_1975;
wire uc_1976;
wire uc_1977;
wire uc_1978;
wire uc_1979;
wire uc_1980;
wire uc_1981;
wire uc_1982;
wire uc_1983;
wire uc_1984;
wire uc_1985;
wire uc_1986;
wire uc_1987;
wire uc_1988;
wire uc_1989;
wire uc_1990;
wire uc_1991;
wire uc_1992;
wire uc_1993;
wire uc_1994;
wire uc_1995;
wire uc_1996;
wire uc_1997;
wire uc_1998;
wire uc_1999;
wire uc_2000;
wire uc_2001;
wire uc_2002;
wire uc_2003;
wire uc_2004;
wire uc_2005;
wire uc_2006;
wire uc_2007;
wire uc_2008;
wire uc_2009;
wire uc_2010;
wire uc_2011;
wire uc_2012;
wire uc_2013;
wire uc_2014;
wire uc_2015;
wire uc_2016;
wire uc_2017;
wire uc_2018;
wire uc_2019;
wire uc_2020;
wire uc_2021;
wire uc_2022;
wire uc_2023;
wire uc_2024;
wire uc_2025;
wire uc_2026;
wire uc_2027;
wire uc_2028;
wire uc_2029;
wire uc_2030;
wire uc_2031;
wire uc_2032;
wire uc_2033;
wire uc_2034;
wire uc_2035;
wire uc_2036;
wire uc_2037;
wire uc_2038;
wire uc_2039;
wire uc_2040;
wire uc_2041;
wire uc_2042;
wire uc_2043;
wire uc_2044;
wire uc_2045;
wire uc_2046;
wire uc_2047;
wire uc_2048;
wire uc_2049;
wire uc_2050;
wire uc_2051;
wire uc_2052;
wire uc_2053;
wire uc_2054;
wire uc_2055;
wire uc_2056;
wire uc_2057;
wire uc_2058;
wire uc_2059;
wire uc_2060;
wire uc_2061;
wire uc_2062;
wire uc_2063;
wire uc_2064;
wire uc_2065;
wire uc_2066;
wire uc_2067;
wire uc_2068;
wire uc_2069;
wire uc_2070;
wire uc_2071;
wire uc_2072;
wire uc_2073;
wire uc_2074;
wire uc_2075;
wire uc_2076;
wire uc_2077;
wire uc_2078;
wire uc_2079;
wire uc_2080;
wire uc_2081;
wire uc_2082;
wire uc_2083;
wire uc_2084;
wire uc_2085;
wire uc_2086;
wire uc_2087;
wire uc_2088;
wire uc_2089;
wire uc_2090;
wire uc_2091;
wire uc_2092;
wire uc_2093;
wire uc_2094;
wire uc_2095;
wire uc_2096;
wire uc_2097;
wire uc_2098;
wire uc_2099;
wire uc_2100;
wire uc_2101;
wire uc_2102;
wire uc_2103;
wire uc_2104;
wire uc_2105;
wire uc_2106;
wire uc_2107;
wire uc_2108;
wire uc_2109;
wire uc_2110;
wire uc_2111;
wire uc_2112;
wire uc_2113;
wire uc_2114;
wire uc_2115;
wire uc_2116;
wire uc_2117;
wire uc_2118;
wire uc_2119;
wire uc_2120;
wire uc_2121;
wire uc_2122;
wire uc_2123;
wire uc_2124;
wire uc_2125;
wire uc_2126;
wire uc_2127;
wire uc_2128;
wire uc_2129;
wire uc_2130;
wire uc_2131;
wire uc_2132;
wire uc_2133;
wire uc_2134;
wire uc_2135;
wire uc_2136;
wire uc_2137;
wire uc_2138;
wire uc_2139;
wire uc_2140;
wire uc_2141;
wire uc_2142;
wire uc_2143;
wire uc_2144;
wire uc_2145;
wire uc_2146;
wire uc_2147;
wire uc_2148;
wire uc_2149;
wire uc_2150;
wire uc_2151;
wire uc_2152;
wire uc_2153;
wire uc_2154;
wire uc_2155;
wire uc_2156;
wire uc_2157;
wire uc_2158;
wire uc_2159;
wire uc_2160;
wire uc_2161;
wire uc_2162;
wire uc_2163;
wire uc_2164;
wire uc_2165;
wire uc_2166;
wire uc_2167;
wire uc_2168;
wire uc_2169;
wire uc_2170;
wire uc_2171;
wire uc_2172;
wire uc_2173;
wire uc_2174;
wire uc_2175;
wire uc_2176;
wire uc_2177;
wire uc_2178;
wire uc_2179;
wire uc_2180;
wire uc_2181;
wire uc_2182;
wire uc_2183;
wire uc_2184;
wire uc_2185;
wire uc_2186;
wire uc_2187;
wire uc_2188;
wire uc_2189;
wire uc_2190;
wire uc_2191;
wire uc_2192;
wire uc_2193;
wire uc_2194;
wire uc_2195;
wire uc_2196;
wire uc_2197;
wire uc_2198;
wire uc_2199;
wire uc_2200;
wire uc_2201;
wire uc_2202;
wire uc_2203;
wire uc_2204;
wire uc_2205;
wire uc_2206;
wire uc_2207;
wire uc_2208;
wire uc_2209;
wire uc_2210;
wire uc_2211;
wire uc_2212;
wire uc_2213;
wire uc_2214;
wire uc_2215;
wire uc_2216;
wire uc_2217;
wire uc_2218;
wire uc_2219;
wire uc_2220;
wire uc_2221;
wire uc_2222;
wire uc_2223;
wire uc_2224;
wire uc_2225;
wire uc_2226;
wire uc_2227;
wire uc_2228;
wire uc_2229;
wire uc_2230;
wire uc_2231;
wire uc_2232;
wire uc_2233;
wire uc_2234;
wire uc_2235;
wire uc_2236;
wire uc_2237;
wire uc_2238;
wire uc_2239;
wire uc_2240;
wire uc_2241;
wire uc_2242;
wire uc_2243;
wire uc_2244;
wire uc_2245;
wire uc_2246;
wire uc_2247;
wire uc_2248;
wire uc_2249;
wire uc_2250;
wire uc_2251;
wire uc_2252;
wire uc_2253;
wire uc_2254;
wire uc_2255;
wire uc_2256;
wire uc_2257;
wire uc_2258;
wire uc_2259;
wire uc_2260;
wire uc_2261;
wire uc_2262;
wire uc_2263;
wire uc_2264;
wire uc_2265;
wire uc_2266;
wire uc_2267;
wire uc_2268;
wire uc_2269;
wire uc_2270;
wire uc_2271;
wire uc_2272;
wire uc_2273;
wire uc_2274;
wire uc_2275;
wire uc_2276;
wire uc_2277;
wire uc_2278;
wire uc_2279;
wire uc_2280;
wire uc_2281;
wire uc_2282;
wire uc_2283;
wire uc_2284;
wire uc_2285;
wire uc_2286;
wire uc_2287;
wire uc_2288;
wire uc_2289;
wire uc_2290;
wire uc_2291;
wire uc_2292;
wire uc_2293;
wire uc_2294;
wire uc_2295;
wire uc_2296;
wire uc_2297;
wire uc_2298;
wire uc_2299;
wire uc_2300;
wire uc_2301;
wire uc_2302;
wire uc_2303;
wire uc_2304;
wire uc_2305;
wire uc_2306;
wire uc_2307;
wire uc_2308;
wire uc_2309;
wire uc_2310;
wire uc_2311;
wire uc_2312;
wire uc_2313;
wire uc_2314;
wire uc_2315;
wire uc_2316;
wire uc_2317;
wire uc_2318;
wire uc_2319;
wire uc_2320;
wire uc_2321;
wire uc_2322;
wire uc_2323;
wire uc_2324;
wire uc_2325;
wire uc_2326;
wire uc_2327;
wire uc_2328;
wire uc_2329;
wire uc_2330;
wire uc_2331;
wire uc_2332;
wire uc_2333;
wire uc_2334;
wire uc_2335;
wire uc_2336;
wire uc_2337;
wire uc_2338;
wire uc_2339;
wire uc_2340;
wire uc_2341;
wire uc_2342;
wire uc_2343;
wire uc_2344;
wire uc_2345;
wire uc_2346;
wire uc_2347;
wire uc_2348;
wire uc_2349;
wire uc_2350;
wire uc_2351;
wire uc_2352;
wire uc_2353;
wire uc_2354;
wire uc_2355;
wire uc_2356;
wire uc_2357;
wire uc_2358;
wire uc_2359;
wire uc_2360;
wire uc_2361;
wire uc_2362;
wire uc_2363;
wire uc_2364;
wire uc_2365;
wire uc_2366;
wire uc_2367;
wire uc_2368;
wire uc_2369;
wire uc_2370;
wire uc_2371;
wire uc_2372;
wire uc_2373;
wire uc_2374;
wire uc_2375;
wire uc_2376;
wire uc_2377;
wire uc_2378;
wire uc_2379;
wire uc_2380;
wire uc_2381;
wire uc_2382;
wire uc_2383;
wire uc_2384;
wire uc_2385;
wire uc_2386;
wire uc_2387;
wire uc_2388;
wire uc_2389;
wire uc_2390;
wire uc_2391;
wire uc_2392;
wire uc_2393;
wire uc_2394;
wire uc_2395;
wire uc_2396;
wire uc_2397;
wire uc_2398;
wire uc_2399;
wire uc_2400;
wire uc_2401;
wire uc_2402;
wire uc_2403;
wire uc_2404;
wire uc_2405;
wire uc_2406;
wire uc_2407;
wire uc_2408;
wire uc_2409;
wire uc_2410;
wire uc_2411;
wire uc_2412;
wire uc_2413;
wire uc_2414;
wire uc_2415;
wire uc_2416;
wire uc_2417;
wire uc_2418;
wire uc_2419;
wire uc_2420;
wire uc_2421;
wire uc_2422;
wire uc_2423;
wire uc_2424;
wire uc_2425;
wire uc_2426;
wire uc_2427;
wire uc_2428;
wire uc_2429;
wire uc_2430;
wire uc_2431;
wire uc_2432;
wire uc_2433;
wire uc_2434;
wire uc_2435;
wire uc_2436;
wire uc_2437;
wire uc_2438;
wire uc_2439;
wire uc_2440;
wire uc_2441;
wire uc_2442;
wire uc_2443;
wire uc_2444;
wire uc_2445;
wire uc_2446;
wire uc_2447;
wire uc_2448;
wire uc_2449;
wire uc_2450;
wire uc_2451;
wire uc_2452;
wire uc_2453;
wire uc_2454;
wire uc_2455;
wire uc_2456;
wire uc_2457;
wire uc_2458;
wire uc_2459;
wire uc_2460;
wire uc_2461;
wire uc_2462;
wire uc_2463;
wire uc_2464;
wire uc_2465;
wire uc_2466;
wire uc_2467;
wire uc_2468;
wire uc_2469;
wire uc_2470;
wire uc_2471;
wire uc_2472;
wire uc_2473;
wire uc_2474;
wire uc_2475;
wire uc_2476;
wire uc_2477;
wire uc_2478;
wire uc_2479;
wire uc_2480;
wire uc_2481;
wire uc_2482;
wire uc_2483;
wire uc_2484;
wire uc_2485;
wire uc_2486;
wire uc_2487;
wire uc_2488;
wire uc_2489;
wire uc_2490;
wire uc_2491;
wire uc_2492;
wire uc_2493;
wire uc_2494;
wire uc_2495;
wire uc_2496;
wire uc_2497;
wire uc_2498;
wire uc_2499;
wire uc_2500;
wire uc_2501;
wire uc_2502;
wire uc_2503;
wire uc_2504;
wire uc_2505;
wire uc_2506;
wire uc_2507;
wire uc_2508;
wire uc_2509;
wire uc_2510;
wire uc_2511;
wire uc_2512;
wire uc_2513;
wire uc_2514;
wire uc_2515;
wire uc_2516;
wire uc_2517;
wire uc_2518;
wire uc_2519;
wire uc_2520;
wire uc_2521;
wire uc_2522;
wire uc_2523;
wire uc_2524;
wire uc_2525;
wire uc_2526;
wire uc_2527;
wire uc_2528;
wire uc_2529;
wire uc_2530;
wire uc_2531;
wire uc_2532;
wire uc_2533;
wire uc_2534;
wire uc_2535;
wire uc_2536;
wire uc_2537;
wire uc_2538;
wire uc_2539;
wire uc_2540;
wire uc_2541;
wire uc_2542;
wire uc_2543;
wire uc_2544;
wire uc_2545;
wire uc_2546;
wire uc_2547;
wire uc_2548;
wire uc_2549;
wire uc_2550;
wire uc_2551;
wire uc_2552;
wire uc_2553;
wire uc_2554;
wire uc_2555;
wire uc_2556;
wire uc_2557;
wire uc_2558;
wire uc_2559;
wire uc_2560;
wire uc_2561;
wire uc_2562;
wire uc_2563;
wire uc_2564;
wire uc_2565;
wire uc_2566;
wire uc_2567;
wire uc_2568;
wire uc_2569;
wire uc_2570;
wire uc_2571;
wire uc_2572;
wire uc_2573;
wire uc_2574;
wire uc_2575;
wire uc_2576;
wire uc_2577;
wire uc_2578;
wire uc_2579;
wire uc_2580;
wire uc_2581;
wire uc_2582;
wire uc_2583;
wire uc_2584;
wire uc_2585;
wire uc_2586;
wire uc_2587;
wire uc_2588;
wire uc_2589;
wire uc_2590;
wire uc_2591;
wire uc_2592;
wire uc_2593;
wire uc_2594;
wire uc_2595;
wire uc_2596;
wire uc_2597;
wire uc_2598;
wire uc_2599;
wire uc_2600;
wire uc_2601;
wire uc_2602;
wire uc_2603;
wire uc_2604;
wire uc_2605;
wire uc_2606;
wire uc_2607;
wire uc_2608;
wire uc_2609;
wire uc_2610;
wire uc_2611;
wire uc_2612;
wire uc_2613;
wire uc_2614;
wire uc_2615;
wire uc_2616;
wire uc_2617;
wire uc_2618;
wire uc_2619;
wire uc_2620;
wire uc_2621;
wire uc_2622;
wire uc_2623;
wire uc_2624;
wire uc_2625;
wire uc_2626;
wire uc_2627;
wire uc_2628;
wire uc_2629;
wire uc_2630;
wire uc_2631;
wire uc_2632;
wire uc_2633;
wire uc_2634;
wire uc_2635;
wire uc_2636;
wire uc_2637;
wire uc_2638;
wire uc_2639;
wire uc_2640;
wire uc_2641;
wire uc_2642;
wire uc_2643;
wire uc_2644;
wire uc_2645;
wire uc_2646;
wire uc_2647;
wire uc_2648;
wire uc_2649;
wire uc_2650;
wire uc_2651;
wire uc_2652;
wire uc_2653;
wire uc_2654;
wire uc_2655;
wire uc_2656;
wire uc_2657;
wire uc_2658;
wire uc_2659;
wire uc_2660;
wire uc_2661;
wire uc_2662;
wire uc_2663;
wire uc_2664;
wire uc_2665;
wire uc_2666;
wire uc_2667;
wire uc_2668;
wire uc_2669;
wire uc_2670;
wire uc_2671;
wire uc_2672;
wire uc_2673;
wire uc_2674;
wire uc_2675;
wire uc_2676;
wire uc_2677;
wire uc_2678;
wire uc_2679;
wire uc_2680;
wire uc_2681;
wire uc_2682;
wire uc_2683;
wire uc_2684;
wire uc_2685;
wire uc_2686;
wire uc_2687;
wire uc_2688;
wire uc_2689;
wire uc_2690;
wire uc_2691;
wire uc_2692;
wire uc_2693;
wire uc_2694;
wire uc_2695;
wire uc_2696;
wire uc_2697;
wire uc_2698;
wire uc_2699;
wire uc_2700;
wire uc_2701;
wire uc_2702;
wire uc_2703;
wire uc_2704;
wire uc_2705;
wire uc_2706;
wire uc_2707;
wire uc_2708;
wire uc_2709;
wire uc_2710;
wire uc_2711;
wire uc_2712;
wire uc_2713;
wire uc_2714;
wire uc_2715;
wire uc_2716;
wire uc_2717;
wire uc_2718;
wire uc_2719;
wire uc_2720;
wire uc_2721;
wire uc_2722;
wire uc_2723;
wire uc_2724;
wire uc_2725;
wire uc_2726;
wire uc_2727;
wire uc_2728;
wire uc_2729;
wire uc_2730;
wire uc_2731;
wire uc_2732;
wire uc_2733;
wire uc_2734;
wire uc_2735;
wire uc_2736;
wire uc_2737;
wire uc_2738;
wire uc_2739;
wire uc_2740;
wire uc_2741;
wire uc_2742;
wire uc_2743;
wire uc_2744;
wire uc_2745;
wire uc_2746;
wire uc_2747;
wire uc_2748;
wire uc_2749;
wire uc_2750;
wire uc_2751;
wire uc_2752;
wire uc_2753;
wire uc_2754;
wire uc_2755;
wire uc_2756;
wire uc_2757;
wire uc_2758;
wire uc_2759;
wire uc_2760;
wire uc_2761;
wire uc_2762;
wire uc_2763;
wire uc_2764;
wire uc_2765;
wire uc_2766;
wire uc_2767;
wire uc_2768;
wire uc_2769;
wire uc_2770;
wire uc_2771;
wire uc_2772;
wire uc_2773;
wire uc_2774;
wire uc_2775;
wire uc_2776;
wire uc_2777;
wire uc_2778;
wire uc_2779;
wire uc_2780;
wire uc_2781;
wire uc_2782;
wire uc_2783;
wire uc_2784;
wire uc_2785;
wire uc_2786;
wire uc_2787;
wire uc_2788;
wire uc_2789;
wire uc_2790;
wire uc_2791;
wire uc_2792;
wire uc_2793;
wire uc_2794;
wire uc_2795;
wire uc_2796;
wire uc_2797;
wire uc_2798;
wire uc_2799;
wire uc_2800;
wire uc_2801;
wire uc_2802;
wire uc_2803;
wire uc_2804;
wire uc_2805;
wire uc_2806;
wire uc_2807;
wire uc_2808;
wire uc_2809;
wire uc_2810;
wire uc_2811;
wire uc_2812;
wire uc_2813;
wire uc_2814;
wire uc_2815;
wire uc_2816;
wire uc_2817;
wire uc_2818;
wire uc_2819;
wire uc_2820;
wire uc_2821;
wire uc_2822;
wire uc_2823;
wire uc_2824;
wire uc_2825;
wire uc_2826;
wire uc_2827;
wire uc_2828;
wire uc_2829;
wire uc_2830;
wire uc_2831;
wire uc_2832;
wire uc_2833;
wire uc_2834;
wire uc_2835;
wire uc_2836;
wire uc_2837;
wire uc_2838;
wire uc_2839;
wire uc_2840;
wire uc_2841;
wire uc_2842;
wire uc_2843;
wire uc_2844;
wire uc_2845;
wire uc_2846;
wire uc_2847;
wire uc_2848;
wire uc_2849;
wire uc_2850;
wire uc_2851;
wire uc_2852;
wire uc_2853;
wire uc_2854;
wire uc_2855;
wire uc_2856;
wire uc_2857;
wire uc_2858;
wire uc_2859;
wire uc_2860;
wire uc_2861;
wire uc_2862;
wire uc_2863;
wire uc_2864;
wire uc_2865;
wire uc_2866;
wire uc_2867;
wire uc_2868;
wire uc_2869;
wire uc_2870;
wire uc_2871;
wire uc_2872;
wire uc_2873;
wire uc_2874;
wire uc_2875;
wire uc_2876;
wire uc_2877;
wire uc_2878;
wire uc_2879;
wire uc_2880;
wire uc_2881;
wire uc_2882;
wire uc_2883;
wire uc_2884;
wire uc_2885;
wire uc_2886;
wire uc_2887;
wire uc_2888;
wire uc_2889;
wire uc_2890;
wire uc_2891;
wire uc_2892;
wire uc_2893;
wire uc_2894;
wire uc_2895;
wire uc_2896;
wire uc_2897;
wire uc_2898;
wire uc_2899;
wire uc_2900;
wire uc_2901;
wire uc_2902;
wire uc_2903;
wire uc_2904;
wire uc_2905;
wire uc_2906;
wire uc_2907;
wire uc_2908;
wire uc_2909;
wire uc_2910;
wire uc_2911;
wire uc_2912;
wire uc_2913;
wire uc_2914;
wire uc_2915;
wire uc_2916;
wire uc_2917;
wire uc_2918;
wire uc_2919;
wire uc_2920;
wire uc_2921;
wire uc_2922;
wire uc_2923;
wire uc_2924;
wire uc_2925;
wire uc_2926;
wire uc_2927;
wire uc_2928;
wire uc_2929;
wire uc_2930;
wire uc_2931;
wire uc_2932;
wire uc_2933;
wire uc_2934;
wire uc_2935;
wire uc_2936;
wire uc_2937;
wire uc_2938;
wire uc_2939;
wire uc_2940;
wire uc_2941;
wire uc_2942;
wire uc_2943;
wire uc_2944;
wire uc_2945;
wire uc_2946;
wire uc_2947;
wire uc_2948;
wire uc_2949;
wire uc_2950;
wire uc_2951;
wire uc_2952;
wire uc_2953;
wire uc_2954;
wire uc_2955;
wire uc_2956;
wire uc_2957;
wire uc_2958;
wire uc_2959;
wire uc_2960;
wire uc_2961;
wire uc_2962;
wire uc_2963;
wire uc_2964;
wire uc_2965;
wire uc_2966;
wire uc_2967;
wire uc_2968;
wire uc_2969;
wire uc_2970;
wire uc_2971;
wire uc_2972;
wire uc_2973;
wire uc_2974;
wire uc_2975;
wire uc_2976;
wire uc_2977;
wire uc_2978;
wire uc_2979;
wire uc_2980;
wire uc_2981;
wire uc_2982;
wire uc_2983;
wire uc_2984;
wire uc_2985;
wire uc_2986;
wire uc_2987;
wire uc_2988;
wire uc_2989;
wire uc_2990;
wire uc_2991;
wire uc_2992;
wire uc_2993;
wire uc_2994;
wire uc_2995;
wire uc_2996;
wire uc_2997;
wire uc_2998;
wire uc_2999;
wire uc_3000;
wire uc_3001;
wire uc_3002;
wire uc_3003;
wire uc_3004;
wire uc_3005;
wire uc_3006;
wire uc_3007;
wire uc_3008;
wire uc_3009;
wire uc_3010;
wire uc_3011;
wire uc_3012;
wire uc_3013;
wire uc_3014;
wire uc_3015;
wire uc_3016;
wire uc_3017;
wire uc_3018;
wire uc_3019;
wire uc_3020;
wire uc_3021;
wire uc_3022;
wire uc_3023;
wire uc_3024;
wire uc_3025;
wire uc_3026;
wire uc_3027;
wire uc_3028;
wire uc_3029;
wire uc_3030;
wire uc_3031;
wire uc_3032;
wire uc_3033;
wire uc_3034;
wire uc_3035;
wire uc_3036;
wire uc_3037;
wire uc_3038;
wire uc_3039;
wire uc_3040;
wire uc_3041;
wire uc_3042;
wire uc_3043;
wire uc_3044;
wire uc_3045;
wire uc_3046;
wire uc_3047;
wire uc_3048;
wire uc_3049;
wire uc_3050;
wire uc_3051;
wire uc_3052;
wire uc_3053;
wire uc_3054;
wire uc_3055;
wire uc_3056;
wire uc_3057;
wire uc_3058;
wire uc_3059;
wire uc_3060;
wire uc_3061;
wire uc_3062;
wire uc_3063;
wire uc_3064;
wire uc_3065;
wire uc_3066;
wire uc_3067;
wire uc_3068;
wire uc_3069;
wire uc_3070;
wire uc_3071;
wire uc_3072;
wire uc_3073;
wire uc_3074;
wire uc_3075;
wire uc_3076;
wire uc_3077;
wire uc_3078;
wire uc_3079;
wire uc_3080;
wire uc_3081;
wire uc_3082;
wire uc_3083;
wire uc_3084;
wire uc_3085;
wire uc_3086;
wire uc_3087;
wire uc_3088;
wire uc_3089;
wire uc_3090;
wire uc_3091;
wire uc_3092;
wire uc_3093;
wire uc_3094;
wire uc_3095;
wire uc_3096;
wire uc_3097;
wire uc_3098;
wire uc_3099;
wire uc_3100;
wire uc_3101;
wire uc_3102;
wire uc_3103;
wire uc_3104;
wire uc_3105;
wire uc_3106;
wire uc_3107;
wire uc_3108;
wire uc_3109;
wire uc_3110;
wire uc_3111;
wire uc_3112;
wire uc_3113;
wire uc_3114;
wire uc_3115;
wire uc_3116;
wire uc_3117;
wire uc_3118;
wire uc_3119;
wire uc_3120;
wire uc_3121;
wire uc_3122;
wire uc_3123;
wire uc_3124;
wire uc_3125;
wire uc_3126;
wire uc_3127;
wire uc_3128;
wire uc_3129;
wire uc_3130;
wire uc_3131;
wire uc_3132;
wire uc_3133;
wire uc_3134;
wire uc_3135;
wire uc_3136;
wire uc_3137;
wire uc_3138;
wire uc_3139;
wire uc_3140;
wire uc_3141;
wire uc_3142;
wire uc_3143;
wire uc_3144;
wire uc_3145;
wire uc_3146;
wire uc_3147;
wire uc_3148;
wire uc_3149;
wire uc_3150;
wire uc_3151;
wire uc_3152;
wire uc_3153;
wire uc_3154;
wire uc_3155;
wire uc_3156;
wire uc_3157;
wire uc_3158;
wire uc_3159;
wire uc_3160;
wire uc_3161;
wire uc_3162;
wire uc_3163;
wire uc_3164;
wire uc_3165;
wire uc_3166;
wire uc_3167;
wire uc_3168;
wire uc_3169;
wire uc_3170;
wire uc_3171;
wire uc_3172;
wire uc_3173;
wire uc_3174;
wire uc_3175;
wire uc_3176;
wire uc_3177;
wire uc_3178;
wire uc_3179;
wire uc_3180;
wire uc_3181;
wire uc_3182;
wire uc_3183;
wire uc_3184;
wire uc_3185;
wire uc_3186;
wire uc_3187;
wire uc_3188;
wire uc_3189;
wire uc_3190;
wire uc_3191;
wire uc_3192;
wire uc_3193;
wire uc_3194;
wire uc_3195;
wire uc_3196;
wire uc_3197;
wire uc_3198;
wire uc_3199;
wire uc_3200;
wire uc_3201;
wire uc_3202;
wire uc_3203;
wire uc_3204;
wire uc_3205;
wire uc_3206;
wire uc_3207;
wire uc_3208;
wire uc_3209;
wire uc_3210;
wire uc_3211;
wire uc_3212;
wire uc_3213;
wire uc_3214;
wire uc_3215;
wire uc_3216;
wire uc_3217;
wire uc_3218;
wire uc_3219;
wire uc_3220;
wire uc_3221;
wire uc_3222;
wire uc_3223;
wire uc_3224;
wire uc_3225;
wire uc_3226;
wire uc_3227;
wire uc_3228;
wire uc_3229;
wire uc_3230;
wire uc_3231;
wire uc_3232;
wire uc_3233;
wire uc_3234;
wire uc_3235;
wire uc_3236;
wire uc_3237;
wire uc_3238;
wire uc_3239;
wire uc_3240;
wire uc_3241;
wire uc_3242;
wire uc_3243;
wire uc_3244;
wire uc_3245;
wire uc_3246;
wire uc_3247;
wire uc_3248;
wire uc_3249;
wire uc_3250;
wire uc_3251;
wire uc_3252;
wire uc_3253;
wire uc_3254;
wire uc_3255;
wire uc_3256;
wire uc_3257;
wire uc_3258;
wire uc_3259;
wire uc_3260;
wire uc_3261;
wire uc_3262;
wire uc_3263;
wire uc_3264;
wire uc_3265;
wire uc_3266;
wire uc_3267;
wire uc_3268;
wire uc_3269;
wire uc_3270;
wire uc_3271;
wire uc_3272;
wire uc_3273;
wire uc_3274;
wire uc_3275;
wire uc_3276;
wire uc_3277;
wire uc_3278;
wire uc_3279;
wire uc_3280;
wire uc_3281;
wire uc_3282;
wire uc_3283;
wire uc_3284;
wire uc_3285;
wire uc_3286;
wire uc_3287;
wire uc_3288;
wire uc_3289;
wire uc_3290;
wire uc_3291;
wire uc_3292;
wire uc_3293;
wire uc_3294;
wire uc_3295;
wire uc_3296;
wire uc_3297;
wire uc_3298;
wire uc_3299;
wire uc_3300;
wire uc_3301;
wire uc_3302;
wire uc_3303;
wire uc_3304;
wire uc_3305;
wire uc_3306;
wire uc_3307;
wire uc_3308;
wire uc_3309;
wire uc_3310;
wire uc_3311;
wire uc_3312;
wire uc_3313;
wire uc_3314;
wire uc_3315;
wire uc_3316;
wire uc_3317;
wire uc_3318;
wire uc_3319;
wire uc_3320;
wire uc_3321;
wire uc_3322;
wire uc_3323;
wire uc_3324;
wire uc_3325;
wire uc_3326;
wire uc_3327;
wire uc_3328;
wire uc_3329;
wire uc_3330;
wire uc_3331;
wire uc_3332;
wire uc_3333;
wire uc_3334;
wire uc_3335;
wire uc_3336;
wire uc_3337;
wire uc_3338;
wire uc_3339;
wire uc_3340;
wire uc_3341;
wire uc_3342;
wire uc_3343;
wire uc_3344;
wire uc_3345;
wire uc_3346;
wire uc_3347;
wire uc_3348;
wire uc_3349;
wire uc_3350;
wire uc_3351;
wire uc_3352;
wire uc_3353;
wire uc_3354;
wire uc_3355;
wire uc_3356;
wire uc_3357;
wire uc_3358;
wire uc_3359;
wire uc_3360;
wire uc_3361;
wire uc_3362;
wire uc_3363;
wire uc_3364;
wire uc_3365;
wire uc_3366;
wire uc_3367;
wire uc_3368;
wire uc_3369;
wire uc_3370;
wire uc_3371;
wire uc_3372;
wire uc_3373;
wire uc_3374;
wire uc_3375;
wire uc_3376;
wire uc_3377;
wire uc_3378;
wire uc_3379;
wire uc_3380;
wire uc_3381;
wire uc_3382;
wire uc_3383;
wire uc_3384;
wire uc_3385;
wire uc_3386;
wire uc_3387;
wire uc_3388;
wire uc_3389;
wire uc_3390;
wire uc_3391;
wire uc_3392;
wire uc_3393;
wire uc_3394;
wire uc_3395;
wire uc_3396;
wire uc_3397;
wire uc_3398;
wire uc_3399;
wire uc_3400;
wire uc_3401;
wire uc_3402;
wire uc_3403;
wire uc_3404;
wire uc_3405;
wire uc_3406;
wire uc_3407;
wire uc_3408;
wire uc_3409;
wire uc_3410;
wire uc_3411;
wire uc_3412;
wire uc_3413;
wire uc_3414;
wire uc_3415;
wire uc_3416;
wire uc_3417;
wire uc_3418;
wire uc_3419;
wire uc_3420;
wire uc_3421;
wire uc_3422;
wire uc_3423;
wire uc_3424;
wire uc_3425;
wire uc_3426;
wire uc_3427;
wire uc_3428;
wire uc_3429;
wire uc_3430;
wire uc_3431;
wire uc_3432;
wire uc_3433;
wire uc_3434;
wire uc_3435;
wire uc_3436;
wire uc_3437;
wire uc_3438;
wire uc_3439;
wire uc_3440;
wire uc_3441;
wire uc_3442;
wire uc_3443;
wire uc_3444;
wire uc_3445;
wire uc_3446;
wire uc_3447;
wire uc_3448;
wire uc_3449;
wire uc_3450;
wire uc_3451;
wire uc_3452;
wire uc_3453;
wire uc_3454;
wire uc_3455;
wire uc_3456;
wire uc_3457;
wire uc_3458;
wire uc_3459;
wire uc_3460;
wire uc_3461;
wire uc_3462;
wire uc_3463;
wire uc_3464;
wire uc_3465;
wire uc_3466;
wire uc_3467;
wire uc_3468;
wire uc_3469;
wire uc_3470;
wire uc_3471;
wire uc_3472;
wire uc_3473;
wire uc_3474;
wire uc_3475;
wire uc_3476;
wire uc_3477;
wire uc_3478;
wire uc_3479;
wire uc_3480;
wire uc_3481;
wire uc_3482;
wire uc_3483;
wire uc_3484;
wire uc_3485;
wire uc_3486;
wire uc_3487;
wire uc_3488;
wire uc_3489;
wire uc_3490;
wire uc_3491;
wire uc_3492;
wire uc_3493;
wire uc_3494;
wire uc_3495;
wire uc_3496;
wire uc_3497;
wire uc_3498;
wire uc_3499;
wire uc_3500;
wire uc_3501;
wire uc_3502;
wire uc_3503;
wire uc_3504;
wire uc_3505;
wire uc_3506;
wire uc_3507;
wire uc_3508;
wire uc_3509;
wire uc_3510;
wire uc_3511;
wire uc_3512;
wire uc_3513;
wire uc_3514;
wire uc_3515;
wire uc_3516;
wire uc_3517;
wire uc_3518;
wire uc_3519;
wire uc_3520;
wire uc_3521;
wire uc_3522;
wire uc_3523;
wire uc_3524;
wire uc_3525;
wire uc_3526;
wire uc_3527;
wire uc_3528;
wire uc_3529;
wire uc_3530;
wire uc_3531;
wire uc_3532;
wire uc_3533;
wire uc_3534;
wire uc_3535;
wire uc_3536;
wire uc_3537;
wire uc_3538;
wire uc_3539;
wire uc_3540;
wire uc_3541;
wire uc_3542;
wire uc_3543;
wire uc_3544;
wire uc_3545;
wire uc_3546;
wire uc_3547;
wire uc_3548;
wire uc_3549;
wire uc_3550;
wire uc_3551;
wire uc_3552;
wire uc_3553;
wire uc_3554;
wire uc_3555;
wire uc_3556;
wire uc_3557;
wire uc_3558;
wire uc_3559;
wire uc_3560;
wire uc_3561;
wire uc_3562;
wire uc_3563;
wire uc_3564;
wire uc_3565;
wire uc_3566;
wire uc_3567;
wire uc_3568;
wire uc_3569;
wire uc_3570;
wire uc_3571;
wire uc_3572;
wire uc_3573;
wire uc_3574;
wire uc_3575;
wire uc_3576;
wire uc_3577;
wire uc_3578;
wire uc_3579;
wire uc_3580;
wire uc_3581;
wire uc_3582;
wire uc_3583;
wire uc_3584;
wire uc_3585;
wire uc_3586;
wire uc_3587;
wire uc_3588;
wire uc_3589;
wire uc_3590;
wire uc_3591;
wire uc_3592;
wire uc_3593;
wire uc_3594;
wire uc_3595;
wire uc_3596;
wire uc_3597;
wire uc_3598;
wire uc_3599;
wire uc_3600;
wire uc_3601;
wire uc_3602;
wire uc_3603;
wire uc_3604;
wire uc_3605;
wire uc_3606;
wire uc_3607;
wire uc_3608;
wire uc_3609;
wire uc_3610;
wire uc_3611;
wire uc_3612;
wire uc_3613;
wire uc_3614;
wire uc_3615;
wire uc_3616;
wire uc_3617;
wire uc_3618;
wire uc_3619;
wire uc_3620;
wire uc_3621;
wire uc_3622;
wire uc_3623;
wire uc_3624;
wire uc_3625;
wire uc_3626;
wire uc_3627;
wire uc_3628;
wire uc_3629;
wire uc_3630;
wire uc_3631;
wire uc_3632;
wire uc_3633;
wire uc_3634;
wire uc_3635;
wire uc_3636;
wire uc_3637;
wire uc_3638;
wire uc_3639;
wire uc_3640;
wire uc_3641;
wire uc_3642;
wire uc_3643;
wire uc_3644;
wire uc_3645;
wire uc_3646;
wire uc_3647;
wire uc_3648;
wire uc_3649;
wire uc_3650;
wire uc_3651;
wire uc_3652;
wire uc_3653;
wire uc_3654;
wire uc_3655;
wire uc_3656;
wire uc_3657;
wire uc_3658;
wire uc_3659;
wire uc_3660;
wire uc_3661;
wire uc_3662;
wire uc_3663;
wire uc_3664;
wire uc_3665;
wire uc_3666;
wire uc_3667;
wire uc_3668;
wire uc_3669;
wire uc_3670;
wire uc_3671;
wire uc_3672;
wire uc_3673;
wire uc_3674;
wire uc_3675;
wire uc_3676;
wire uc_3677;
wire uc_3678;
wire uc_3679;
wire uc_3680;
wire uc_3681;
wire uc_3682;
wire uc_3683;
wire uc_3684;
wire uc_3685;
wire uc_3686;
wire uc_3687;
wire uc_3688;
wire uc_3689;
wire uc_3690;
wire uc_3691;
wire uc_3692;
wire uc_3693;
wire uc_3694;
wire uc_3695;
wire uc_3696;
wire uc_3697;
wire uc_3698;
wire uc_3699;
wire uc_3700;
wire uc_3701;
wire uc_3702;
wire uc_3703;
wire uc_3704;
wire uc_3705;
wire uc_3706;
wire uc_3707;
wire uc_3708;
wire uc_3709;
wire uc_3710;
wire uc_3711;
wire uc_3712;
wire uc_3713;
wire uc_3714;
wire uc_3715;
wire uc_3716;
wire uc_3717;
wire uc_3718;
wire uc_3719;
wire uc_3720;
wire uc_3721;
wire uc_3722;
wire uc_3723;
wire uc_3724;
wire uc_3725;
wire uc_3726;
wire uc_3727;
wire uc_3728;
wire uc_3729;
wire uc_3730;
wire uc_3731;
wire uc_3732;
wire uc_3733;
wire uc_3734;
wire uc_3735;
wire uc_3736;
wire uc_3737;
wire uc_3738;
wire uc_3739;
wire uc_3740;
wire uc_3741;
wire uc_3742;
wire uc_3743;
wire uc_3744;
wire uc_3745;
wire uc_3746;
wire uc_3747;
wire uc_3748;
wire uc_3749;
wire uc_3750;
wire uc_3751;
wire uc_3752;
wire uc_3753;
wire uc_3754;
wire uc_3755;
wire uc_3756;
wire uc_3757;
wire uc_3758;
wire uc_3759;
wire uc_3760;
wire uc_3761;
wire uc_3762;
wire uc_3763;
wire uc_3764;
wire uc_3765;
wire uc_3766;
wire uc_3767;
wire uc_3768;
wire uc_3769;
wire uc_3770;
wire uc_3771;
wire uc_3772;
wire uc_3773;
wire uc_3774;
wire uc_3775;
wire uc_3776;
wire uc_3777;
wire uc_3778;
wire uc_3779;
wire uc_3780;
wire uc_3781;
wire uc_3782;
wire uc_3783;
wire uc_3784;
wire uc_3785;
wire uc_3786;
wire uc_3787;
wire uc_3788;
wire uc_3789;
wire uc_3790;
wire uc_3791;
wire uc_3792;
wire uc_3793;
wire uc_3794;
wire uc_3795;
wire uc_3796;
wire uc_3797;
wire uc_3798;
wire uc_3799;
wire uc_3800;
wire uc_3801;
wire uc_3802;
wire uc_3803;
wire uc_3804;
wire uc_3805;
wire uc_3806;
wire uc_3807;
wire uc_3808;
wire uc_3809;
wire uc_3810;
wire uc_3811;
wire uc_3812;
wire uc_3813;
wire uc_3814;
wire uc_3815;
wire uc_3816;
wire uc_3817;
wire uc_3818;
wire uc_3819;
wire uc_3820;
wire uc_3821;
wire uc_3822;
wire uc_3823;
wire uc_3824;
wire uc_3825;
wire uc_3826;
wire uc_3827;
wire uc_3828;
wire uc_3829;
wire uc_3830;
wire uc_3831;
wire uc_3832;
wire uc_3833;
wire uc_3834;
wire uc_3835;
wire uc_3836;
wire uc_3837;
wire uc_3838;
wire uc_3839;
wire uc_3840;
wire uc_3841;
wire uc_3842;
wire uc_3843;
wire uc_3844;
wire uc_3845;
wire uc_3846;
wire uc_3847;
wire uc_3848;
wire uc_3849;
wire uc_3850;
wire uc_3851;
wire uc_3852;
wire uc_3853;
wire uc_3854;
wire uc_3855;
wire uc_3856;
wire uc_3857;
wire uc_3858;
wire uc_3859;
wire uc_3860;
wire uc_3861;
wire uc_3862;
wire uc_3863;
wire uc_3864;
wire uc_3865;
wire uc_3866;
wire uc_3867;
wire uc_3868;
wire uc_3869;
wire uc_3870;
wire uc_3871;
wire uc_3872;
wire uc_3873;
wire uc_3874;
wire uc_3875;
wire uc_3876;
wire uc_3877;
wire uc_3878;
wire uc_3879;
wire uc_3880;
wire uc_3881;
wire uc_3882;
wire uc_3883;
wire uc_3884;
wire uc_3885;
wire uc_3886;
wire uc_3887;
wire uc_3888;
wire uc_3889;
wire uc_3890;
wire uc_3891;
wire uc_3892;
wire uc_3893;
wire uc_3894;
wire uc_3895;
wire uc_3896;
wire uc_3897;
wire uc_3898;
wire uc_3899;
wire uc_3900;
wire uc_3901;
wire uc_3902;
wire uc_3903;
wire uc_3904;
wire uc_3905;
wire uc_3906;
wire uc_3907;
wire uc_3908;
wire uc_3909;
wire uc_3910;
wire uc_3911;
wire uc_3912;
wire uc_3913;
wire uc_3914;
wire uc_3915;
wire uc_3916;
wire uc_3917;
wire uc_3918;
wire uc_3919;
wire uc_3920;
wire uc_3921;
wire uc_3922;
wire uc_3923;
wire uc_3924;
wire uc_3925;
wire uc_3926;
wire uc_3927;
wire uc_3928;
wire uc_3929;
wire uc_3930;
wire uc_3931;
wire uc_3932;
wire uc_3933;
wire uc_3934;
wire uc_3935;
wire uc_3936;
wire uc_3937;
wire uc_3938;
wire uc_3939;
wire uc_3940;
wire uc_3941;
wire uc_3942;
wire uc_3943;
wire uc_3944;
wire uc_3945;
wire uc_3946;
wire uc_3947;
wire uc_3948;
wire uc_3949;
wire uc_3950;
wire uc_3951;
wire uc_3952;
wire uc_3953;
wire uc_3954;
wire uc_3955;
wire uc_3956;
wire uc_3957;
wire uc_3958;
wire uc_3959;
wire uc_3960;
wire uc_3961;
wire uc_3962;
wire uc_3963;
wire uc_3964;
wire uc_3965;
wire uc_3966;
wire uc_3967;
wire uc_3968;
wire uc_3969;
wire uc_3970;
wire uc_3971;
wire uc_3972;
wire uc_3973;
wire uc_3974;
wire uc_3975;
wire uc_3976;
wire uc_3977;
wire uc_3978;
wire uc_3979;
wire uc_3980;
wire uc_3981;
wire uc_3982;
wire uc_3983;
wire uc_3984;
wire uc_3985;
wire uc_3986;
wire uc_3987;
wire uc_3988;
wire uc_3989;
wire uc_3990;
wire uc_3991;
wire uc_3992;
wire uc_3993;
wire uc_3994;
wire uc_3995;
wire uc_3996;
wire uc_3997;
wire uc_3998;
wire uc_3999;
wire uc_4000;
wire uc_4001;
wire uc_4002;
wire uc_4003;
wire uc_4004;
wire uc_4005;
wire uc_4006;
wire uc_4007;
wire uc_4008;
wire uc_4009;
wire uc_4010;
wire uc_4011;
wire uc_4012;
wire uc_4013;
wire uc_4014;
wire uc_4015;
wire uc_4016;
wire uc_4017;
wire uc_4018;
wire uc_4019;
wire uc_4020;
wire uc_4021;
wire uc_4022;
wire uc_4023;
wire uc_4024;
wire uc_4025;
wire uc_4026;
wire uc_4027;
wire uc_4028;
wire uc_4029;
wire uc_4030;
wire uc_4031;
wire uc_4032;
wire uc_4033;
wire uc_4034;
wire uc_4035;
wire uc_4036;
wire uc_4037;
wire uc_4038;
wire uc_4039;
wire uc_4040;
wire uc_4041;
wire uc_4042;
wire uc_4043;
wire uc_4044;
wire uc_4045;
wire uc_4046;
wire uc_4047;
wire uc_4048;
wire uc_4049;
wire uc_4050;
wire uc_4051;
wire uc_4052;
wire uc_4053;
wire uc_4054;
wire uc_4055;
wire uc_4056;
wire uc_4057;
wire uc_4058;
wire uc_4059;
wire uc_4060;
wire uc_4061;
wire uc_4062;
wire uc_4063;
wire uc_4064;
wire uc_4065;
wire uc_4066;
wire uc_4067;
wire uc_4068;
wire uc_4069;
wire uc_4070;
wire uc_4071;
wire uc_4072;
wire uc_4073;
wire uc_4074;
wire uc_4075;
wire uc_4076;
wire uc_4077;
wire uc_4078;
wire uc_4079;
wire uc_4080;
wire uc_4081;
wire uc_4082;
wire uc_4083;
wire uc_4084;
wire uc_4085;
wire uc_4086;
wire uc_4087;
wire uc_4088;
wire uc_4089;
wire uc_4090;
wire uc_4091;
wire uc_4092;
wire uc_4093;
wire uc_4094;
wire uc_4095;
wire uc_4096;
wire uc_4097;
wire uc_4098;
wire uc_4099;
wire uc_4100;
wire uc_4101;
wire uc_4102;
wire uc_4103;
wire uc_4104;
wire uc_4105;
wire uc_4106;
wire uc_4107;
wire uc_4108;
wire uc_4109;
wire uc_4110;
wire uc_4111;
wire uc_4112;
wire uc_4113;
wire uc_4114;
wire uc_4115;
wire uc_4116;
wire uc_4117;
wire uc_4118;
wire uc_4119;
wire uc_4120;
wire uc_4121;
wire uc_4122;
wire uc_4123;
wire uc_4124;
wire uc_4125;
wire uc_4126;
wire uc_4127;
wire uc_4128;
wire uc_4129;
wire uc_4130;
wire uc_4131;
wire uc_4132;
wire uc_4133;
wire uc_4134;
wire uc_4135;
wire uc_4136;
wire uc_4137;
wire uc_4138;
wire uc_4139;
wire uc_4140;
wire uc_4141;
wire uc_4142;
wire uc_4143;
wire uc_4144;
wire uc_4145;
wire uc_4146;
wire uc_4147;
wire uc_4148;
wire uc_4149;
wire uc_4150;
wire uc_4151;
wire uc_4152;
wire uc_4153;
wire uc_4154;
wire uc_4155;
wire uc_4156;
wire uc_4157;
wire uc_4158;
wire uc_4159;
wire uc_4160;
wire uc_4161;
wire uc_4162;
wire uc_4163;
wire uc_4164;
wire uc_4165;
wire uc_4166;
wire uc_4167;
wire uc_4168;
wire uc_4169;
wire uc_4170;
wire uc_4171;
wire uc_4172;
wire uc_4173;
wire uc_4174;
wire uc_4175;
wire uc_4176;
wire uc_4177;
wire uc_4178;
wire uc_4179;
wire uc_4180;
wire uc_4181;
wire uc_4182;
wire uc_4183;
wire uc_4184;
wire uc_4185;
wire uc_4186;
wire uc_4187;
wire uc_4188;
wire uc_4189;
wire uc_4190;
wire uc_4191;
wire uc_4192;
wire uc_4193;
wire uc_4194;
wire uc_4195;
wire uc_4196;
wire uc_4197;
wire uc_4198;
wire uc_4199;
wire uc_4200;
wire uc_4201;
wire uc_4202;
wire uc_4203;
wire uc_4204;
wire uc_4205;
wire uc_4206;
wire uc_4207;
wire uc_4208;
wire uc_4209;
wire uc_4210;
wire uc_4211;
wire uc_4212;
wire uc_4213;
wire uc_4214;
wire uc_4215;
wire uc_4216;
wire uc_4217;
wire uc_4218;
wire uc_4219;
wire uc_4220;
wire uc_4221;
wire uc_4222;
wire uc_4223;
wire uc_4224;
wire uc_4225;
wire uc_4226;
wire uc_4227;
wire uc_4228;
wire uc_4229;
wire uc_4230;
wire uc_4231;
wire uc_4232;
wire uc_4233;
wire uc_4234;
wire uc_4235;
wire uc_4236;
wire uc_4237;
wire uc_4238;
wire uc_4239;
wire uc_4240;
wire uc_4241;
wire uc_4242;
wire uc_4243;
wire uc_4244;
wire uc_4245;
wire uc_4246;
wire uc_4247;
wire uc_4248;
wire uc_4249;
wire uc_4250;
wire uc_4251;
wire uc_4252;
wire uc_4253;
wire uc_4254;
wire uc_4255;
wire uc_4256;
wire uc_4257;
wire uc_4258;
wire uc_4259;
wire uc_4260;
wire uc_4261;
wire uc_4262;
wire uc_4263;
wire uc_4264;
wire uc_4265;
wire uc_4266;
wire uc_4267;
wire uc_4268;
wire uc_4269;
wire uc_4270;
wire uc_4271;
wire uc_4272;
wire uc_4273;
wire uc_4274;
wire uc_4275;
wire uc_4276;
wire uc_4277;
wire uc_4278;
wire uc_4279;
wire uc_4280;
wire uc_4281;
wire uc_4282;
wire uc_4283;
wire uc_4284;
wire uc_4285;
wire uc_4286;
wire uc_4287;
wire uc_4288;
wire uc_4289;
wire uc_4290;
wire uc_4291;
wire uc_4292;
wire uc_4293;
wire uc_4294;
wire uc_4295;
wire uc_4296;
wire uc_4297;
wire uc_4298;
wire uc_4299;
wire uc_4300;
wire uc_4301;
wire uc_4302;
wire uc_4303;
wire uc_4304;
wire uc_4305;
wire uc_4306;
wire uc_4307;
wire uc_4308;
wire uc_4309;
wire uc_4310;
wire uc_4311;
wire uc_4312;
wire uc_4313;
wire uc_4314;
wire uc_4315;
wire uc_4316;
wire uc_4317;
wire uc_4318;
wire uc_4319;
wire uc_4320;
wire uc_4321;
wire uc_4322;
wire uc_4323;
wire uc_4324;
wire uc_4325;
wire uc_4326;
wire uc_4327;
wire uc_4328;
wire uc_4329;
wire uc_4330;
wire uc_4331;
wire uc_4332;
wire uc_4333;
wire uc_4334;
wire uc_4335;
wire uc_4336;
wire uc_4337;
wire uc_4338;
wire uc_4339;
wire uc_4340;
wire uc_4341;
wire uc_4342;
wire uc_4343;
wire uc_4344;
wire uc_4345;
wire uc_4346;
wire uc_4347;
wire uc_4348;
wire uc_4349;
wire uc_4350;
wire uc_4351;
wire uc_4352;
wire uc_4353;
wire uc_4354;
wire uc_4355;
wire uc_4356;
wire uc_4357;
wire uc_4358;
wire uc_4359;
wire uc_4360;
wire uc_4361;
wire uc_4362;
wire uc_4363;
wire uc_4364;
wire uc_4365;
wire uc_4366;
wire uc_4367;
wire uc_4368;
wire uc_4369;
wire uc_4370;
wire uc_4371;
wire uc_4372;
wire uc_4373;
wire uc_4374;
wire uc_4375;
wire uc_4376;
wire uc_4377;
wire uc_4378;
wire uc_4379;
wire uc_4380;
wire uc_4381;
wire uc_4382;
wire uc_4383;
wire uc_4384;
wire uc_4385;
wire uc_4386;
wire uc_4387;
wire uc_4388;
wire uc_4389;
wire uc_4390;
wire uc_4391;
wire uc_4392;
wire uc_4393;
wire uc_4394;
wire uc_4395;
wire uc_4396;
wire uc_4397;
wire uc_4398;
wire uc_4399;
wire uc_4400;
wire uc_4401;
wire uc_4402;
wire uc_4403;
wire uc_4404;
wire uc_4405;
wire uc_4406;
wire uc_4407;
wire uc_4408;
wire uc_4409;
wire uc_4410;
wire uc_4411;
wire uc_4412;
wire uc_4413;
wire uc_4414;
wire uc_4415;
wire uc_4416;
wire uc_4417;
wire uc_4418;
wire uc_4419;
wire uc_4420;
wire uc_4421;
wire uc_4422;
wire uc_4423;
wire uc_4424;
wire uc_4425;
wire uc_4426;
wire uc_4427;
wire uc_4428;
wire uc_4429;
wire uc_4430;
wire uc_4431;
wire uc_4432;
wire uc_4433;
wire uc_4434;
wire uc_4435;
wire uc_4436;
wire uc_4437;
wire uc_4438;
wire uc_4439;
wire uc_4440;
wire uc_4441;
wire uc_4442;
wire uc_4443;
wire uc_4444;
wire uc_4445;
wire uc_4446;
wire uc_4447;
wire uc_4448;
wire uc_4449;
wire uc_4450;
wire uc_4451;
wire uc_4452;
wire uc_4453;
wire uc_4454;
wire uc_4455;
wire uc_4456;
wire uc_4457;
wire uc_4458;
wire uc_4459;
wire uc_4460;
wire uc_4461;
wire uc_4462;
wire uc_4463;
wire uc_4464;
wire uc_4465;
wire uc_4466;
wire uc_4467;
wire uc_4468;
wire uc_4469;
wire uc_4470;
wire uc_4471;
wire uc_4472;
wire uc_4473;
wire uc_4474;
wire uc_4475;
wire uc_4476;
wire uc_4477;
wire uc_4478;
wire uc_4479;
wire uc_4480;
wire uc_4481;
wire uc_4482;
wire uc_4483;
wire uc_4484;
wire uc_4485;
wire uc_4486;
wire uc_4487;
wire uc_4488;
wire uc_4489;


CSAlike genblk9_0_finalStage (.carry ({uc_4429, carry[62], carry[61], carry[60], 
    carry[59], carry[58], carry[57], carry[56], carry[55], carry[54], carry[53], 
    carry[52], carry[51], carry[50], carry[49], carry[48], carry[47], carry[46], 
    carry[45], carry[44], carry[43], carry[42], carry[41], carry[40], carry[39], 
    carry[38], carry[37], carry[36], carry[35], carry[34], carry[33], carry[32], 
    carry[31], carry[30], carry[29], carry[28], carry[27], carry[26], carry[25], 
    carry[24], carry[23], carry[22], carry[21], carry[20], carry[19], carry[18], 
    carry[17], carry[16], carry[15], carry[14], carry[13], carry[12], carry[11], 
    carry[10], carry[9], uc_4430, uc_4431, uc_4432, uc_4433, uc_4434, uc_4435, uc_4436, 
    uc_4437, uc_4438}), .result ({uc_4419, uc_4420, Res[61], Res[60], Res[59], Res[58], 
    Res[57], Res[56], Res[55], Res[54], Res[53], Res[52], Res[51], Res[50], Res[49], 
    Res[48], Res[47], Res[46], Res[45], Res[44], Res[43], Res[42], Res[41], Res[40], 
    Res[39], Res[38], Res[37], Res[36], Res[35], Res[34], Res[33], Res[32], Res[31], 
    Res[30], Res[29], Res[28], Res[27], Res[26], Res[25], Res[24], Res[23], Res[22], 
    Res[21], Res[20], Res[19], Res[18], Res[17], Res[16], Res[15], Res[14], Res[13], 
    Res[12], Res[11], Res[10], Res[9], Res[8], uc_4421, uc_4422, uc_4423, uc_4424, 
    uc_4425, uc_4426, uc_4427, uc_4428}), .A ({1'b0 , uc_4439, normalizedWires[2045], 
    \intermediateWiresStage3[8][60] , \intermediateWiresStage7[0][59] , \intermediateWiresStage7[0][58] , 
    \intermediateWiresStage7[0][57] , \intermediateWiresStage7[0][56] , \intermediateWiresStage7[0][55] , 
    \intermediateWiresStage7[0][54] , \intermediateWiresStage7[0][53] , \intermediateWiresStage7[0][52] , 
    \intermediateWiresStage7[0][51] , \intermediateWiresStage7[0][50] , \intermediateWiresStage7[0][49] , 
    \intermediateWiresStage7[0][48] , \intermediateWiresStage7[0][47] , \intermediateWiresStage7[0][46] , 
    \intermediateWiresStage7[0][45] , \intermediateWiresStage7[0][44] , \intermediateWiresStage7[0][43] , 
    \intermediateWiresStage7[0][42] , \intermediateWiresStage7[0][41] , \intermediateWiresStage7[0][40] , 
    \intermediateWiresStage7[0][39] , \intermediateWiresStage7[0][38] , \intermediateWiresStage7[0][37] , 
    \intermediateWiresStage7[0][36] , \intermediateWiresStage7[0][35] , \intermediateWiresStage7[0][34] , 
    \intermediateWiresStage7[0][33] , \intermediateWiresStage7[0][32] , \intermediateWiresStage7[0][31] , 
    \intermediateWiresStage7[0][30] , \intermediateWiresStage7[0][29] , \intermediateWiresStage7[0][28] , 
    \intermediateWiresStage7[0][27] , \intermediateWiresStage7[0][26] , \intermediateWiresStage7[0][25] , 
    \intermediateWiresStage7[0][24] , \intermediateWiresStage7[0][23] , \intermediateWiresStage7[0][22] , 
    \intermediateWiresStage7[0][21] , \intermediateWiresStage7[0][20] , \intermediateWiresStage7[0][19] , 
    \intermediateWiresStage7[0][18] , \intermediateWiresStage7[0][17] , \intermediateWiresStage7[0][16] , 
    \intermediateWiresStage7[0][15] , \intermediateWiresStage7[0][14] , \intermediateWiresStage7[0][13] , 
    \intermediateWiresStage7[0][12] , \intermediateWiresStage7[0][11] , \intermediateWiresStage7[0][10] , 
    \intermediateWiresStage7[0][9] , \intermediateWiresStage7[0][8] , uc_4440, uc_4441, 
    uc_4442, uc_4443, uc_4444, uc_4445, uc_4446, uc_4447}), .B ({1'b0 , uc_4448, 
    uc_4449, \intermediateWiresStage7[1][60] , \intermediateWiresStage7[1][59] , 
    \intermediateWiresStage7[1][58] , \intermediateWiresStage7[1][57] , \intermediateWiresStage7[1][56] , 
    \intermediateWiresStage7[1][55] , \intermediateWiresStage7[1][54] , \intermediateWiresStage7[1][53] , 
    \intermediateWiresStage7[1][52] , \intermediateWiresStage7[1][51] , \intermediateWiresStage7[1][50] , 
    \intermediateWiresStage7[1][49] , \intermediateWiresStage7[1][48] , \intermediateWiresStage7[1][47] , 
    \intermediateWiresStage7[1][46] , \intermediateWiresStage7[1][45] , \intermediateWiresStage7[1][44] , 
    \intermediateWiresStage7[1][43] , \intermediateWiresStage7[1][42] , \intermediateWiresStage7[1][41] , 
    \intermediateWiresStage7[1][40] , \intermediateWiresStage7[1][39] , \intermediateWiresStage7[1][38] , 
    \intermediateWiresStage7[1][37] , \intermediateWiresStage7[1][36] , \intermediateWiresStage7[1][35] , 
    \intermediateWiresStage7[1][34] , \intermediateWiresStage7[1][33] , \intermediateWiresStage7[1][32] , 
    \intermediateWiresStage7[1][31] , \intermediateWiresStage7[1][30] , \intermediateWiresStage7[1][29] , 
    \intermediateWiresStage7[1][28] , \intermediateWiresStage7[1][27] , \intermediateWiresStage7[1][26] , 
    \intermediateWiresStage7[1][25] , \intermediateWiresStage7[1][24] , \intermediateWiresStage7[1][23] , 
    \intermediateWiresStage7[1][22] , \intermediateWiresStage7[1][21] , \intermediateWiresStage7[1][20] , 
    \intermediateWiresStage7[1][19] , \intermediateWiresStage7[1][18] , \intermediateWiresStage7[1][17] , 
    \intermediateWiresStage7[1][16] , \intermediateWiresStage7[1][15] , \intermediateWiresStage7[1][14] , 
    \intermediateWiresStage7[1][13] , \intermediateWiresStage7[1][12] , \intermediateWiresStage7[1][11] , 
    \intermediateWiresStage7[1][10] , \intermediateWiresStage7[1][9] , \intermediateWiresStage7[1][8] , 
    uc_4450, uc_4451, uc_4452, uc_4453, uc_4454, uc_4455, uc_4456, uc_4457}), .C ({
    1'b0 , uc_4458, \intermediateWiresStage3[9][61] , \intermediateWiresStage3[9][60] , 
    \intermediateWiresStage3[9][59] , \intermediateWiresStage3[9][58] , \intermediateWiresStage3[9][57] , 
    \intermediateWiresStage3[9][56] , \intermediateWiresStage3[9][55] , \intermediateWiresStage3[9][54] , 
    \intermediateWiresStage3[9][53] , \intermediateWiresStage3[9][52] , \intermediateWiresStage3[9][51] , 
    \intermediateWiresStage3[9][50] , \intermediateWiresStage3[9][49] , \intermediateWiresStage3[9][48] , 
    \intermediateWiresStage3[9][47] , \intermediateWiresStage3[9][46] , \intermediateWiresStage3[9][45] , 
    \intermediateWiresStage3[9][44] , \intermediateWiresStage3[9][43] , \intermediateWiresStage3[9][42] , 
    \intermediateWiresStage3[9][41] , \intermediateWiresStage3[9][40] , \intermediateWiresStage3[9][39] , 
    \intermediateWiresStage3[9][38] , \intermediateWiresStage3[9][37] , \intermediateWiresStage3[9][36] , 
    \intermediateWiresStage3[9][35] , \intermediateWiresStage3[9][34] , \intermediateWiresStage3[9][33] , 
    \intermediateWiresStage3[9][32] , \intermediateWiresStage3[9][31] , uc_4459, 
    uc_4460, uc_4461, uc_4462, uc_4463, uc_4464, uc_4465, uc_4466, uc_4467, uc_4468, 
    uc_4469, uc_4470, uc_4471, uc_4472, uc_4473, uc_4474, uc_4475, uc_4476, uc_4477, 
    uc_4478, uc_4479, uc_4480, uc_4481, uc_4482, uc_4483, uc_4484, uc_4485, uc_4486, 
    uc_4487, uc_4488, uc_4489}));
CSAlike__4_2018 genblk8_0_parallelAdderStage7 (.carry ({uc_4358, uc_4359, uc_4360, 
    \intermediateWiresStage7[1][60] , \intermediateWiresStage7[1][59] , \intermediateWiresStage7[1][58] , 
    \intermediateWiresStage7[1][57] , \intermediateWiresStage7[1][56] , \intermediateWiresStage7[1][55] , 
    \intermediateWiresStage7[1][54] , \intermediateWiresStage7[1][53] , \intermediateWiresStage7[1][52] , 
    \intermediateWiresStage7[1][51] , \intermediateWiresStage7[1][50] , \intermediateWiresStage7[1][49] , 
    \intermediateWiresStage7[1][48] , \intermediateWiresStage7[1][47] , \intermediateWiresStage7[1][46] , 
    \intermediateWiresStage7[1][45] , \intermediateWiresStage7[1][44] , \intermediateWiresStage7[1][43] , 
    \intermediateWiresStage7[1][42] , \intermediateWiresStage7[1][41] , \intermediateWiresStage7[1][40] , 
    \intermediateWiresStage7[1][39] , \intermediateWiresStage7[1][38] , \intermediateWiresStage7[1][37] , 
    \intermediateWiresStage7[1][36] , \intermediateWiresStage7[1][35] , \intermediateWiresStage7[1][34] , 
    \intermediateWiresStage7[1][33] , \intermediateWiresStage7[1][32] , \intermediateWiresStage7[1][31] , 
    \intermediateWiresStage7[1][30] , \intermediateWiresStage7[1][29] , \intermediateWiresStage7[1][28] , 
    \intermediateWiresStage7[1][27] , \intermediateWiresStage7[1][26] , \intermediateWiresStage7[1][25] , 
    \intermediateWiresStage7[1][24] , \intermediateWiresStage7[1][23] , \intermediateWiresStage7[1][22] , 
    \intermediateWiresStage7[1][21] , \intermediateWiresStage7[1][20] , \intermediateWiresStage7[1][19] , 
    \intermediateWiresStage7[1][18] , \intermediateWiresStage7[1][17] , \intermediateWiresStage7[1][16] , 
    \intermediateWiresStage7[1][15] , \intermediateWiresStage7[1][14] , \intermediateWiresStage7[1][13] , 
    \intermediateWiresStage7[1][12] , \intermediateWiresStage7[1][11] , \intermediateWiresStage7[1][10] , 
    \intermediateWiresStage7[1][9] , \intermediateWiresStage7[1][8] , uc_4361, uc_4362, 
    uc_4363, uc_4364, uc_4365, uc_4366, uc_4367, uc_4368}), .result ({uc_4347, uc_4348, 
    uc_4349, uc_4350, \intermediateWiresStage7[0][59] , \intermediateWiresStage7[0][58] , 
    \intermediateWiresStage7[0][57] , \intermediateWiresStage7[0][56] , \intermediateWiresStage7[0][55] , 
    \intermediateWiresStage7[0][54] , \intermediateWiresStage7[0][53] , \intermediateWiresStage7[0][52] , 
    \intermediateWiresStage7[0][51] , \intermediateWiresStage7[0][50] , \intermediateWiresStage7[0][49] , 
    \intermediateWiresStage7[0][48] , \intermediateWiresStage7[0][47] , \intermediateWiresStage7[0][46] , 
    \intermediateWiresStage7[0][45] , \intermediateWiresStage7[0][44] , \intermediateWiresStage7[0][43] , 
    \intermediateWiresStage7[0][42] , \intermediateWiresStage7[0][41] , \intermediateWiresStage7[0][40] , 
    \intermediateWiresStage7[0][39] , \intermediateWiresStage7[0][38] , \intermediateWiresStage7[0][37] , 
    \intermediateWiresStage7[0][36] , \intermediateWiresStage7[0][35] , \intermediateWiresStage7[0][34] , 
    \intermediateWiresStage7[0][33] , \intermediateWiresStage7[0][32] , \intermediateWiresStage7[0][31] , 
    \intermediateWiresStage7[0][30] , \intermediateWiresStage7[0][29] , \intermediateWiresStage7[0][28] , 
    \intermediateWiresStage7[0][27] , \intermediateWiresStage7[0][26] , \intermediateWiresStage7[0][25] , 
    \intermediateWiresStage7[0][24] , \intermediateWiresStage7[0][23] , \intermediateWiresStage7[0][22] , 
    \intermediateWiresStage7[0][21] , \intermediateWiresStage7[0][20] , \intermediateWiresStage7[0][19] , 
    \intermediateWiresStage7[0][18] , \intermediateWiresStage7[0][17] , \intermediateWiresStage7[0][16] , 
    \intermediateWiresStage7[0][15] , \intermediateWiresStage7[0][14] , \intermediateWiresStage7[0][13] , 
    \intermediateWiresStage7[0][12] , \intermediateWiresStage7[0][11] , \intermediateWiresStage7[0][10] , 
    \intermediateWiresStage7[0][9] , \intermediateWiresStage7[0][8] , Res[7], uc_4351, 
    uc_4352, uc_4353, uc_4354, uc_4355, uc_4356, uc_4357}), .A ({1'b0 , uc_4369, 
    uc_4370, uc_4371, \intermediateWiresStage3[8][59] , \intermediateWiresStage5[2][58] , 
    \intermediateWiresStage5[2][57] , \intermediateWiresStage5[2][56] , \intermediateWiresStage5[2][55] , 
    \intermediateWiresStage5[2][54] , \intermediateWiresStage6[0][53] , \intermediateWiresStage6[0][52] , 
    \intermediateWiresStage6[0][51] , \intermediateWiresStage6[0][50] , \intermediateWiresStage6[0][49] , 
    \intermediateWiresStage6[0][48] , \intermediateWiresStage6[0][47] , \intermediateWiresStage6[0][46] , 
    \intermediateWiresStage6[0][45] , \intermediateWiresStage6[0][44] , \intermediateWiresStage6[0][43] , 
    \intermediateWiresStage6[0][42] , \intermediateWiresStage6[0][41] , \intermediateWiresStage6[0][40] , 
    \intermediateWiresStage6[0][39] , \intermediateWiresStage6[0][38] , \intermediateWiresStage6[0][37] , 
    \intermediateWiresStage6[0][36] , \intermediateWiresStage6[0][35] , \intermediateWiresStage6[0][34] , 
    \intermediateWiresStage6[0][33] , \intermediateWiresStage6[0][32] , \intermediateWiresStage6[0][31] , 
    \intermediateWiresStage6[0][30] , \intermediateWiresStage6[0][29] , \intermediateWiresStage6[0][28] , 
    \intermediateWiresStage6[0][27] , \intermediateWiresStage6[0][26] , \intermediateWiresStage6[0][25] , 
    \intermediateWiresStage6[0][24] , \intermediateWiresStage6[0][23] , \intermediateWiresStage6[0][22] , 
    \intermediateWiresStage6[0][21] , \intermediateWiresStage6[0][20] , \intermediateWiresStage6[0][19] , 
    \intermediateWiresStage6[0][18] , \intermediateWiresStage6[0][17] , \intermediateWiresStage6[0][16] , 
    \intermediateWiresStage6[0][15] , \intermediateWiresStage6[0][14] , \intermediateWiresStage6[0][13] , 
    \intermediateWiresStage6[0][12] , \intermediateWiresStage6[0][11] , \intermediateWiresStage6[0][10] , 
    \intermediateWiresStage6[0][9] , \intermediateWiresStage6[0][8] , \intermediateWiresStage6[0][7] , 
    uc_4372, uc_4373, uc_4374, uc_4375, uc_4376, uc_4377, uc_4378}), .B ({1'b0 , 
    uc_4379, uc_4380, uc_4381, uc_4382, uc_4383, uc_4384, uc_4385, uc_4386, \intermediateWiresStage6[1][54] , 
    \intermediateWiresStage6[1][53] , \intermediateWiresStage6[1][52] , \intermediateWiresStage6[1][51] , 
    \intermediateWiresStage6[1][50] , \intermediateWiresStage6[1][49] , \intermediateWiresStage6[1][48] , 
    \intermediateWiresStage6[1][47] , \intermediateWiresStage6[1][46] , \intermediateWiresStage6[1][45] , 
    \intermediateWiresStage6[1][44] , \intermediateWiresStage6[1][43] , \intermediateWiresStage6[1][42] , 
    \intermediateWiresStage6[1][41] , \intermediateWiresStage6[1][40] , \intermediateWiresStage6[1][39] , 
    \intermediateWiresStage6[1][38] , \intermediateWiresStage6[1][37] , \intermediateWiresStage6[1][36] , 
    \intermediateWiresStage6[1][35] , \intermediateWiresStage6[1][34] , \intermediateWiresStage6[1][33] , 
    \intermediateWiresStage6[1][32] , \intermediateWiresStage6[1][31] , \intermediateWiresStage6[1][30] , 
    \intermediateWiresStage6[1][29] , \intermediateWiresStage6[1][28] , \intermediateWiresStage6[1][27] , 
    \intermediateWiresStage6[1][26] , \intermediateWiresStage6[1][25] , \intermediateWiresStage6[1][24] , 
    \intermediateWiresStage6[1][23] , \intermediateWiresStage6[1][22] , \intermediateWiresStage6[1][21] , 
    \intermediateWiresStage6[1][20] , \intermediateWiresStage6[1][19] , \intermediateWiresStage6[1][18] , 
    \intermediateWiresStage6[1][17] , \intermediateWiresStage6[1][16] , \intermediateWiresStage6[1][15] , 
    \intermediateWiresStage6[1][14] , \intermediateWiresStage6[1][13] , \intermediateWiresStage6[1][12] , 
    \intermediateWiresStage6[1][11] , \intermediateWiresStage6[1][10] , \intermediateWiresStage6[1][9] , 
    \intermediateWiresStage6[1][8] , \intermediateWiresStage6[1][7] , uc_4387, uc_4388, 
    uc_4389, uc_4390, uc_4391, uc_4392, uc_4393}), .C ({1'b0 , uc_4394, uc_4395, 
    uc_4396, \intermediateWiresStage5[3][59] , \intermediateWiresStage5[3][58] , 
    \intermediateWiresStage5[3][57] , \intermediateWiresStage5[3][56] , \intermediateWiresStage5[3][55] , 
    \intermediateWiresStage5[3][54] , \intermediateWiresStage5[3][53] , \intermediateWiresStage5[3][52] , 
    \intermediateWiresStage5[3][51] , \intermediateWiresStage5[3][50] , \intermediateWiresStage5[3][49] , 
    \intermediateWiresStage5[3][48] , \intermediateWiresStage5[3][47] , \intermediateWiresStage5[3][46] , 
    \intermediateWiresStage5[3][45] , \intermediateWiresStage5[3][44] , \intermediateWiresStage5[3][43] , 
    \intermediateWiresStage5[3][42] , \intermediateWiresStage5[3][41] , \intermediateWiresStage5[3][40] , 
    \intermediateWiresStage5[3][39] , \intermediateWiresStage5[3][38] , \intermediateWiresStage5[3][37] , 
    \intermediateWiresStage5[3][36] , \intermediateWiresStage5[3][35] , \intermediateWiresStage5[3][34] , 
    \intermediateWiresStage5[3][33] , \intermediateWiresStage5[3][32] , \intermediateWiresStage5[3][31] , 
    \intermediateWiresStage5[3][30] , \intermediateWiresStage5[3][29] , \intermediateWiresStage5[3][28] , 
    \intermediateWiresStage5[3][27] , \intermediateWiresStage5[3][26] , \intermediateWiresStage5[3][25] , 
    \intermediateWiresStage5[3][24] , \intermediateWiresStage5[3][23] , \intermediateWiresStage5[3][22] , 
    uc_4397, uc_4398, uc_4399, uc_4400, uc_4401, uc_4402, uc_4403, uc_4404, uc_4405, 
    uc_4406, uc_4407, uc_4408, uc_4409, uc_4410, uc_4411, uc_4412, uc_4413, uc_4414, 
    uc_4415, uc_4416, uc_4417, uc_4418}));
CSAlike__4_1765 genblk7_0_parallelAdderStage6 (.carry ({uc_4269, uc_4270, uc_4271, 
    uc_4272, uc_4273, uc_4274, uc_4275, uc_4276, uc_4277, \intermediateWiresStage6[1][54] , 
    \intermediateWiresStage6[1][53] , \intermediateWiresStage6[1][52] , \intermediateWiresStage6[1][51] , 
    \intermediateWiresStage6[1][50] , \intermediateWiresStage6[1][49] , \intermediateWiresStage6[1][48] , 
    \intermediateWiresStage6[1][47] , \intermediateWiresStage6[1][46] , \intermediateWiresStage6[1][45] , 
    \intermediateWiresStage6[1][44] , \intermediateWiresStage6[1][43] , \intermediateWiresStage6[1][42] , 
    \intermediateWiresStage6[1][41] , \intermediateWiresStage6[1][40] , \intermediateWiresStage6[1][39] , 
    \intermediateWiresStage6[1][38] , \intermediateWiresStage6[1][37] , \intermediateWiresStage6[1][36] , 
    \intermediateWiresStage6[1][35] , \intermediateWiresStage6[1][34] , \intermediateWiresStage6[1][33] , 
    \intermediateWiresStage6[1][32] , \intermediateWiresStage6[1][31] , \intermediateWiresStage6[1][30] , 
    \intermediateWiresStage6[1][29] , \intermediateWiresStage6[1][28] , \intermediateWiresStage6[1][27] , 
    \intermediateWiresStage6[1][26] , \intermediateWiresStage6[1][25] , \intermediateWiresStage6[1][24] , 
    \intermediateWiresStage6[1][23] , \intermediateWiresStage6[1][22] , \intermediateWiresStage6[1][21] , 
    \intermediateWiresStage6[1][20] , \intermediateWiresStage6[1][19] , \intermediateWiresStage6[1][18] , 
    \intermediateWiresStage6[1][17] , \intermediateWiresStage6[1][16] , \intermediateWiresStage6[1][15] , 
    \intermediateWiresStage6[1][14] , \intermediateWiresStage6[1][13] , \intermediateWiresStage6[1][12] , 
    \intermediateWiresStage6[1][11] , \intermediateWiresStage6[1][10] , \intermediateWiresStage6[1][9] , 
    \intermediateWiresStage6[1][8] , \intermediateWiresStage6[1][7] , uc_4278, uc_4279, 
    uc_4280, uc_4281, uc_4282, uc_4283, uc_4284}), .result ({uc_4253, uc_4254, uc_4255, 
    uc_4256, uc_4257, uc_4258, uc_4259, uc_4260, uc_4261, uc_4262, \intermediateWiresStage6[0][53] , 
    \intermediateWiresStage6[0][52] , \intermediateWiresStage6[0][51] , \intermediateWiresStage6[0][50] , 
    \intermediateWiresStage6[0][49] , \intermediateWiresStage6[0][48] , \intermediateWiresStage6[0][47] , 
    \intermediateWiresStage6[0][46] , \intermediateWiresStage6[0][45] , \intermediateWiresStage6[0][44] , 
    \intermediateWiresStage6[0][43] , \intermediateWiresStage6[0][42] , \intermediateWiresStage6[0][41] , 
    \intermediateWiresStage6[0][40] , \intermediateWiresStage6[0][39] , \intermediateWiresStage6[0][38] , 
    \intermediateWiresStage6[0][37] , \intermediateWiresStage6[0][36] , \intermediateWiresStage6[0][35] , 
    \intermediateWiresStage6[0][34] , \intermediateWiresStage6[0][33] , \intermediateWiresStage6[0][32] , 
    \intermediateWiresStage6[0][31] , \intermediateWiresStage6[0][30] , \intermediateWiresStage6[0][29] , 
    \intermediateWiresStage6[0][28] , \intermediateWiresStage6[0][27] , \intermediateWiresStage6[0][26] , 
    \intermediateWiresStage6[0][25] , \intermediateWiresStage6[0][24] , \intermediateWiresStage6[0][23] , 
    \intermediateWiresStage6[0][22] , \intermediateWiresStage6[0][21] , \intermediateWiresStage6[0][20] , 
    \intermediateWiresStage6[0][19] , \intermediateWiresStage6[0][18] , \intermediateWiresStage6[0][17] , 
    \intermediateWiresStage6[0][16] , \intermediateWiresStage6[0][15] , \intermediateWiresStage6[0][14] , 
    \intermediateWiresStage6[0][13] , \intermediateWiresStage6[0][12] , \intermediateWiresStage6[0][11] , 
    \intermediateWiresStage6[0][10] , \intermediateWiresStage6[0][9] , \intermediateWiresStage6[0][8] , 
    \intermediateWiresStage6[0][7] , Res[6], uc_4263, uc_4264, uc_4265, uc_4266, 
    uc_4267, uc_4268}), .A ({1'b0 , uc_4285, uc_4286, uc_4287, uc_4288, uc_4289, 
    uc_4290, uc_4291, uc_4292, uc_4293, normalizedWires[1525], \intermediateWiresStage1[14][52] , 
    \intermediateWiresStage1[14][51] , \intermediateWiresStage2[8][50] , \intermediateWiresStage4[2][49] , 
    \intermediateWiresStage4[2][48] , \intermediateWiresStage4[2][47] , \intermediateWiresStage4[2][46] , 
    \intermediateWiresStage4[2][45] , \intermediateWiresStage5[0][44] , \intermediateWiresStage5[0][43] , 
    \intermediateWiresStage5[0][42] , \intermediateWiresStage5[0][41] , \intermediateWiresStage5[0][40] , 
    \intermediateWiresStage5[0][39] , \intermediateWiresStage5[0][38] , \intermediateWiresStage5[0][37] , 
    \intermediateWiresStage5[0][36] , \intermediateWiresStage5[0][35] , \intermediateWiresStage5[0][34] , 
    \intermediateWiresStage5[0][33] , \intermediateWiresStage5[0][32] , \intermediateWiresStage5[0][31] , 
    \intermediateWiresStage5[0][30] , \intermediateWiresStage5[0][29] , \intermediateWiresStage5[0][28] , 
    \intermediateWiresStage5[0][27] , \intermediateWiresStage5[0][26] , \intermediateWiresStage5[0][25] , 
    \intermediateWiresStage5[0][24] , \intermediateWiresStage5[0][23] , \intermediateWiresStage5[0][22] , 
    \intermediateWiresStage5[0][21] , \intermediateWiresStage5[0][20] , \intermediateWiresStage5[0][19] , 
    \intermediateWiresStage5[0][18] , \intermediateWiresStage5[0][17] , \intermediateWiresStage5[0][16] , 
    \intermediateWiresStage5[0][15] , \intermediateWiresStage5[0][14] , \intermediateWiresStage5[0][13] , 
    \intermediateWiresStage5[0][12] , \intermediateWiresStage5[0][11] , \intermediateWiresStage5[0][10] , 
    \intermediateWiresStage5[0][9] , \intermediateWiresStage5[0][8] , \intermediateWiresStage5[0][7] , 
    \intermediateWiresStage5[0][6] , uc_4294, uc_4295, uc_4296, uc_4297, uc_4298, 
    uc_4299}), .B ({1'b0 , uc_4300, uc_4301, uc_4302, uc_4303, uc_4304, uc_4305, 
    uc_4306, uc_4307, uc_4308, uc_4309, uc_4310, uc_4311, uc_4312, uc_4313, uc_4314, 
    uc_4315, uc_4316, \intermediateWiresStage5[1][45] , \intermediateWiresStage5[1][44] , 
    \intermediateWiresStage5[1][43] , \intermediateWiresStage5[1][42] , \intermediateWiresStage5[1][41] , 
    \intermediateWiresStage5[1][40] , \intermediateWiresStage5[1][39] , \intermediateWiresStage5[1][38] , 
    \intermediateWiresStage5[1][37] , \intermediateWiresStage5[1][36] , \intermediateWiresStage5[1][35] , 
    \intermediateWiresStage5[1][34] , \intermediateWiresStage5[1][33] , \intermediateWiresStage5[1][32] , 
    \intermediateWiresStage5[1][31] , \intermediateWiresStage5[1][30] , \intermediateWiresStage5[1][29] , 
    \intermediateWiresStage5[1][28] , \intermediateWiresStage5[1][27] , \intermediateWiresStage5[1][26] , 
    \intermediateWiresStage5[1][25] , \intermediateWiresStage5[1][24] , \intermediateWiresStage5[1][23] , 
    \intermediateWiresStage5[1][22] , \intermediateWiresStage5[1][21] , \intermediateWiresStage5[1][20] , 
    \intermediateWiresStage5[1][19] , \intermediateWiresStage5[1][18] , \intermediateWiresStage5[1][17] , 
    \intermediateWiresStage5[1][16] , \intermediateWiresStage5[1][15] , \intermediateWiresStage5[1][14] , 
    \intermediateWiresStage5[1][13] , \intermediateWiresStage5[1][12] , \intermediateWiresStage5[1][11] , 
    \intermediateWiresStage5[1][10] , \intermediateWiresStage5[1][9] , \intermediateWiresStage5[1][8] , 
    \intermediateWiresStage5[1][7] , \intermediateWiresStage5[1][6] , uc_4317, uc_4318, 
    uc_4319, uc_4320, uc_4321, uc_4322}), .C ({1'b0 , uc_4323, uc_4324, uc_4325, 
    uc_4326, uc_4327, uc_4328, uc_4329, uc_4330, uc_4331, \intermediateWiresStage5[2][53] , 
    \intermediateWiresStage5[2][52] , \intermediateWiresStage5[2][51] , \intermediateWiresStage5[2][50] , 
    \intermediateWiresStage5[2][49] , \intermediateWiresStage5[2][48] , \intermediateWiresStage5[2][47] , 
    \intermediateWiresStage5[2][46] , \intermediateWiresStage5[2][45] , \intermediateWiresStage5[2][44] , 
    \intermediateWiresStage5[2][43] , \intermediateWiresStage5[2][42] , \intermediateWiresStage5[2][41] , 
    \intermediateWiresStage5[2][40] , \intermediateWiresStage5[2][39] , \intermediateWiresStage5[2][38] , 
    \intermediateWiresStage5[2][37] , \intermediateWiresStage5[2][36] , \intermediateWiresStage5[2][35] , 
    \intermediateWiresStage5[2][34] , \intermediateWiresStage5[2][33] , \intermediateWiresStage5[2][32] , 
    \intermediateWiresStage5[2][31] , \intermediateWiresStage5[2][30] , \intermediateWiresStage5[2][29] , 
    \intermediateWiresStage5[2][28] , \intermediateWiresStage5[2][27] , \intermediateWiresStage5[2][26] , 
    \intermediateWiresStage5[2][25] , \intermediateWiresStage5[2][24] , \intermediateWiresStage5[2][23] , 
    \intermediateWiresStage5[2][22] , \intermediateWiresStage5[2][21] , \intermediateWiresStage4[3][20] , 
    \intermediateWiresStage4[3][19] , \intermediateWiresStage4[3][18] , \intermediateWiresStage4[3][17] , 
    \intermediateWiresStage4[3][16] , \intermediateWiresStage4[3][15] , uc_4332, 
    uc_4333, uc_4334, uc_4335, uc_4336, uc_4337, uc_4338, uc_4339, uc_4340, uc_4341, 
    uc_4342, uc_4343, uc_4344, uc_4345, uc_4346}));
CSAlike__4_1512 genblk6_0_parallelAdderStage5 (.carry ({uc_4150, uc_4151, uc_4152, 
    uc_4153, uc_4154, uc_4155, uc_4156, uc_4157, uc_4158, uc_4159, uc_4160, uc_4161, 
    uc_4162, uc_4163, uc_4164, uc_4165, uc_4166, uc_4167, \intermediateWiresStage5[1][45] , 
    \intermediateWiresStage5[1][44] , \intermediateWiresStage5[1][43] , \intermediateWiresStage5[1][42] , 
    \intermediateWiresStage5[1][41] , \intermediateWiresStage5[1][40] , \intermediateWiresStage5[1][39] , 
    \intermediateWiresStage5[1][38] , \intermediateWiresStage5[1][37] , \intermediateWiresStage5[1][36] , 
    \intermediateWiresStage5[1][35] , \intermediateWiresStage5[1][34] , \intermediateWiresStage5[1][33] , 
    \intermediateWiresStage5[1][32] , \intermediateWiresStage5[1][31] , \intermediateWiresStage5[1][30] , 
    \intermediateWiresStage5[1][29] , \intermediateWiresStage5[1][28] , \intermediateWiresStage5[1][27] , 
    \intermediateWiresStage5[1][26] , \intermediateWiresStage5[1][25] , \intermediateWiresStage5[1][24] , 
    \intermediateWiresStage5[1][23] , \intermediateWiresStage5[1][22] , \intermediateWiresStage5[1][21] , 
    \intermediateWiresStage5[1][20] , \intermediateWiresStage5[1][19] , \intermediateWiresStage5[1][18] , 
    \intermediateWiresStage5[1][17] , \intermediateWiresStage5[1][16] , \intermediateWiresStage5[1][15] , 
    \intermediateWiresStage5[1][14] , \intermediateWiresStage5[1][13] , \intermediateWiresStage5[1][12] , 
    \intermediateWiresStage5[1][11] , \intermediateWiresStage5[1][10] , \intermediateWiresStage5[1][9] , 
    \intermediateWiresStage5[1][8] , \intermediateWiresStage5[1][7] , \intermediateWiresStage5[1][6] , 
    uc_4168, uc_4169, uc_4170, uc_4171, uc_4172, uc_4173}), .result ({uc_4126, uc_4127, 
    uc_4128, uc_4129, uc_4130, uc_4131, uc_4132, uc_4133, uc_4134, uc_4135, uc_4136, 
    uc_4137, uc_4138, uc_4139, uc_4140, uc_4141, uc_4142, uc_4143, uc_4144, \intermediateWiresStage5[0][44] , 
    \intermediateWiresStage5[0][43] , \intermediateWiresStage5[0][42] , \intermediateWiresStage5[0][41] , 
    \intermediateWiresStage5[0][40] , \intermediateWiresStage5[0][39] , \intermediateWiresStage5[0][38] , 
    \intermediateWiresStage5[0][37] , \intermediateWiresStage5[0][36] , \intermediateWiresStage5[0][35] , 
    \intermediateWiresStage5[0][34] , \intermediateWiresStage5[0][33] , \intermediateWiresStage5[0][32] , 
    \intermediateWiresStage5[0][31] , \intermediateWiresStage5[0][30] , \intermediateWiresStage5[0][29] , 
    \intermediateWiresStage5[0][28] , \intermediateWiresStage5[0][27] , \intermediateWiresStage5[0][26] , 
    \intermediateWiresStage5[0][25] , \intermediateWiresStage5[0][24] , \intermediateWiresStage5[0][23] , 
    \intermediateWiresStage5[0][22] , \intermediateWiresStage5[0][21] , \intermediateWiresStage5[0][20] , 
    \intermediateWiresStage5[0][19] , \intermediateWiresStage5[0][18] , \intermediateWiresStage5[0][17] , 
    \intermediateWiresStage5[0][16] , \intermediateWiresStage5[0][15] , \intermediateWiresStage5[0][14] , 
    \intermediateWiresStage5[0][13] , \intermediateWiresStage5[0][12] , \intermediateWiresStage5[0][11] , 
    \intermediateWiresStage5[0][10] , \intermediateWiresStage5[0][9] , \intermediateWiresStage5[0][8] , 
    \intermediateWiresStage5[0][7] , \intermediateWiresStage5[0][6] , Res[5], uc_4145, 
    uc_4146, uc_4147, uc_4148, uc_4149}), .A ({1'b0 , uc_4174, uc_4175, uc_4176, 
    uc_4177, uc_4178, uc_4179, uc_4180, uc_4181, uc_4182, uc_4183, uc_4184, uc_4185, 
    uc_4186, uc_4187, uc_4188, uc_4189, uc_4190, uc_4191, normalizedWires[940], \intermediateWiresStage1[8][43] , 
    \intermediateWiresStage3[2][42] , \intermediateWiresStage3[2][41] , \intermediateWiresStage3[2][40] , 
    \intermediateWiresStage3[2][39] , \intermediateWiresStage4[0][38] , \intermediateWiresStage4[0][37] , 
    \intermediateWiresStage4[0][36] , \intermediateWiresStage4[0][35] , \intermediateWiresStage4[0][34] , 
    \intermediateWiresStage4[0][33] , \intermediateWiresStage4[0][32] , \intermediateWiresStage4[0][31] , 
    \intermediateWiresStage4[0][30] , \intermediateWiresStage4[0][29] , \intermediateWiresStage4[0][28] , 
    \intermediateWiresStage4[0][27] , \intermediateWiresStage4[0][26] , \intermediateWiresStage4[0][25] , 
    \intermediateWiresStage4[0][24] , \intermediateWiresStage4[0][23] , \intermediateWiresStage4[0][22] , 
    \intermediateWiresStage4[0][21] , \intermediateWiresStage4[0][20] , \intermediateWiresStage4[0][19] , 
    \intermediateWiresStage4[0][18] , \intermediateWiresStage4[0][17] , \intermediateWiresStage4[0][16] , 
    \intermediateWiresStage4[0][15] , \intermediateWiresStage4[0][14] , \intermediateWiresStage4[0][13] , 
    \intermediateWiresStage4[0][12] , \intermediateWiresStage4[0][11] , \intermediateWiresStage4[0][10] , 
    \intermediateWiresStage4[0][9] , \intermediateWiresStage4[0][8] , \intermediateWiresStage4[0][7] , 
    \intermediateWiresStage4[0][6] , \intermediateWiresStage4[0][5] , uc_4192, uc_4193, 
    uc_4194, uc_4195, uc_4196}), .B ({1'b0 , uc_4197, uc_4198, uc_4199, uc_4200, 
    uc_4201, uc_4202, uc_4203, uc_4204, uc_4205, uc_4206, uc_4207, uc_4208, uc_4209, 
    uc_4210, uc_4211, uc_4212, uc_4213, uc_4214, uc_4215, uc_4216, uc_4217, uc_4218, 
    uc_4219, \intermediateWiresStage4[1][39] , \intermediateWiresStage4[1][38] , 
    \intermediateWiresStage4[1][37] , \intermediateWiresStage4[1][36] , \intermediateWiresStage4[1][35] , 
    \intermediateWiresStage4[1][34] , \intermediateWiresStage4[1][33] , \intermediateWiresStage4[1][32] , 
    \intermediateWiresStage4[1][31] , \intermediateWiresStage4[1][30] , \intermediateWiresStage4[1][29] , 
    \intermediateWiresStage4[1][28] , \intermediateWiresStage4[1][27] , \intermediateWiresStage4[1][26] , 
    \intermediateWiresStage4[1][25] , \intermediateWiresStage4[1][24] , \intermediateWiresStage4[1][23] , 
    \intermediateWiresStage4[1][22] , \intermediateWiresStage4[1][21] , \intermediateWiresStage4[1][20] , 
    \intermediateWiresStage4[1][19] , \intermediateWiresStage4[1][18] , \intermediateWiresStage4[1][17] , 
    \intermediateWiresStage4[1][16] , \intermediateWiresStage4[1][15] , \intermediateWiresStage4[1][14] , 
    \intermediateWiresStage4[1][13] , \intermediateWiresStage4[1][12] , \intermediateWiresStage4[1][11] , 
    \intermediateWiresStage4[1][10] , \intermediateWiresStage4[1][9] , \intermediateWiresStage4[1][8] , 
    \intermediateWiresStage4[1][7] , \intermediateWiresStage4[1][6] , \intermediateWiresStage4[1][5] , 
    uc_4220, uc_4221, uc_4222, uc_4223, uc_4224}), .C ({1'b0 , uc_4225, uc_4226, 
    uc_4227, uc_4228, uc_4229, uc_4230, uc_4231, uc_4232, uc_4233, uc_4234, uc_4235, 
    uc_4236, uc_4237, uc_4238, uc_4239, uc_4240, uc_4241, uc_4242, \intermediateWiresStage4[2][44] , 
    \intermediateWiresStage4[2][43] , \intermediateWiresStage4[2][42] , \intermediateWiresStage4[2][41] , 
    \intermediateWiresStage4[2][40] , \intermediateWiresStage4[2][39] , \intermediateWiresStage4[2][38] , 
    \intermediateWiresStage4[2][37] , \intermediateWiresStage4[2][36] , \intermediateWiresStage4[2][35] , 
    \intermediateWiresStage4[2][34] , \intermediateWiresStage4[2][33] , \intermediateWiresStage4[2][32] , 
    \intermediateWiresStage4[2][31] , \intermediateWiresStage4[2][30] , \intermediateWiresStage4[2][29] , 
    \intermediateWiresStage4[2][28] , \intermediateWiresStage4[2][27] , \intermediateWiresStage4[2][26] , 
    \intermediateWiresStage4[2][25] , \intermediateWiresStage4[2][24] , \intermediateWiresStage4[2][23] , 
    \intermediateWiresStage4[2][22] , \intermediateWiresStage4[2][21] , \intermediateWiresStage4[2][20] , 
    \intermediateWiresStage4[2][19] , \intermediateWiresStage4[2][18] , \intermediateWiresStage4[2][17] , 
    \intermediateWiresStage4[2][16] , \intermediateWiresStage4[2][15] , \intermediateWiresStage4[2][14] , 
    \intermediateWiresStage3[3][13] , \intermediateWiresStage3[3][12] , \intermediateWiresStage3[3][11] , 
    \intermediateWiresStage3[3][10] , uc_4243, uc_4244, uc_4245, uc_4246, uc_4247, 
    uc_4248, uc_4249, uc_4250, uc_4251, uc_4252}));
CSAlike__4_1259 genblk6_1_parallelAdderStage5 (.carry ({uc_4013, uc_4014, uc_4015, 
    uc_4016, \intermediateWiresStage5[3][59] , \intermediateWiresStage5[3][58] , 
    \intermediateWiresStage5[3][57] , \intermediateWiresStage5[3][56] , \intermediateWiresStage5[3][55] , 
    \intermediateWiresStage5[3][54] , \intermediateWiresStage5[3][53] , \intermediateWiresStage5[3][52] , 
    \intermediateWiresStage5[3][51] , \intermediateWiresStage5[3][50] , \intermediateWiresStage5[3][49] , 
    \intermediateWiresStage5[3][48] , \intermediateWiresStage5[3][47] , \intermediateWiresStage5[3][46] , 
    \intermediateWiresStage5[3][45] , \intermediateWiresStage5[3][44] , \intermediateWiresStage5[3][43] , 
    \intermediateWiresStage5[3][42] , \intermediateWiresStage5[3][41] , \intermediateWiresStage5[3][40] , 
    \intermediateWiresStage5[3][39] , \intermediateWiresStage5[3][38] , \intermediateWiresStage5[3][37] , 
    \intermediateWiresStage5[3][36] , \intermediateWiresStage5[3][35] , \intermediateWiresStage5[3][34] , 
    \intermediateWiresStage5[3][33] , \intermediateWiresStage5[3][32] , \intermediateWiresStage5[3][31] , 
    \intermediateWiresStage5[3][30] , \intermediateWiresStage5[3][29] , \intermediateWiresStage5[3][28] , 
    \intermediateWiresStage5[3][27] , \intermediateWiresStage5[3][26] , \intermediateWiresStage5[3][25] , 
    \intermediateWiresStage5[3][24] , \intermediateWiresStage5[3][23] , \intermediateWiresStage5[3][22] , 
    uc_4017, uc_4018, uc_4019, uc_4020, uc_4021, uc_4022, uc_4023, uc_4024, uc_4025, 
    uc_4026, uc_4027, uc_4028, uc_4029, uc_4030, uc_4031, uc_4032, uc_4033, uc_4034, 
    uc_4035, uc_4036, uc_4037, uc_4038}), .result ({uc_3987, uc_3988, uc_3989, uc_3990, 
    uc_3991, \intermediateWiresStage5[2][58] , \intermediateWiresStage5[2][57] , 
    \intermediateWiresStage5[2][56] , \intermediateWiresStage5[2][55] , \intermediateWiresStage5[2][54] , 
    \intermediateWiresStage5[2][53] , \intermediateWiresStage5[2][52] , \intermediateWiresStage5[2][51] , 
    \intermediateWiresStage5[2][50] , \intermediateWiresStage5[2][49] , \intermediateWiresStage5[2][48] , 
    \intermediateWiresStage5[2][47] , \intermediateWiresStage5[2][46] , \intermediateWiresStage5[2][45] , 
    \intermediateWiresStage5[2][44] , \intermediateWiresStage5[2][43] , \intermediateWiresStage5[2][42] , 
    \intermediateWiresStage5[2][41] , \intermediateWiresStage5[2][40] , \intermediateWiresStage5[2][39] , 
    \intermediateWiresStage5[2][38] , \intermediateWiresStage5[2][37] , \intermediateWiresStage5[2][36] , 
    \intermediateWiresStage5[2][35] , \intermediateWiresStage5[2][34] , \intermediateWiresStage5[2][33] , 
    \intermediateWiresStage5[2][32] , \intermediateWiresStage5[2][31] , \intermediateWiresStage5[2][30] , 
    \intermediateWiresStage5[2][29] , \intermediateWiresStage5[2][28] , \intermediateWiresStage5[2][27] , 
    \intermediateWiresStage5[2][26] , \intermediateWiresStage5[2][25] , \intermediateWiresStage5[2][24] , 
    \intermediateWiresStage5[2][23] , \intermediateWiresStage5[2][22] , \intermediateWiresStage5[2][21] , 
    uc_3992, uc_3993, uc_3994, uc_3995, uc_3996, uc_3997, uc_3998, uc_3999, uc_4000, 
    uc_4001, uc_4002, uc_4003, uc_4004, uc_4005, uc_4006, uc_4007, uc_4008, uc_4009, 
    uc_4010, uc_4011, uc_4012}), .A ({1'b0 , uc_4039, uc_4040, uc_4041, uc_4042, 
    uc_4043, uc_4044, uc_4045, uc_4046, uc_4047, uc_4048, uc_4049, uc_4050, \intermediateWiresStage4[3][50] , 
    \intermediateWiresStage4[3][49] , \intermediateWiresStage4[3][48] , \intermediateWiresStage4[3][47] , 
    \intermediateWiresStage4[3][46] , \intermediateWiresStage4[3][45] , \intermediateWiresStage4[3][44] , 
    \intermediateWiresStage4[3][43] , \intermediateWiresStage4[3][42] , \intermediateWiresStage4[3][41] , 
    \intermediateWiresStage4[3][40] , \intermediateWiresStage4[3][39] , \intermediateWiresStage4[3][38] , 
    \intermediateWiresStage4[3][37] , \intermediateWiresStage4[3][36] , \intermediateWiresStage4[3][35] , 
    \intermediateWiresStage4[3][34] , \intermediateWiresStage4[3][33] , \intermediateWiresStage4[3][32] , 
    \intermediateWiresStage4[3][31] , \intermediateWiresStage4[3][30] , \intermediateWiresStage4[3][29] , 
    \intermediateWiresStage4[3][28] , \intermediateWiresStage4[3][27] , \intermediateWiresStage4[3][26] , 
    \intermediateWiresStage4[3][25] , \intermediateWiresStage4[3][24] , \intermediateWiresStage4[3][23] , 
    \intermediateWiresStage4[3][22] , \intermediateWiresStage4[3][21] , uc_4051, 
    uc_4052, uc_4053, uc_4054, uc_4055, uc_4056, uc_4057, uc_4058, uc_4059, uc_4060, 
    uc_4061, uc_4062, uc_4063, uc_4064, uc_4065, uc_4066, uc_4067, uc_4068, uc_4069, 
    uc_4070, uc_4071}), .B ({1'b0 , uc_4072, uc_4073, uc_4074, uc_4075, \intermediateWiresStage3[8][58] , 
    \intermediateWiresStage4[4][57] , \intermediateWiresStage4[4][56] , \intermediateWiresStage4[4][55] , 
    \intermediateWiresStage4[4][54] , \intermediateWiresStage4[4][53] , \intermediateWiresStage4[4][52] , 
    \intermediateWiresStage4[4][51] , \intermediateWiresStage4[4][50] , \intermediateWiresStage4[4][49] , 
    \intermediateWiresStage4[4][48] , \intermediateWiresStage4[4][47] , \intermediateWiresStage4[4][46] , 
    \intermediateWiresStage4[4][45] , \intermediateWiresStage4[4][44] , \intermediateWiresStage4[4][43] , 
    \intermediateWiresStage4[4][42] , \intermediateWiresStage4[4][41] , \intermediateWiresStage4[4][40] , 
    \intermediateWiresStage4[4][39] , \intermediateWiresStage4[4][38] , \intermediateWiresStage4[4][37] , 
    \intermediateWiresStage4[4][36] , \intermediateWiresStage4[4][35] , \intermediateWiresStage4[4][34] , 
    \intermediateWiresStage4[4][33] , \intermediateWiresStage4[4][32] , \intermediateWiresStage4[4][31] , 
    \intermediateWiresStage4[4][30] , \intermediateWiresStage4[4][29] , \intermediateWiresStage4[4][28] , 
    \intermediateWiresStage4[4][27] , \intermediateWiresStage4[4][26] , \intermediateWiresStage4[4][25] , 
    \intermediateWiresStage4[4][24] , \intermediateWiresStage3[6][23] , \intermediateWiresStage2[9][22] , 
    \intermediateWiresStage2[9][21] , uc_4076, uc_4077, uc_4078, uc_4079, uc_4080, 
    uc_4081, uc_4082, uc_4083, uc_4084, uc_4085, uc_4086, uc_4087, uc_4088, uc_4089, 
    uc_4090, uc_4091, uc_4092, uc_4093, uc_4094, uc_4095, uc_4096}), .C ({1'b0 , 
    uc_4097, uc_4098, uc_4099, uc_4100, \intermediateWiresStage4[5][58] , \intermediateWiresStage4[5][57] , 
    \intermediateWiresStage4[5][56] , \intermediateWiresStage4[5][55] , \intermediateWiresStage4[5][54] , 
    \intermediateWiresStage4[5][53] , \intermediateWiresStage4[5][52] , \intermediateWiresStage4[5][51] , 
    \intermediateWiresStage4[5][50] , \intermediateWiresStage4[5][49] , \intermediateWiresStage4[5][48] , 
    \intermediateWiresStage4[5][47] , \intermediateWiresStage4[5][46] , \intermediateWiresStage4[5][45] , 
    \intermediateWiresStage4[5][44] , \intermediateWiresStage4[5][43] , \intermediateWiresStage4[5][42] , 
    \intermediateWiresStage4[5][41] , \intermediateWiresStage4[5][40] , \intermediateWiresStage4[5][39] , 
    \intermediateWiresStage4[5][38] , \intermediateWiresStage4[5][37] , \intermediateWiresStage4[5][36] , 
    \intermediateWiresStage4[5][35] , \intermediateWiresStage4[5][34] , \intermediateWiresStage4[5][33] , 
    \intermediateWiresStage4[5][32] , \intermediateWiresStage4[5][31] , \intermediateWiresStage4[5][30] , 
    \intermediateWiresStage4[5][29] , \intermediateWiresStage4[5][28] , \intermediateWiresStage4[5][27] , 
    \intermediateWiresStage4[5][26] , \intermediateWiresStage4[5][25] , uc_4101, 
    uc_4102, uc_4103, uc_4104, uc_4105, uc_4106, uc_4107, uc_4108, uc_4109, uc_4110, 
    uc_4111, uc_4112, uc_4113, uc_4114, uc_4115, uc_4116, uc_4117, uc_4118, uc_4119, 
    uc_4120, uc_4121, uc_4122, uc_4123, uc_4124, uc_4125}));
CSAlike__4_1006 genblk5_0_parallelAdderStage4 (.carry ({uc_3869, uc_3870, uc_3871, 
    uc_3872, uc_3873, uc_3874, uc_3875, uc_3876, uc_3877, uc_3878, uc_3879, uc_3880, 
    uc_3881, uc_3882, uc_3883, uc_3884, uc_3885, uc_3886, uc_3887, uc_3888, uc_3889, 
    uc_3890, uc_3891, uc_3892, \intermediateWiresStage4[1][39] , \intermediateWiresStage4[1][38] , 
    \intermediateWiresStage4[1][37] , \intermediateWiresStage4[1][36] , \intermediateWiresStage4[1][35] , 
    \intermediateWiresStage4[1][34] , \intermediateWiresStage4[1][33] , \intermediateWiresStage4[1][32] , 
    \intermediateWiresStage4[1][31] , \intermediateWiresStage4[1][30] , \intermediateWiresStage4[1][29] , 
    \intermediateWiresStage4[1][28] , \intermediateWiresStage4[1][27] , \intermediateWiresStage4[1][26] , 
    \intermediateWiresStage4[1][25] , \intermediateWiresStage4[1][24] , \intermediateWiresStage4[1][23] , 
    \intermediateWiresStage4[1][22] , \intermediateWiresStage4[1][21] , \intermediateWiresStage4[1][20] , 
    \intermediateWiresStage4[1][19] , \intermediateWiresStage4[1][18] , \intermediateWiresStage4[1][17] , 
    \intermediateWiresStage4[1][16] , \intermediateWiresStage4[1][15] , \intermediateWiresStage4[1][14] , 
    \intermediateWiresStage4[1][13] , \intermediateWiresStage4[1][12] , \intermediateWiresStage4[1][11] , 
    \intermediateWiresStage4[1][10] , \intermediateWiresStage4[1][9] , \intermediateWiresStage4[1][8] , 
    \intermediateWiresStage4[1][7] , \intermediateWiresStage4[1][6] , \intermediateWiresStage4[1][5] , 
    uc_3893, uc_3894, uc_3895, uc_3896, uc_3897}), .result ({uc_3840, uc_3841, uc_3842, 
    uc_3843, uc_3844, uc_3845, uc_3846, uc_3847, uc_3848, uc_3849, uc_3850, uc_3851, 
    uc_3852, uc_3853, uc_3854, uc_3855, uc_3856, uc_3857, uc_3858, uc_3859, uc_3860, 
    uc_3861, uc_3862, uc_3863, uc_3864, \intermediateWiresStage4[0][38] , \intermediateWiresStage4[0][37] , 
    \intermediateWiresStage4[0][36] , \intermediateWiresStage4[0][35] , \intermediateWiresStage4[0][34] , 
    \intermediateWiresStage4[0][33] , \intermediateWiresStage4[0][32] , \intermediateWiresStage4[0][31] , 
    \intermediateWiresStage4[0][30] , \intermediateWiresStage4[0][29] , \intermediateWiresStage4[0][28] , 
    \intermediateWiresStage4[0][27] , \intermediateWiresStage4[0][26] , \intermediateWiresStage4[0][25] , 
    \intermediateWiresStage4[0][24] , \intermediateWiresStage4[0][23] , \intermediateWiresStage4[0][22] , 
    \intermediateWiresStage4[0][21] , \intermediateWiresStage4[0][20] , \intermediateWiresStage4[0][19] , 
    \intermediateWiresStage4[0][18] , \intermediateWiresStage4[0][17] , \intermediateWiresStage4[0][16] , 
    \intermediateWiresStage4[0][15] , \intermediateWiresStage4[0][14] , \intermediateWiresStage4[0][13] , 
    \intermediateWiresStage4[0][12] , \intermediateWiresStage4[0][11] , \intermediateWiresStage4[0][10] , 
    \intermediateWiresStage4[0][9] , \intermediateWiresStage4[0][8] , \intermediateWiresStage4[0][7] , 
    \intermediateWiresStage4[0][6] , \intermediateWiresStage4[0][5] , Res[4], uc_3865, 
    uc_3866, uc_3867, uc_3868}), .A ({1'b0 , uc_3898, uc_3899, uc_3900, uc_3901, 
    uc_3902, uc_3903, uc_3904, uc_3905, uc_3906, uc_3907, uc_3908, uc_3909, uc_3910, 
    uc_3911, uc_3912, uc_3913, uc_3914, uc_3915, uc_3916, uc_3917, uc_3918, uc_3919, 
    uc_3920, uc_3921, \intermediateWiresStage2[2][38] , \intermediateWiresStage2[2][37] , 
    \intermediateWiresStage2[2][36] , \intermediateWiresStage3[0][35] , \intermediateWiresStage3[0][34] , 
    \intermediateWiresStage3[0][33] , \intermediateWiresStage3[0][32] , \intermediateWiresStage3[0][31] , 
    \intermediateWiresStage3[0][30] , \intermediateWiresStage3[0][29] , \intermediateWiresStage3[0][28] , 
    \intermediateWiresStage3[0][27] , \intermediateWiresStage3[0][26] , \intermediateWiresStage3[0][25] , 
    \intermediateWiresStage3[0][24] , \intermediateWiresStage3[0][23] , \intermediateWiresStage3[0][22] , 
    \intermediateWiresStage3[0][21] , \intermediateWiresStage3[0][20] , \intermediateWiresStage3[0][19] , 
    \intermediateWiresStage3[0][18] , \intermediateWiresStage3[0][17] , \intermediateWiresStage3[0][16] , 
    \intermediateWiresStage3[0][15] , \intermediateWiresStage3[0][14] , \intermediateWiresStage3[0][13] , 
    \intermediateWiresStage3[0][12] , \intermediateWiresStage3[0][11] , \intermediateWiresStage3[0][10] , 
    \intermediateWiresStage3[0][9] , \intermediateWiresStage3[0][8] , \intermediateWiresStage3[0][7] , 
    \intermediateWiresStage3[0][6] , \intermediateWiresStage3[0][5] , \intermediateWiresStage3[0][4] , 
    uc_3922, uc_3923, uc_3924, uc_3925}), .B ({1'b0 , uc_3926, uc_3927, uc_3928, 
    uc_3929, uc_3930, uc_3931, uc_3932, uc_3933, uc_3934, uc_3935, uc_3936, uc_3937, 
    uc_3938, uc_3939, uc_3940, uc_3941, uc_3942, uc_3943, uc_3944, uc_3945, uc_3946, 
    uc_3947, uc_3948, uc_3949, uc_3950, uc_3951, \intermediateWiresStage3[1][36] , 
    \intermediateWiresStage3[1][35] , \intermediateWiresStage3[1][34] , \intermediateWiresStage3[1][33] , 
    \intermediateWiresStage3[1][32] , \intermediateWiresStage3[1][31] , \intermediateWiresStage3[1][30] , 
    \intermediateWiresStage3[1][29] , \intermediateWiresStage3[1][28] , \intermediateWiresStage3[1][27] , 
    \intermediateWiresStage3[1][26] , \intermediateWiresStage3[1][25] , \intermediateWiresStage3[1][24] , 
    \intermediateWiresStage3[1][23] , \intermediateWiresStage3[1][22] , \intermediateWiresStage3[1][21] , 
    \intermediateWiresStage3[1][20] , \intermediateWiresStage3[1][19] , \intermediateWiresStage3[1][18] , 
    \intermediateWiresStage3[1][17] , \intermediateWiresStage3[1][16] , \intermediateWiresStage3[1][15] , 
    \intermediateWiresStage3[1][14] , \intermediateWiresStage3[1][13] , \intermediateWiresStage3[1][12] , 
    \intermediateWiresStage3[1][11] , \intermediateWiresStage3[1][10] , \intermediateWiresStage3[1][9] , 
    \intermediateWiresStage3[1][8] , \intermediateWiresStage3[1][7] , \intermediateWiresStage3[1][6] , 
    \intermediateWiresStage3[1][5] , \intermediateWiresStage3[1][4] , uc_3952, uc_3953, 
    uc_3954, uc_3955}), .C ({1'b0 , uc_3956, uc_3957, uc_3958, uc_3959, uc_3960, 
    uc_3961, uc_3962, uc_3963, uc_3964, uc_3965, uc_3966, uc_3967, uc_3968, uc_3969, 
    uc_3970, uc_3971, uc_3972, uc_3973, uc_3974, uc_3975, uc_3976, uc_3977, uc_3978, 
    uc_3979, \intermediateWiresStage3[2][38] , \intermediateWiresStage3[2][37] , 
    \intermediateWiresStage3[2][36] , \intermediateWiresStage3[2][35] , \intermediateWiresStage3[2][34] , 
    \intermediateWiresStage3[2][33] , \intermediateWiresStage3[2][32] , \intermediateWiresStage3[2][31] , 
    \intermediateWiresStage3[2][30] , \intermediateWiresStage3[2][29] , \intermediateWiresStage3[2][28] , 
    \intermediateWiresStage3[2][27] , \intermediateWiresStage3[2][26] , \intermediateWiresStage3[2][25] , 
    \intermediateWiresStage3[2][24] , \intermediateWiresStage3[2][23] , \intermediateWiresStage3[2][22] , 
    \intermediateWiresStage3[2][21] , \intermediateWiresStage3[2][20] , \intermediateWiresStage3[2][19] , 
    \intermediateWiresStage3[2][18] , \intermediateWiresStage3[2][17] , \intermediateWiresStage3[2][16] , 
    \intermediateWiresStage3[2][15] , \intermediateWiresStage3[2][14] , \intermediateWiresStage3[2][13] , 
    \intermediateWiresStage3[2][12] , \intermediateWiresStage3[2][11] , \intermediateWiresStage3[2][10] , 
    \intermediateWiresStage3[2][9] , \intermediateWiresStage2[3][8] , \intermediateWiresStage2[3][7] , 
    uc_3980, uc_3981, uc_3982, uc_3983, uc_3984, uc_3985, uc_3986}));
CSAlike__4_753 genblk5_1_parallelAdderStage4 (.carry ({uc_3722, uc_3723, uc_3724, 
    uc_3725, uc_3726, uc_3727, uc_3728, uc_3729, uc_3730, uc_3731, uc_3732, uc_3733, 
    uc_3734, \intermediateWiresStage4[3][50] , \intermediateWiresStage4[3][49] , 
    \intermediateWiresStage4[3][48] , \intermediateWiresStage4[3][47] , \intermediateWiresStage4[3][46] , 
    \intermediateWiresStage4[3][45] , \intermediateWiresStage4[3][44] , \intermediateWiresStage4[3][43] , 
    \intermediateWiresStage4[3][42] , \intermediateWiresStage4[3][41] , \intermediateWiresStage4[3][40] , 
    \intermediateWiresStage4[3][39] , \intermediateWiresStage4[3][38] , \intermediateWiresStage4[3][37] , 
    \intermediateWiresStage4[3][36] , \intermediateWiresStage4[3][35] , \intermediateWiresStage4[3][34] , 
    \intermediateWiresStage4[3][33] , \intermediateWiresStage4[3][32] , \intermediateWiresStage4[3][31] , 
    \intermediateWiresStage4[3][30] , \intermediateWiresStage4[3][29] , \intermediateWiresStage4[3][28] , 
    \intermediateWiresStage4[3][27] , \intermediateWiresStage4[3][26] , \intermediateWiresStage4[3][25] , 
    \intermediateWiresStage4[3][24] , \intermediateWiresStage4[3][23] , \intermediateWiresStage4[3][22] , 
    \intermediateWiresStage4[3][21] , \intermediateWiresStage4[3][20] , \intermediateWiresStage4[3][19] , 
    \intermediateWiresStage4[3][18] , \intermediateWiresStage4[3][17] , \intermediateWiresStage4[3][16] , 
    \intermediateWiresStage4[3][15] , uc_3735, uc_3736, uc_3737, uc_3738, uc_3739, 
    uc_3740, uc_3741, uc_3742, uc_3743, uc_3744, uc_3745, uc_3746, uc_3747, uc_3748, 
    uc_3749}), .result ({uc_3694, uc_3695, uc_3696, uc_3697, uc_3698, uc_3699, uc_3700, 
    uc_3701, uc_3702, uc_3703, uc_3704, uc_3705, uc_3706, uc_3707, \intermediateWiresStage4[2][49] , 
    \intermediateWiresStage4[2][48] , \intermediateWiresStage4[2][47] , \intermediateWiresStage4[2][46] , 
    \intermediateWiresStage4[2][45] , \intermediateWiresStage4[2][44] , \intermediateWiresStage4[2][43] , 
    \intermediateWiresStage4[2][42] , \intermediateWiresStage4[2][41] , \intermediateWiresStage4[2][40] , 
    \intermediateWiresStage4[2][39] , \intermediateWiresStage4[2][38] , \intermediateWiresStage4[2][37] , 
    \intermediateWiresStage4[2][36] , \intermediateWiresStage4[2][35] , \intermediateWiresStage4[2][34] , 
    \intermediateWiresStage4[2][33] , \intermediateWiresStage4[2][32] , \intermediateWiresStage4[2][31] , 
    \intermediateWiresStage4[2][30] , \intermediateWiresStage4[2][29] , \intermediateWiresStage4[2][28] , 
    \intermediateWiresStage4[2][27] , \intermediateWiresStage4[2][26] , \intermediateWiresStage4[2][25] , 
    \intermediateWiresStage4[2][24] , \intermediateWiresStage4[2][23] , \intermediateWiresStage4[2][22] , 
    \intermediateWiresStage4[2][21] , \intermediateWiresStage4[2][20] , \intermediateWiresStage4[2][19] , 
    \intermediateWiresStage4[2][18] , \intermediateWiresStage4[2][17] , \intermediateWiresStage4[2][16] , 
    \intermediateWiresStage4[2][15] , \intermediateWiresStage4[2][14] , uc_3708, 
    uc_3709, uc_3710, uc_3711, uc_3712, uc_3713, uc_3714, uc_3715, uc_3716, uc_3717, 
    uc_3718, uc_3719, uc_3720, uc_3721}), .A ({1'b0 , uc_3750, uc_3751, uc_3752, 
    uc_3753, uc_3754, uc_3755, uc_3756, uc_3757, uc_3758, uc_3759, uc_3760, uc_3761, 
    uc_3762, uc_3763, uc_3764, uc_3765, uc_3766, uc_3767, uc_3768, \intermediateWiresStage3[3][43] , 
    \intermediateWiresStage3[3][42] , \intermediateWiresStage3[3][41] , \intermediateWiresStage3[3][40] , 
    \intermediateWiresStage3[3][39] , \intermediateWiresStage3[3][38] , \intermediateWiresStage3[3][37] , 
    \intermediateWiresStage3[3][36] , \intermediateWiresStage3[3][35] , \intermediateWiresStage3[3][34] , 
    \intermediateWiresStage3[3][33] , \intermediateWiresStage3[3][32] , \intermediateWiresStage3[3][31] , 
    \intermediateWiresStage3[3][30] , \intermediateWiresStage3[3][29] , \intermediateWiresStage3[3][28] , 
    \intermediateWiresStage3[3][27] , \intermediateWiresStage3[3][26] , \intermediateWiresStage3[3][25] , 
    \intermediateWiresStage3[3][24] , \intermediateWiresStage3[3][23] , \intermediateWiresStage3[3][22] , 
    \intermediateWiresStage3[3][21] , \intermediateWiresStage3[3][20] , \intermediateWiresStage3[3][19] , 
    \intermediateWiresStage3[3][18] , \intermediateWiresStage3[3][17] , \intermediateWiresStage3[3][16] , 
    \intermediateWiresStage3[3][15] , \intermediateWiresStage3[3][14] , uc_3769, 
    uc_3770, uc_3771, uc_3772, uc_3773, uc_3774, uc_3775, uc_3776, uc_3777, uc_3778, 
    uc_3779, uc_3780, uc_3781, uc_3782}), .B ({1'b0 , uc_3783, uc_3784, uc_3785, 
    uc_3786, uc_3787, uc_3788, uc_3789, uc_3790, uc_3791, uc_3792, uc_3793, uc_3794, 
    uc_3795, \intermediateWiresStage2[8][49] , \intermediateWiresStage3[4][48] , 
    \intermediateWiresStage3[4][47] , \intermediateWiresStage3[4][46] , \intermediateWiresStage3[4][45] , 
    \intermediateWiresStage3[4][44] , \intermediateWiresStage3[4][43] , \intermediateWiresStage3[4][42] , 
    \intermediateWiresStage3[4][41] , \intermediateWiresStage3[4][40] , \intermediateWiresStage3[4][39] , 
    \intermediateWiresStage3[4][38] , \intermediateWiresStage3[4][37] , \intermediateWiresStage3[4][36] , 
    \intermediateWiresStage3[4][35] , \intermediateWiresStage3[4][34] , \intermediateWiresStage3[4][33] , 
    \intermediateWiresStage3[4][32] , \intermediateWiresStage3[4][31] , \intermediateWiresStage3[4][30] , 
    \intermediateWiresStage3[4][29] , \intermediateWiresStage3[4][28] , \intermediateWiresStage3[4][27] , 
    \intermediateWiresStage3[4][26] , \intermediateWiresStage3[4][25] , \intermediateWiresStage3[4][24] , 
    \intermediateWiresStage3[4][23] , \intermediateWiresStage3[4][22] , \intermediateWiresStage3[4][21] , 
    \intermediateWiresStage3[4][20] , \intermediateWiresStage3[4][19] , \intermediateWiresStage3[4][18] , 
    \intermediateWiresStage3[4][17] , \intermediateWiresStage3[4][16] , \intermediateWiresStage2[6][15] , 
    \intermediateWiresStage1[9][14] , uc_3796, uc_3797, uc_3798, uc_3799, uc_3800, 
    uc_3801, uc_3802, uc_3803, uc_3804, uc_3805, uc_3806, uc_3807, uc_3808, uc_3809})
    , .C ({1'b0 , uc_3810, uc_3811, uc_3812, uc_3813, uc_3814, uc_3815, uc_3816, 
    uc_3817, uc_3818, uc_3819, uc_3820, uc_3821, uc_3822, \intermediateWiresStage3[5][49] , 
    \intermediateWiresStage3[5][48] , \intermediateWiresStage3[5][47] , \intermediateWiresStage3[5][46] , 
    \intermediateWiresStage3[5][45] , \intermediateWiresStage3[5][44] , \intermediateWiresStage3[5][43] , 
    \intermediateWiresStage3[5][42] , \intermediateWiresStage3[5][41] , \intermediateWiresStage3[5][40] , 
    \intermediateWiresStage3[5][39] , \intermediateWiresStage3[5][38] , \intermediateWiresStage3[5][37] , 
    \intermediateWiresStage3[5][36] , \intermediateWiresStage3[5][35] , \intermediateWiresStage3[5][34] , 
    \intermediateWiresStage3[5][33] , \intermediateWiresStage3[5][32] , \intermediateWiresStage3[5][31] , 
    \intermediateWiresStage3[5][30] , \intermediateWiresStage3[5][29] , \intermediateWiresStage3[5][28] , 
    \intermediateWiresStage3[5][27] , \intermediateWiresStage3[5][26] , \intermediateWiresStage3[5][25] , 
    \intermediateWiresStage3[5][24] , \intermediateWiresStage3[5][23] , \intermediateWiresStage3[5][22] , 
    \intermediateWiresStage3[5][21] , \intermediateWiresStage3[5][20] , \intermediateWiresStage3[5][19] , 
    \intermediateWiresStage3[5][18] , \intermediateWiresStage3[5][17] , uc_3823, 
    uc_3824, uc_3825, uc_3826, uc_3827, uc_3828, uc_3829, uc_3830, uc_3831, uc_3832, 
    uc_3833, uc_3834, uc_3835, uc_3836, uc_3837, uc_3838, uc_3839}));
CSAlike__4_500 genblk5_2_parallelAdderStage4 (.carry ({uc_3574, uc_3575, uc_3576, 
    uc_3577, uc_3578, \intermediateWiresStage4[5][58] , \intermediateWiresStage4[5][57] , 
    \intermediateWiresStage4[5][56] , \intermediateWiresStage4[5][55] , \intermediateWiresStage4[5][54] , 
    \intermediateWiresStage4[5][53] , \intermediateWiresStage4[5][52] , \intermediateWiresStage4[5][51] , 
    \intermediateWiresStage4[5][50] , \intermediateWiresStage4[5][49] , \intermediateWiresStage4[5][48] , 
    \intermediateWiresStage4[5][47] , \intermediateWiresStage4[5][46] , \intermediateWiresStage4[5][45] , 
    \intermediateWiresStage4[5][44] , \intermediateWiresStage4[5][43] , \intermediateWiresStage4[5][42] , 
    \intermediateWiresStage4[5][41] , \intermediateWiresStage4[5][40] , \intermediateWiresStage4[5][39] , 
    \intermediateWiresStage4[5][38] , \intermediateWiresStage4[5][37] , \intermediateWiresStage4[5][36] , 
    \intermediateWiresStage4[5][35] , \intermediateWiresStage4[5][34] , \intermediateWiresStage4[5][33] , 
    \intermediateWiresStage4[5][32] , \intermediateWiresStage4[5][31] , \intermediateWiresStage4[5][30] , 
    \intermediateWiresStage4[5][29] , \intermediateWiresStage4[5][28] , \intermediateWiresStage4[5][27] , 
    \intermediateWiresStage4[5][26] , \intermediateWiresStage4[5][25] , uc_3579, 
    uc_3580, uc_3581, uc_3582, uc_3583, uc_3584, uc_3585, uc_3586, uc_3587, uc_3588, 
    uc_3589, uc_3590, uc_3591, uc_3592, uc_3593, uc_3594, uc_3595, uc_3596, uc_3597, 
    uc_3598, uc_3599, uc_3600, uc_3601, uc_3602, uc_3603}), .result ({uc_3544, uc_3545, 
    uc_3546, uc_3547, uc_3548, uc_3549, \intermediateWiresStage4[4][57] , \intermediateWiresStage4[4][56] , 
    \intermediateWiresStage4[4][55] , \intermediateWiresStage4[4][54] , \intermediateWiresStage4[4][53] , 
    \intermediateWiresStage4[4][52] , \intermediateWiresStage4[4][51] , \intermediateWiresStage4[4][50] , 
    \intermediateWiresStage4[4][49] , \intermediateWiresStage4[4][48] , \intermediateWiresStage4[4][47] , 
    \intermediateWiresStage4[4][46] , \intermediateWiresStage4[4][45] , \intermediateWiresStage4[4][44] , 
    \intermediateWiresStage4[4][43] , \intermediateWiresStage4[4][42] , \intermediateWiresStage4[4][41] , 
    \intermediateWiresStage4[4][40] , \intermediateWiresStage4[4][39] , \intermediateWiresStage4[4][38] , 
    \intermediateWiresStage4[4][37] , \intermediateWiresStage4[4][36] , \intermediateWiresStage4[4][35] , 
    \intermediateWiresStage4[4][34] , \intermediateWiresStage4[4][33] , \intermediateWiresStage4[4][32] , 
    \intermediateWiresStage4[4][31] , \intermediateWiresStage4[4][30] , \intermediateWiresStage4[4][29] , 
    \intermediateWiresStage4[4][28] , \intermediateWiresStage4[4][27] , \intermediateWiresStage4[4][26] , 
    \intermediateWiresStage4[4][25] , \intermediateWiresStage4[4][24] , uc_3550, 
    uc_3551, uc_3552, uc_3553, uc_3554, uc_3555, uc_3556, uc_3557, uc_3558, uc_3559, 
    uc_3560, uc_3561, uc_3562, uc_3563, uc_3564, uc_3565, uc_3566, uc_3567, uc_3568, 
    uc_3569, uc_3570, uc_3571, uc_3572, uc_3573}), .A ({1'b0 , uc_3604, uc_3605, 
    uc_3606, uc_3607, uc_3608, \intermediateWiresStage2[11][57] , \intermediateWiresStage3[6][56] , 
    \intermediateWiresStage3[6][55] , \intermediateWiresStage3[6][54] , \intermediateWiresStage3[6][53] , 
    \intermediateWiresStage3[6][52] , \intermediateWiresStage3[6][51] , \intermediateWiresStage3[6][50] , 
    \intermediateWiresStage3[6][49] , \intermediateWiresStage3[6][48] , \intermediateWiresStage3[6][47] , 
    \intermediateWiresStage3[6][46] , \intermediateWiresStage3[6][45] , \intermediateWiresStage3[6][44] , 
    \intermediateWiresStage3[6][43] , \intermediateWiresStage3[6][42] , \intermediateWiresStage3[6][41] , 
    \intermediateWiresStage3[6][40] , \intermediateWiresStage3[6][39] , \intermediateWiresStage3[6][38] , 
    \intermediateWiresStage3[6][37] , \intermediateWiresStage3[6][36] , \intermediateWiresStage3[6][35] , 
    \intermediateWiresStage3[6][34] , \intermediateWiresStage3[6][33] , \intermediateWiresStage3[6][32] , 
    \intermediateWiresStage3[6][31] , \intermediateWiresStage3[6][30] , \intermediateWiresStage3[6][29] , 
    \intermediateWiresStage3[6][28] , \intermediateWiresStage3[6][27] , \intermediateWiresStage3[6][26] , 
    \intermediateWiresStage3[6][25] , \intermediateWiresStage3[6][24] , uc_3609, 
    uc_3610, uc_3611, uc_3612, uc_3613, uc_3614, uc_3615, uc_3616, uc_3617, uc_3618, 
    uc_3619, uc_3620, uc_3621, uc_3622, uc_3623, uc_3624, uc_3625, uc_3626, uc_3627, 
    uc_3628, uc_3629, uc_3630, uc_3631, uc_3632}), .B ({1'b0 , uc_3633, uc_3634, 
    uc_3635, uc_3636, uc_3637, \intermediateWiresStage3[7][57] , \intermediateWiresStage3[7][56] , 
    \intermediateWiresStage3[7][55] , \intermediateWiresStage3[7][54] , \intermediateWiresStage3[7][53] , 
    \intermediateWiresStage3[7][52] , \intermediateWiresStage3[7][51] , \intermediateWiresStage3[7][50] , 
    \intermediateWiresStage3[7][49] , \intermediateWiresStage3[7][48] , \intermediateWiresStage3[7][47] , 
    \intermediateWiresStage3[7][46] , \intermediateWiresStage3[7][45] , \intermediateWiresStage3[7][44] , 
    \intermediateWiresStage3[7][43] , \intermediateWiresStage3[7][42] , \intermediateWiresStage3[7][41] , 
    \intermediateWiresStage3[7][40] , \intermediateWiresStage3[7][39] , \intermediateWiresStage3[7][38] , 
    \intermediateWiresStage3[7][37] , \intermediateWiresStage3[7][36] , \intermediateWiresStage3[7][35] , 
    \intermediateWiresStage3[7][34] , \intermediateWiresStage3[7][33] , \intermediateWiresStage3[7][32] , 
    \intermediateWiresStage3[7][31] , \intermediateWiresStage3[7][30] , \intermediateWiresStage3[7][29] , 
    \intermediateWiresStage3[7][28] , \intermediateWiresStage3[7][27] , \intermediateWiresStage3[7][26] , 
    \intermediateWiresStage3[7][25] , \intermediateWiresStage3[7][24] , uc_3638, 
    uc_3639, uc_3640, uc_3641, uc_3642, uc_3643, uc_3644, uc_3645, uc_3646, uc_3647, 
    uc_3648, uc_3649, uc_3650, uc_3651, uc_3652, uc_3653, uc_3654, uc_3655, uc_3656, 
    uc_3657, uc_3658, uc_3659, uc_3660, uc_3661}), .C ({1'b0 , uc_3662, uc_3663, 
    uc_3664, uc_3665, uc_3666, \intermediateWiresStage3[8][57] , \intermediateWiresStage3[8][56] , 
    \intermediateWiresStage3[8][55] , \intermediateWiresStage3[8][54] , \intermediateWiresStage3[8][53] , 
    \intermediateWiresStage3[8][52] , \intermediateWiresStage3[8][51] , \intermediateWiresStage3[8][50] , 
    \intermediateWiresStage3[8][49] , \intermediateWiresStage3[8][48] , \intermediateWiresStage3[8][47] , 
    \intermediateWiresStage3[8][46] , \intermediateWiresStage3[8][45] , \intermediateWiresStage3[8][44] , 
    \intermediateWiresStage3[8][43] , \intermediateWiresStage3[8][42] , \intermediateWiresStage3[8][41] , 
    \intermediateWiresStage3[8][40] , \intermediateWiresStage3[8][39] , \intermediateWiresStage3[8][38] , 
    \intermediateWiresStage3[8][37] , \intermediateWiresStage3[8][36] , \intermediateWiresStage3[8][35] , 
    \intermediateWiresStage3[8][34] , \intermediateWiresStage3[8][33] , \intermediateWiresStage3[8][32] , 
    \intermediateWiresStage3[8][31] , \intermediateWiresStage3[8][30] , \intermediateWiresStage2[12][29] , 
    \intermediateWiresStage1[18][28] , normalizedWires[1755], uc_3667, uc_3668, uc_3669, 
    uc_3670, uc_3671, uc_3672, uc_3673, uc_3674, uc_3675, uc_3676, uc_3677, uc_3678, 
    uc_3679, uc_3680, uc_3681, uc_3682, uc_3683, uc_3684, uc_3685, uc_3686, uc_3687, 
    uc_3688, uc_3689, uc_3690, uc_3691, uc_3692, uc_3693}));
CSAlike__0_118 genblk4_0_parallelAdderStage3 (.carry ({uc_3419, uc_3420, uc_3421, 
    uc_3422, uc_3423, uc_3424, uc_3425, uc_3426, uc_3427, uc_3428, uc_3429, uc_3430, 
    uc_3431, uc_3432, uc_3433, uc_3434, uc_3435, uc_3436, uc_3437, uc_3438, uc_3439, 
    uc_3440, uc_3441, uc_3442, uc_3443, uc_3444, uc_3445, \intermediateWiresStage3[1][36] , 
    \intermediateWiresStage3[1][35] , \intermediateWiresStage3[1][34] , \intermediateWiresStage3[1][33] , 
    \intermediateWiresStage3[1][32] , \intermediateWiresStage3[1][31] , \intermediateWiresStage3[1][30] , 
    \intermediateWiresStage3[1][29] , \intermediateWiresStage3[1][28] , \intermediateWiresStage3[1][27] , 
    \intermediateWiresStage3[1][26] , \intermediateWiresStage3[1][25] , \intermediateWiresStage3[1][24] , 
    \intermediateWiresStage3[1][23] , \intermediateWiresStage3[1][22] , \intermediateWiresStage3[1][21] , 
    \intermediateWiresStage3[1][20] , \intermediateWiresStage3[1][19] , \intermediateWiresStage3[1][18] , 
    \intermediateWiresStage3[1][17] , \intermediateWiresStage3[1][16] , \intermediateWiresStage3[1][15] , 
    \intermediateWiresStage3[1][14] , \intermediateWiresStage3[1][13] , \intermediateWiresStage3[1][12] , 
    \intermediateWiresStage3[1][11] , \intermediateWiresStage3[1][10] , \intermediateWiresStage3[1][9] , 
    \intermediateWiresStage3[1][8] , \intermediateWiresStage3[1][7] , \intermediateWiresStage3[1][6] , 
    \intermediateWiresStage3[1][5] , \intermediateWiresStage3[1][4] , uc_3446, uc_3447, 
    uc_3448, uc_3449}), .result ({uc_3388, uc_3389, uc_3390, uc_3391, uc_3392, uc_3393, 
    uc_3394, uc_3395, uc_3396, uc_3397, uc_3398, uc_3399, uc_3400, uc_3401, uc_3402, 
    uc_3403, uc_3404, uc_3405, uc_3406, uc_3407, uc_3408, uc_3409, uc_3410, uc_3411, 
    uc_3412, uc_3413, uc_3414, uc_3415, \intermediateWiresStage3[0][35] , \intermediateWiresStage3[0][34] , 
    \intermediateWiresStage3[0][33] , \intermediateWiresStage3[0][32] , \intermediateWiresStage3[0][31] , 
    \intermediateWiresStage3[0][30] , \intermediateWiresStage3[0][29] , \intermediateWiresStage3[0][28] , 
    \intermediateWiresStage3[0][27] , \intermediateWiresStage3[0][26] , \intermediateWiresStage3[0][25] , 
    \intermediateWiresStage3[0][24] , \intermediateWiresStage3[0][23] , \intermediateWiresStage3[0][22] , 
    \intermediateWiresStage3[0][21] , \intermediateWiresStage3[0][20] , \intermediateWiresStage3[0][19] , 
    \intermediateWiresStage3[0][18] , \intermediateWiresStage3[0][17] , \intermediateWiresStage3[0][16] , 
    \intermediateWiresStage3[0][15] , \intermediateWiresStage3[0][14] , \intermediateWiresStage3[0][13] , 
    \intermediateWiresStage3[0][12] , \intermediateWiresStage3[0][11] , \intermediateWiresStage3[0][10] , 
    \intermediateWiresStage3[0][9] , \intermediateWiresStage3[0][8] , \intermediateWiresStage3[0][7] , 
    \intermediateWiresStage3[0][6] , \intermediateWiresStage3[0][5] , \intermediateWiresStage3[0][4] , 
    Res[3], uc_3416, uc_3417, uc_3418}), .A ({1'b0 , uc_3450, uc_3451, uc_3452, uc_3453, 
    uc_3454, uc_3455, uc_3456, uc_3457, uc_3458, uc_3459, uc_3460, uc_3461, uc_3462, 
    uc_3463, uc_3464, uc_3465, uc_3466, uc_3467, uc_3468, uc_3469, uc_3470, uc_3471, 
    uc_3472, uc_3473, uc_3474, uc_3475, uc_3476, normalizedWires[355], \intermediateWiresStage1[2][34] , 
    \intermediateWiresStage1[2][33] , \intermediateWiresStage2[0][32] , \intermediateWiresStage2[0][31] , 
    \intermediateWiresStage2[0][30] , \intermediateWiresStage2[0][29] , \intermediateWiresStage2[0][28] , 
    \intermediateWiresStage2[0][27] , \intermediateWiresStage2[0][26] , \intermediateWiresStage2[0][25] , 
    \intermediateWiresStage2[0][24] , \intermediateWiresStage2[0][23] , \intermediateWiresStage2[0][22] , 
    \intermediateWiresStage2[0][21] , \intermediateWiresStage2[0][20] , \intermediateWiresStage2[0][19] , 
    \intermediateWiresStage2[0][18] , \intermediateWiresStage2[0][17] , \intermediateWiresStage2[0][16] , 
    \intermediateWiresStage2[0][15] , \intermediateWiresStage2[0][14] , \intermediateWiresStage2[0][13] , 
    \intermediateWiresStage2[0][12] , \intermediateWiresStage2[0][11] , \intermediateWiresStage2[0][10] , 
    \intermediateWiresStage2[0][9] , \intermediateWiresStage2[0][8] , \intermediateWiresStage2[0][7] , 
    \intermediateWiresStage2[0][6] , \intermediateWiresStage2[0][5] , \intermediateWiresStage2[0][4] , 
    \intermediateWiresStage2[0][3] , uc_3477, uc_3478, uc_3479}), .B ({1'b0 , uc_3480, 
    uc_3481, uc_3482, uc_3483, uc_3484, uc_3485, uc_3486, uc_3487, uc_3488, uc_3489, 
    uc_3490, uc_3491, uc_3492, uc_3493, uc_3494, uc_3495, uc_3496, uc_3497, uc_3498, 
    uc_3499, uc_3500, uc_3501, uc_3502, uc_3503, uc_3504, uc_3505, uc_3506, uc_3507, 
    uc_3508, \intermediateWiresStage2[1][33] , \intermediateWiresStage2[1][32] , 
    \intermediateWiresStage2[1][31] , \intermediateWiresStage2[1][30] , \intermediateWiresStage2[1][29] , 
    \intermediateWiresStage2[1][28] , \intermediateWiresStage2[1][27] , \intermediateWiresStage2[1][26] , 
    \intermediateWiresStage2[1][25] , \intermediateWiresStage2[1][24] , \intermediateWiresStage2[1][23] , 
    \intermediateWiresStage2[1][22] , \intermediateWiresStage2[1][21] , \intermediateWiresStage2[1][20] , 
    \intermediateWiresStage2[1][19] , \intermediateWiresStage2[1][18] , \intermediateWiresStage2[1][17] , 
    \intermediateWiresStage2[1][16] , \intermediateWiresStage2[1][15] , \intermediateWiresStage2[1][14] , 
    \intermediateWiresStage2[1][13] , \intermediateWiresStage2[1][12] , \intermediateWiresStage2[1][11] , 
    \intermediateWiresStage2[1][10] , \intermediateWiresStage2[1][9] , \intermediateWiresStage2[1][8] , 
    \intermediateWiresStage2[1][7] , \intermediateWiresStage2[1][6] , \intermediateWiresStage2[1][5] , 
    \intermediateWiresStage2[1][4] , \intermediateWiresStage2[1][3] , uc_3509, uc_3510, 
    uc_3511}), .C ({1'b0 , uc_3512, uc_3513, uc_3514, uc_3515, uc_3516, uc_3517, 
    uc_3518, uc_3519, uc_3520, uc_3521, uc_3522, uc_3523, uc_3524, uc_3525, uc_3526, 
    uc_3527, uc_3528, uc_3529, uc_3530, uc_3531, uc_3532, uc_3533, uc_3534, uc_3535, 
    uc_3536, uc_3537, uc_3538, \intermediateWiresStage2[2][35] , \intermediateWiresStage2[2][34] , 
    \intermediateWiresStage2[2][33] , \intermediateWiresStage2[2][32] , \intermediateWiresStage2[2][31] , 
    \intermediateWiresStage2[2][30] , \intermediateWiresStage2[2][29] , \intermediateWiresStage2[2][28] , 
    \intermediateWiresStage2[2][27] , \intermediateWiresStage2[2][26] , \intermediateWiresStage2[2][25] , 
    \intermediateWiresStage2[2][24] , \intermediateWiresStage2[2][23] , \intermediateWiresStage2[2][22] , 
    \intermediateWiresStage2[2][21] , \intermediateWiresStage2[2][20] , \intermediateWiresStage2[2][19] , 
    \intermediateWiresStage2[2][18] , \intermediateWiresStage2[2][17] , \intermediateWiresStage2[2][16] , 
    \intermediateWiresStage2[2][15] , \intermediateWiresStage2[2][14] , \intermediateWiresStage2[2][13] , 
    \intermediateWiresStage2[2][12] , \intermediateWiresStage2[2][11] , \intermediateWiresStage2[2][10] , 
    \intermediateWiresStage2[2][9] , \intermediateWiresStage2[2][8] , \intermediateWiresStage2[2][7] , 
    \intermediateWiresStage2[2][6] , \intermediateWiresStage1[3][5] , uc_3539, uc_3540, 
    uc_3541, uc_3542, uc_3543}));
CSAlike__3_1259 genblk4_1_parallelAdderStage3 (.carry ({uc_3265, uc_3266, uc_3267, 
    uc_3268, uc_3269, uc_3270, uc_3271, uc_3272, uc_3273, uc_3274, uc_3275, uc_3276, 
    uc_3277, uc_3278, uc_3279, uc_3280, uc_3281, uc_3282, uc_3283, uc_3284, \intermediateWiresStage3[3][43] , 
    \intermediateWiresStage3[3][42] , \intermediateWiresStage3[3][41] , \intermediateWiresStage3[3][40] , 
    \intermediateWiresStage3[3][39] , \intermediateWiresStage3[3][38] , \intermediateWiresStage3[3][37] , 
    \intermediateWiresStage3[3][36] , \intermediateWiresStage3[3][35] , \intermediateWiresStage3[3][34] , 
    \intermediateWiresStage3[3][33] , \intermediateWiresStage3[3][32] , \intermediateWiresStage3[3][31] , 
    \intermediateWiresStage3[3][30] , \intermediateWiresStage3[3][29] , \intermediateWiresStage3[3][28] , 
    \intermediateWiresStage3[3][27] , \intermediateWiresStage3[3][26] , \intermediateWiresStage3[3][25] , 
    \intermediateWiresStage3[3][24] , \intermediateWiresStage3[3][23] , \intermediateWiresStage3[3][22] , 
    \intermediateWiresStage3[3][21] , \intermediateWiresStage3[3][20] , \intermediateWiresStage3[3][19] , 
    \intermediateWiresStage3[3][18] , \intermediateWiresStage3[3][17] , \intermediateWiresStage3[3][16] , 
    \intermediateWiresStage3[3][15] , \intermediateWiresStage3[3][14] , \intermediateWiresStage3[3][13] , 
    \intermediateWiresStage3[3][12] , \intermediateWiresStage3[3][11] , \intermediateWiresStage3[3][10] , 
    uc_3285, uc_3286, uc_3287, uc_3288, uc_3289, uc_3290, uc_3291, uc_3292, uc_3293, 
    uc_3294}), .result ({uc_3235, uc_3236, uc_3237, uc_3238, uc_3239, uc_3240, uc_3241, 
    uc_3242, uc_3243, uc_3244, uc_3245, uc_3246, uc_3247, uc_3248, uc_3249, uc_3250, 
    uc_3251, uc_3252, uc_3253, uc_3254, uc_3255, \intermediateWiresStage3[2][42] , 
    \intermediateWiresStage3[2][41] , \intermediateWiresStage3[2][40] , \intermediateWiresStage3[2][39] , 
    \intermediateWiresStage3[2][38] , \intermediateWiresStage3[2][37] , \intermediateWiresStage3[2][36] , 
    \intermediateWiresStage3[2][35] , \intermediateWiresStage3[2][34] , \intermediateWiresStage3[2][33] , 
    \intermediateWiresStage3[2][32] , \intermediateWiresStage3[2][31] , \intermediateWiresStage3[2][30] , 
    \intermediateWiresStage3[2][29] , \intermediateWiresStage3[2][28] , \intermediateWiresStage3[2][27] , 
    \intermediateWiresStage3[2][26] , \intermediateWiresStage3[2][25] , \intermediateWiresStage3[2][24] , 
    \intermediateWiresStage3[2][23] , \intermediateWiresStage3[2][22] , \intermediateWiresStage3[2][21] , 
    \intermediateWiresStage3[2][20] , \intermediateWiresStage3[2][19] , \intermediateWiresStage3[2][18] , 
    \intermediateWiresStage3[2][17] , \intermediateWiresStage3[2][16] , \intermediateWiresStage3[2][15] , 
    \intermediateWiresStage3[2][14] , \intermediateWiresStage3[2][13] , \intermediateWiresStage3[2][12] , 
    \intermediateWiresStage3[2][11] , \intermediateWiresStage3[2][10] , \intermediateWiresStage3[2][9] , 
    uc_3256, uc_3257, uc_3258, uc_3259, uc_3260, uc_3261, uc_3262, uc_3263, uc_3264})
    , .A ({1'b0 , uc_3295, uc_3296, uc_3297, uc_3298, uc_3299, uc_3300, uc_3301, 
    uc_3302, uc_3303, uc_3304, uc_3305, uc_3306, uc_3307, uc_3308, uc_3309, uc_3310, 
    uc_3311, uc_3312, uc_3313, uc_3314, uc_3315, uc_3316, uc_3317, \intermediateWiresStage2[3][39] , 
    \intermediateWiresStage2[3][38] , \intermediateWiresStage2[3][37] , \intermediateWiresStage2[3][36] , 
    \intermediateWiresStage2[3][35] , \intermediateWiresStage2[3][34] , \intermediateWiresStage2[3][33] , 
    \intermediateWiresStage2[3][32] , \intermediateWiresStage2[3][31] , \intermediateWiresStage2[3][30] , 
    \intermediateWiresStage2[3][29] , \intermediateWiresStage2[3][28] , \intermediateWiresStage2[3][27] , 
    \intermediateWiresStage2[3][26] , \intermediateWiresStage2[3][25] , \intermediateWiresStage2[3][24] , 
    \intermediateWiresStage2[3][23] , \intermediateWiresStage2[3][22] , \intermediateWiresStage2[3][21] , 
    \intermediateWiresStage2[3][20] , \intermediateWiresStage2[3][19] , \intermediateWiresStage2[3][18] , 
    \intermediateWiresStage2[3][17] , \intermediateWiresStage2[3][16] , \intermediateWiresStage2[3][15] , 
    \intermediateWiresStage2[3][14] , \intermediateWiresStage2[3][13] , \intermediateWiresStage2[3][12] , 
    \intermediateWiresStage2[3][11] , \intermediateWiresStage2[3][10] , \intermediateWiresStage2[3][9] , 
    uc_3318, uc_3319, uc_3320, uc_3321, uc_3322, uc_3323, uc_3324, uc_3325, uc_3326})
    , .B ({1'b0 , uc_3327, uc_3328, uc_3329, uc_3330, uc_3331, uc_3332, uc_3333, 
    uc_3334, uc_3335, uc_3336, uc_3337, uc_3338, uc_3339, uc_3340, uc_3341, uc_3342, 
    uc_3343, uc_3344, uc_3345, uc_3346, \intermediateWiresStage1[8][42] , \intermediateWiresStage2[4][41] , 
    \intermediateWiresStage2[4][40] , \intermediateWiresStage2[4][39] , \intermediateWiresStage2[4][38] , 
    \intermediateWiresStage2[4][37] , \intermediateWiresStage2[4][36] , \intermediateWiresStage2[4][35] , 
    \intermediateWiresStage2[4][34] , \intermediateWiresStage2[4][33] , \intermediateWiresStage2[4][32] , 
    \intermediateWiresStage2[4][31] , \intermediateWiresStage2[4][30] , \intermediateWiresStage2[4][29] , 
    \intermediateWiresStage2[4][28] , \intermediateWiresStage2[4][27] , \intermediateWiresStage2[4][26] , 
    \intermediateWiresStage2[4][25] , \intermediateWiresStage2[4][24] , \intermediateWiresStage2[4][23] , 
    \intermediateWiresStage2[4][22] , \intermediateWiresStage2[4][21] , \intermediateWiresStage2[4][20] , 
    \intermediateWiresStage2[4][19] , \intermediateWiresStage2[4][18] , \intermediateWiresStage2[4][17] , 
    \intermediateWiresStage2[4][16] , \intermediateWiresStage2[4][15] , \intermediateWiresStage2[4][14] , 
    \intermediateWiresStage2[4][13] , \intermediateWiresStage2[4][12] , \intermediateWiresStage2[4][11] , 
    \intermediateWiresStage1[6][10] , normalizedWires[585], uc_3347, uc_3348, uc_3349, 
    uc_3350, uc_3351, uc_3352, uc_3353, uc_3354, uc_3355}), .C ({1'b0 , uc_3356, 
    uc_3357, uc_3358, uc_3359, uc_3360, uc_3361, uc_3362, uc_3363, uc_3364, uc_3365, 
    uc_3366, uc_3367, uc_3368, uc_3369, uc_3370, uc_3371, uc_3372, uc_3373, uc_3374, 
    uc_3375, \intermediateWiresStage2[5][42] , \intermediateWiresStage2[5][41] , 
    \intermediateWiresStage2[5][40] , \intermediateWiresStage2[5][39] , \intermediateWiresStage2[5][38] , 
    \intermediateWiresStage2[5][37] , \intermediateWiresStage2[5][36] , \intermediateWiresStage2[5][35] , 
    \intermediateWiresStage2[5][34] , \intermediateWiresStage2[5][33] , \intermediateWiresStage2[5][32] , 
    \intermediateWiresStage2[5][31] , \intermediateWiresStage2[5][30] , \intermediateWiresStage2[5][29] , 
    \intermediateWiresStage2[5][28] , \intermediateWiresStage2[5][27] , \intermediateWiresStage2[5][26] , 
    \intermediateWiresStage2[5][25] , \intermediateWiresStage2[5][24] , \intermediateWiresStage2[5][23] , 
    \intermediateWiresStage2[5][22] , \intermediateWiresStage2[5][21] , \intermediateWiresStage2[5][20] , 
    \intermediateWiresStage2[5][19] , \intermediateWiresStage2[5][18] , \intermediateWiresStage2[5][17] , 
    \intermediateWiresStage2[5][16] , \intermediateWiresStage2[5][15] , \intermediateWiresStage2[5][14] , 
    \intermediateWiresStage2[5][13] , \intermediateWiresStage2[5][12] , uc_3376, 
    uc_3377, uc_3378, uc_3379, uc_3380, uc_3381, uc_3382, uc_3383, uc_3384, uc_3385, 
    uc_3386, uc_3387}));
CSAlike__3_1006 genblk4_2_parallelAdderStage3 (.carry ({uc_3111, uc_3112, uc_3113, 
    uc_3114, uc_3115, uc_3116, uc_3117, uc_3118, uc_3119, uc_3120, uc_3121, uc_3122, 
    uc_3123, uc_3124, \intermediateWiresStage3[5][49] , \intermediateWiresStage3[5][48] , 
    \intermediateWiresStage3[5][47] , \intermediateWiresStage3[5][46] , \intermediateWiresStage3[5][45] , 
    \intermediateWiresStage3[5][44] , \intermediateWiresStage3[5][43] , \intermediateWiresStage3[5][42] , 
    \intermediateWiresStage3[5][41] , \intermediateWiresStage3[5][40] , \intermediateWiresStage3[5][39] , 
    \intermediateWiresStage3[5][38] , \intermediateWiresStage3[5][37] , \intermediateWiresStage3[5][36] , 
    \intermediateWiresStage3[5][35] , \intermediateWiresStage3[5][34] , \intermediateWiresStage3[5][33] , 
    \intermediateWiresStage3[5][32] , \intermediateWiresStage3[5][31] , \intermediateWiresStage3[5][30] , 
    \intermediateWiresStage3[5][29] , \intermediateWiresStage3[5][28] , \intermediateWiresStage3[5][27] , 
    \intermediateWiresStage3[5][26] , \intermediateWiresStage3[5][25] , \intermediateWiresStage3[5][24] , 
    \intermediateWiresStage3[5][23] , \intermediateWiresStage3[5][22] , \intermediateWiresStage3[5][21] , 
    \intermediateWiresStage3[5][20] , \intermediateWiresStage3[5][19] , \intermediateWiresStage3[5][18] , 
    \intermediateWiresStage3[5][17] , uc_3125, uc_3126, uc_3127, uc_3128, uc_3129, 
    uc_3130, uc_3131, uc_3132, uc_3133, uc_3134, uc_3135, uc_3136, uc_3137, uc_3138, 
    uc_3139, uc_3140, uc_3141}), .result ({uc_3080, uc_3081, uc_3082, uc_3083, uc_3084, 
    uc_3085, uc_3086, uc_3087, uc_3088, uc_3089, uc_3090, uc_3091, uc_3092, uc_3093, 
    uc_3094, \intermediateWiresStage3[4][48] , \intermediateWiresStage3[4][47] , 
    \intermediateWiresStage3[4][46] , \intermediateWiresStage3[4][45] , \intermediateWiresStage3[4][44] , 
    \intermediateWiresStage3[4][43] , \intermediateWiresStage3[4][42] , \intermediateWiresStage3[4][41] , 
    \intermediateWiresStage3[4][40] , \intermediateWiresStage3[4][39] , \intermediateWiresStage3[4][38] , 
    \intermediateWiresStage3[4][37] , \intermediateWiresStage3[4][36] , \intermediateWiresStage3[4][35] , 
    \intermediateWiresStage3[4][34] , \intermediateWiresStage3[4][33] , \intermediateWiresStage3[4][32] , 
    \intermediateWiresStage3[4][31] , \intermediateWiresStage3[4][30] , \intermediateWiresStage3[4][29] , 
    \intermediateWiresStage3[4][28] , \intermediateWiresStage3[4][27] , \intermediateWiresStage3[4][26] , 
    \intermediateWiresStage3[4][25] , \intermediateWiresStage3[4][24] , \intermediateWiresStage3[4][23] , 
    \intermediateWiresStage3[4][22] , \intermediateWiresStage3[4][21] , \intermediateWiresStage3[4][20] , 
    \intermediateWiresStage3[4][19] , \intermediateWiresStage3[4][18] , \intermediateWiresStage3[4][17] , 
    \intermediateWiresStage3[4][16] , uc_3095, uc_3096, uc_3097, uc_3098, uc_3099, 
    uc_3100, uc_3101, uc_3102, uc_3103, uc_3104, uc_3105, uc_3106, uc_3107, uc_3108, 
    uc_3109, uc_3110}), .A ({1'b0 , uc_3142, uc_3143, uc_3144, uc_3145, uc_3146, 
    uc_3147, uc_3148, uc_3149, uc_3150, uc_3151, uc_3152, uc_3153, uc_3154, uc_3155, 
    uc_3156, \intermediateWiresStage2[6][47] , \intermediateWiresStage2[6][46] , 
    \intermediateWiresStage2[6][45] , \intermediateWiresStage2[6][44] , \intermediateWiresStage2[6][43] , 
    \intermediateWiresStage2[6][42] , \intermediateWiresStage2[6][41] , \intermediateWiresStage2[6][40] , 
    \intermediateWiresStage2[6][39] , \intermediateWiresStage2[6][38] , \intermediateWiresStage2[6][37] , 
    \intermediateWiresStage2[6][36] , \intermediateWiresStage2[6][35] , \intermediateWiresStage2[6][34] , 
    \intermediateWiresStage2[6][33] , \intermediateWiresStage2[6][32] , \intermediateWiresStage2[6][31] , 
    \intermediateWiresStage2[6][30] , \intermediateWiresStage2[6][29] , \intermediateWiresStage2[6][28] , 
    \intermediateWiresStage2[6][27] , \intermediateWiresStage2[6][26] , \intermediateWiresStage2[6][25] , 
    \intermediateWiresStage2[6][24] , \intermediateWiresStage2[6][23] , \intermediateWiresStage2[6][22] , 
    \intermediateWiresStage2[6][21] , \intermediateWiresStage2[6][20] , \intermediateWiresStage2[6][19] , 
    \intermediateWiresStage2[6][18] , \intermediateWiresStage2[6][17] , \intermediateWiresStage2[6][16] , 
    uc_3157, uc_3158, uc_3159, uc_3160, uc_3161, uc_3162, uc_3163, uc_3164, uc_3165, 
    uc_3166, uc_3167, uc_3168, uc_3169, uc_3170, uc_3171, uc_3172}), .B ({1'b0 , 
    uc_3173, uc_3174, uc_3175, uc_3176, uc_3177, uc_3178, uc_3179, uc_3180, uc_3181, 
    uc_3182, uc_3183, uc_3184, uc_3185, uc_3186, \intermediateWiresStage2[7][48] , 
    \intermediateWiresStage2[7][47] , \intermediateWiresStage2[7][46] , \intermediateWiresStage2[7][45] , 
    \intermediateWiresStage2[7][44] , \intermediateWiresStage2[7][43] , \intermediateWiresStage2[7][42] , 
    \intermediateWiresStage2[7][41] , \intermediateWiresStage2[7][40] , \intermediateWiresStage2[7][39] , 
    \intermediateWiresStage2[7][38] , \intermediateWiresStage2[7][37] , \intermediateWiresStage2[7][36] , 
    \intermediateWiresStage2[7][35] , \intermediateWiresStage2[7][34] , \intermediateWiresStage2[7][33] , 
    \intermediateWiresStage2[7][32] , \intermediateWiresStage2[7][31] , \intermediateWiresStage2[7][30] , 
    \intermediateWiresStage2[7][29] , \intermediateWiresStage2[7][28] , \intermediateWiresStage2[7][27] , 
    \intermediateWiresStage2[7][26] , \intermediateWiresStage2[7][25] , \intermediateWiresStage2[7][24] , 
    \intermediateWiresStage2[7][23] , \intermediateWiresStage2[7][22] , \intermediateWiresStage2[7][21] , 
    \intermediateWiresStage2[7][20] , \intermediateWiresStage2[7][19] , \intermediateWiresStage2[7][18] , 
    \intermediateWiresStage2[7][17] , \intermediateWiresStage2[7][16] , uc_3187, 
    uc_3188, uc_3189, uc_3190, uc_3191, uc_3192, uc_3193, uc_3194, uc_3195, uc_3196, 
    uc_3197, uc_3198, uc_3199, uc_3200, uc_3201, uc_3202}), .C ({1'b0 , uc_3203, 
    uc_3204, uc_3205, uc_3206, uc_3207, uc_3208, uc_3209, uc_3210, uc_3211, uc_3212, 
    uc_3213, uc_3214, uc_3215, uc_3216, \intermediateWiresStage2[8][48] , \intermediateWiresStage2[8][47] , 
    \intermediateWiresStage2[8][46] , \intermediateWiresStage2[8][45] , \intermediateWiresStage2[8][44] , 
    \intermediateWiresStage2[8][43] , \intermediateWiresStage2[8][42] , \intermediateWiresStage2[8][41] , 
    \intermediateWiresStage2[8][40] , \intermediateWiresStage2[8][39] , \intermediateWiresStage2[8][38] , 
    \intermediateWiresStage2[8][37] , \intermediateWiresStage2[8][36] , \intermediateWiresStage2[8][35] , 
    \intermediateWiresStage2[8][34] , \intermediateWiresStage2[8][33] , \intermediateWiresStage2[8][32] , 
    \intermediateWiresStage2[8][31] , \intermediateWiresStage2[8][30] , \intermediateWiresStage2[8][29] , 
    \intermediateWiresStage2[8][28] , \intermediateWiresStage2[8][27] , \intermediateWiresStage2[8][26] , 
    \intermediateWiresStage2[8][25] , \intermediateWiresStage2[8][24] , \intermediateWiresStage2[8][23] , 
    \intermediateWiresStage2[8][22] , \intermediateWiresStage2[8][21] , \intermediateWiresStage2[8][20] , 
    \intermediateWiresStage1[12][19] , normalizedWires[1170], uc_3217, uc_3218, uc_3219, 
    uc_3220, uc_3221, uc_3222, uc_3223, uc_3224, uc_3225, uc_3226, uc_3227, uc_3228, 
    uc_3229, uc_3230, uc_3231, uc_3232, uc_3233, uc_3234}));
CSAlike__3_753 genblk4_3_parallelAdderStage3 (.carry ({uc_2956, uc_2957, uc_2958, 
    uc_2959, uc_2960, uc_2961, \intermediateWiresStage3[7][57] , \intermediateWiresStage3[7][56] , 
    \intermediateWiresStage3[7][55] , \intermediateWiresStage3[7][54] , \intermediateWiresStage3[7][53] , 
    \intermediateWiresStage3[7][52] , \intermediateWiresStage3[7][51] , \intermediateWiresStage3[7][50] , 
    \intermediateWiresStage3[7][49] , \intermediateWiresStage3[7][48] , \intermediateWiresStage3[7][47] , 
    \intermediateWiresStage3[7][46] , \intermediateWiresStage3[7][45] , \intermediateWiresStage3[7][44] , 
    \intermediateWiresStage3[7][43] , \intermediateWiresStage3[7][42] , \intermediateWiresStage3[7][41] , 
    \intermediateWiresStage3[7][40] , \intermediateWiresStage3[7][39] , \intermediateWiresStage3[7][38] , 
    \intermediateWiresStage3[7][37] , \intermediateWiresStage3[7][36] , \intermediateWiresStage3[7][35] , 
    \intermediateWiresStage3[7][34] , \intermediateWiresStage3[7][33] , \intermediateWiresStage3[7][32] , 
    \intermediateWiresStage3[7][31] , \intermediateWiresStage3[7][30] , \intermediateWiresStage3[7][29] , 
    \intermediateWiresStage3[7][28] , \intermediateWiresStage3[7][27] , \intermediateWiresStage3[7][26] , 
    \intermediateWiresStage3[7][25] , \intermediateWiresStage3[7][24] , uc_2962, 
    uc_2963, uc_2964, uc_2965, uc_2966, uc_2967, uc_2968, uc_2969, uc_2970, uc_2971, 
    uc_2972, uc_2973, uc_2974, uc_2975, uc_2976, uc_2977, uc_2978, uc_2979, uc_2980, 
    uc_2981, uc_2982, uc_2983, uc_2984, uc_2985}), .result ({uc_2926, uc_2927, uc_2928, 
    uc_2929, uc_2930, uc_2931, uc_2932, \intermediateWiresStage3[6][56] , \intermediateWiresStage3[6][55] , 
    \intermediateWiresStage3[6][54] , \intermediateWiresStage3[6][53] , \intermediateWiresStage3[6][52] , 
    \intermediateWiresStage3[6][51] , \intermediateWiresStage3[6][50] , \intermediateWiresStage3[6][49] , 
    \intermediateWiresStage3[6][48] , \intermediateWiresStage3[6][47] , \intermediateWiresStage3[6][46] , 
    \intermediateWiresStage3[6][45] , \intermediateWiresStage3[6][44] , \intermediateWiresStage3[6][43] , 
    \intermediateWiresStage3[6][42] , \intermediateWiresStage3[6][41] , \intermediateWiresStage3[6][40] , 
    \intermediateWiresStage3[6][39] , \intermediateWiresStage3[6][38] , \intermediateWiresStage3[6][37] , 
    \intermediateWiresStage3[6][36] , \intermediateWiresStage3[6][35] , \intermediateWiresStage3[6][34] , 
    \intermediateWiresStage3[6][33] , \intermediateWiresStage3[6][32] , \intermediateWiresStage3[6][31] , 
    \intermediateWiresStage3[6][30] , \intermediateWiresStage3[6][29] , \intermediateWiresStage3[6][28] , 
    \intermediateWiresStage3[6][27] , \intermediateWiresStage3[6][26] , \intermediateWiresStage3[6][25] , 
    \intermediateWiresStage3[6][24] , \intermediateWiresStage3[6][23] , uc_2933, 
    uc_2934, uc_2935, uc_2936, uc_2937, uc_2938, uc_2939, uc_2940, uc_2941, uc_2942, 
    uc_2943, uc_2944, uc_2945, uc_2946, uc_2947, uc_2948, uc_2949, uc_2950, uc_2951, 
    uc_2952, uc_2953, uc_2954, uc_2955}), .A ({1'b0 , uc_2986, uc_2987, uc_2988, 
    uc_2989, uc_2990, uc_2991, uc_2992, uc_2993, uc_2994, uc_2995, uc_2996, \intermediateWiresStage2[9][51] , 
    \intermediateWiresStage2[9][50] , \intermediateWiresStage2[9][49] , \intermediateWiresStage2[9][48] , 
    \intermediateWiresStage2[9][47] , \intermediateWiresStage2[9][46] , \intermediateWiresStage2[9][45] , 
    \intermediateWiresStage2[9][44] , \intermediateWiresStage2[9][43] , \intermediateWiresStage2[9][42] , 
    \intermediateWiresStage2[9][41] , \intermediateWiresStage2[9][40] , \intermediateWiresStage2[9][39] , 
    \intermediateWiresStage2[9][38] , \intermediateWiresStage2[9][37] , \intermediateWiresStage2[9][36] , 
    \intermediateWiresStage2[9][35] , \intermediateWiresStage2[9][34] , \intermediateWiresStage2[9][33] , 
    \intermediateWiresStage2[9][32] , \intermediateWiresStage2[9][31] , \intermediateWiresStage2[9][30] , 
    \intermediateWiresStage2[9][29] , \intermediateWiresStage2[9][28] , \intermediateWiresStage2[9][27] , 
    \intermediateWiresStage2[9][26] , \intermediateWiresStage2[9][25] , \intermediateWiresStage2[9][24] , 
    \intermediateWiresStage2[9][23] , uc_2997, uc_2998, uc_2999, uc_3000, uc_3001, 
    uc_3002, uc_3003, uc_3004, uc_3005, uc_3006, uc_3007, uc_3008, uc_3009, uc_3010, 
    uc_3011, uc_3012, uc_3013, uc_3014, uc_3015, uc_3016, uc_3017, uc_3018, uc_3019})
    , .B ({1'b0 , uc_3020, uc_3021, uc_3022, uc_3023, uc_3024, uc_3025, \intermediateWiresStage2[10][56] , 
    \intermediateWiresStage2[10][55] , \intermediateWiresStage2[10][54] , \intermediateWiresStage2[10][53] , 
    \intermediateWiresStage2[10][52] , \intermediateWiresStage2[10][51] , \intermediateWiresStage2[10][50] , 
    \intermediateWiresStage2[10][49] , \intermediateWiresStage2[10][48] , \intermediateWiresStage2[10][47] , 
    \intermediateWiresStage2[10][46] , \intermediateWiresStage2[10][45] , \intermediateWiresStage2[10][44] , 
    \intermediateWiresStage2[10][43] , \intermediateWiresStage2[10][42] , \intermediateWiresStage2[10][41] , 
    \intermediateWiresStage2[10][40] , \intermediateWiresStage2[10][39] , \intermediateWiresStage2[10][38] , 
    \intermediateWiresStage2[10][37] , \intermediateWiresStage2[10][36] , \intermediateWiresStage2[10][35] , 
    \intermediateWiresStage2[10][34] , \intermediateWiresStage2[10][33] , \intermediateWiresStage2[10][32] , 
    \intermediateWiresStage2[10][31] , \intermediateWiresStage2[10][30] , \intermediateWiresStage2[10][29] , 
    \intermediateWiresStage2[10][28] , \intermediateWiresStage2[10][27] , \intermediateWiresStage2[10][26] , 
    \intermediateWiresStage2[10][25] , \intermediateWiresStage2[10][24] , \intermediateWiresStage1[15][23] , 
    uc_3026, uc_3027, uc_3028, uc_3029, uc_3030, uc_3031, uc_3032, uc_3033, uc_3034, 
    uc_3035, uc_3036, uc_3037, uc_3038, uc_3039, uc_3040, uc_3041, uc_3042, uc_3043, 
    uc_3044, uc_3045, uc_3046, uc_3047, uc_3048}), .C ({1'b0 , uc_3049, uc_3050, 
    uc_3051, uc_3052, uc_3053, uc_3054, \intermediateWiresStage2[11][56] , \intermediateWiresStage2[11][55] , 
    \intermediateWiresStage2[11][54] , \intermediateWiresStage2[11][53] , \intermediateWiresStage2[11][52] , 
    \intermediateWiresStage2[11][51] , \intermediateWiresStage2[11][50] , \intermediateWiresStage2[11][49] , 
    \intermediateWiresStage2[11][48] , \intermediateWiresStage2[11][47] , \intermediateWiresStage2[11][46] , 
    \intermediateWiresStage2[11][45] , \intermediateWiresStage2[11][44] , \intermediateWiresStage2[11][43] , 
    \intermediateWiresStage2[11][42] , \intermediateWiresStage2[11][41] , \intermediateWiresStage2[11][40] , 
    \intermediateWiresStage2[11][39] , \intermediateWiresStage2[11][38] , \intermediateWiresStage2[11][37] , 
    \intermediateWiresStage2[11][36] , \intermediateWiresStage2[11][35] , \intermediateWiresStage2[11][34] , 
    \intermediateWiresStage2[11][33] , \intermediateWiresStage2[11][32] , \intermediateWiresStage2[11][31] , 
    \intermediateWiresStage2[11][30] , \intermediateWiresStage2[11][29] , \intermediateWiresStage2[11][28] , 
    \intermediateWiresStage2[11][27] , \intermediateWiresStage2[11][26] , \intermediateWiresStage2[11][25] , 
    uc_3055, uc_3056, uc_3057, uc_3058, uc_3059, uc_3060, uc_3061, uc_3062, uc_3063, 
    uc_3064, uc_3065, uc_3066, uc_3067, uc_3068, uc_3069, uc_3070, uc_3071, uc_3072, 
    uc_3073, uc_3074, uc_3075, uc_3076, uc_3077, uc_3078, uc_3079}));
CSAlike__3_500 genblk4_4_parallelAdderStage3 (.carry ({uc_2796, uc_2797, \intermediateWiresStage3[9][61] , 
    \intermediateWiresStage3[9][60] , \intermediateWiresStage3[9][59] , \intermediateWiresStage3[9][58] , 
    \intermediateWiresStage3[9][57] , \intermediateWiresStage3[9][56] , \intermediateWiresStage3[9][55] , 
    \intermediateWiresStage3[9][54] , \intermediateWiresStage3[9][53] , \intermediateWiresStage3[9][52] , 
    \intermediateWiresStage3[9][51] , \intermediateWiresStage3[9][50] , \intermediateWiresStage3[9][49] , 
    \intermediateWiresStage3[9][48] , \intermediateWiresStage3[9][47] , \intermediateWiresStage3[9][46] , 
    \intermediateWiresStage3[9][45] , \intermediateWiresStage3[9][44] , \intermediateWiresStage3[9][43] , 
    \intermediateWiresStage3[9][42] , \intermediateWiresStage3[9][41] , \intermediateWiresStage3[9][40] , 
    \intermediateWiresStage3[9][39] , \intermediateWiresStage3[9][38] , \intermediateWiresStage3[9][37] , 
    \intermediateWiresStage3[9][36] , \intermediateWiresStage3[9][35] , \intermediateWiresStage3[9][34] , 
    \intermediateWiresStage3[9][33] , \intermediateWiresStage3[9][32] , \intermediateWiresStage3[9][31] , 
    uc_2798, uc_2799, uc_2800, uc_2801, uc_2802, uc_2803, uc_2804, uc_2805, uc_2806, 
    uc_2807, uc_2808, uc_2809, uc_2810, uc_2811, uc_2812, uc_2813, uc_2814, uc_2815, 
    uc_2816, uc_2817, uc_2818, uc_2819, uc_2820, uc_2821, uc_2822, uc_2823, uc_2824, 
    uc_2825, uc_2826, uc_2827, uc_2828}), .result ({uc_2763, uc_2764, uc_2765, \intermediateWiresStage3[8][60] , 
    \intermediateWiresStage3[8][59] , \intermediateWiresStage3[8][58] , \intermediateWiresStage3[8][57] , 
    \intermediateWiresStage3[8][56] , \intermediateWiresStage3[8][55] , \intermediateWiresStage3[8][54] , 
    \intermediateWiresStage3[8][53] , \intermediateWiresStage3[8][52] , \intermediateWiresStage3[8][51] , 
    \intermediateWiresStage3[8][50] , \intermediateWiresStage3[8][49] , \intermediateWiresStage3[8][48] , 
    \intermediateWiresStage3[8][47] , \intermediateWiresStage3[8][46] , \intermediateWiresStage3[8][45] , 
    \intermediateWiresStage3[8][44] , \intermediateWiresStage3[8][43] , \intermediateWiresStage3[8][42] , 
    \intermediateWiresStage3[8][41] , \intermediateWiresStage3[8][40] , \intermediateWiresStage3[8][39] , 
    \intermediateWiresStage3[8][38] , \intermediateWiresStage3[8][37] , \intermediateWiresStage3[8][36] , 
    \intermediateWiresStage3[8][35] , \intermediateWiresStage3[8][34] , \intermediateWiresStage3[8][33] , 
    \intermediateWiresStage3[8][32] , \intermediateWiresStage3[8][31] , \intermediateWiresStage3[8][30] , 
    uc_2766, uc_2767, uc_2768, uc_2769, uc_2770, uc_2771, uc_2772, uc_2773, uc_2774, 
    uc_2775, uc_2776, uc_2777, uc_2778, uc_2779, uc_2780, uc_2781, uc_2782, uc_2783, 
    uc_2784, uc_2785, uc_2786, uc_2787, uc_2788, uc_2789, uc_2790, uc_2791, uc_2792, 
    uc_2793, uc_2794, uc_2795}), .A ({1'b0 , uc_2829, uc_2830, normalizedWires[1980], 
    \intermediateWiresStage2[12][59] , \intermediateWiresStage2[12][58] , \intermediateWiresStage2[12][57] , 
    \intermediateWiresStage2[12][56] , \intermediateWiresStage2[12][55] , \intermediateWiresStage2[12][54] , 
    \intermediateWiresStage2[12][53] , \intermediateWiresStage2[12][52] , \intermediateWiresStage2[12][51] , 
    \intermediateWiresStage2[12][50] , \intermediateWiresStage2[12][49] , \intermediateWiresStage2[12][48] , 
    \intermediateWiresStage2[12][47] , \intermediateWiresStage2[12][46] , \intermediateWiresStage2[12][45] , 
    \intermediateWiresStage2[12][44] , \intermediateWiresStage2[12][43] , \intermediateWiresStage2[12][42] , 
    \intermediateWiresStage2[12][41] , \intermediateWiresStage2[12][40] , \intermediateWiresStage2[12][39] , 
    \intermediateWiresStage2[12][38] , \intermediateWiresStage2[12][37] , \intermediateWiresStage2[12][36] , 
    \intermediateWiresStage2[12][35] , \intermediateWiresStage2[12][34] , \intermediateWiresStage2[12][33] , 
    \intermediateWiresStage2[12][32] , \intermediateWiresStage2[12][31] , \intermediateWiresStage2[12][30] , 
    uc_2831, uc_2832, uc_2833, uc_2834, uc_2835, uc_2836, uc_2837, uc_2838, uc_2839, 
    uc_2840, uc_2841, uc_2842, uc_2843, uc_2844, uc_2845, uc_2846, uc_2847, uc_2848, 
    uc_2849, uc_2850, uc_2851, uc_2852, uc_2853, uc_2854, uc_2855, uc_2856, uc_2857, 
    uc_2858, uc_2859, uc_2860}), .B ({1'b0 , uc_2861, uc_2862, \intermediateWiresStage2[13][60] , 
    \intermediateWiresStage2[13][59] , \intermediateWiresStage2[13][58] , \intermediateWiresStage2[13][57] , 
    \intermediateWiresStage2[13][56] , \intermediateWiresStage2[13][55] , \intermediateWiresStage2[13][54] , 
    \intermediateWiresStage2[13][53] , \intermediateWiresStage2[13][52] , \intermediateWiresStage2[13][51] , 
    \intermediateWiresStage2[13][50] , \intermediateWiresStage2[13][49] , \intermediateWiresStage2[13][48] , 
    \intermediateWiresStage2[13][47] , \intermediateWiresStage2[13][46] , \intermediateWiresStage2[13][45] , 
    \intermediateWiresStage2[13][44] , \intermediateWiresStage2[13][43] , \intermediateWiresStage2[13][42] , 
    \intermediateWiresStage2[13][41] , \intermediateWiresStage2[13][40] , \intermediateWiresStage2[13][39] , 
    \intermediateWiresStage2[13][38] , \intermediateWiresStage2[13][37] , \intermediateWiresStage2[13][36] , 
    \intermediateWiresStage2[13][35] , \intermediateWiresStage2[13][34] , \intermediateWiresStage2[13][33] , 
    \intermediateWiresStage2[13][32] , \intermediateWiresStage2[13][31] , \intermediateWiresStage2[13][30] , 
    uc_2863, uc_2864, uc_2865, uc_2866, uc_2867, uc_2868, uc_2869, uc_2870, uc_2871, 
    uc_2872, uc_2873, uc_2874, uc_2875, uc_2876, uc_2877, uc_2878, uc_2879, uc_2880, 
    uc_2881, uc_2882, uc_2883, uc_2884, uc_2885, uc_2886, uc_2887, uc_2888, uc_2889, 
    uc_2890, uc_2891, uc_2892}), .C ({1'b0 , uc_2893, uc_2894, normalizedWires[2044], 
    normalizedWires[2043], normalizedWires[2042], normalizedWires[2041], normalizedWires[2040], 
    normalizedWires[2039], normalizedWires[2038], normalizedWires[2037], normalizedWires[2036], 
    normalizedWires[2035], normalizedWires[2034], normalizedWires[2033], normalizedWires[2032], 
    normalizedWires[2031], normalizedWires[2030], normalizedWires[2029], normalizedWires[2028], 
    normalizedWires[2027], normalizedWires[2026], normalizedWires[2025], normalizedWires[2024], 
    normalizedWires[2023], normalizedWires[2022], normalizedWires[2021], normalizedWires[2020], 
    normalizedWires[2019], normalizedWires[2018], normalizedWires[2017], normalizedWires[2016], 
    normalizedWires[2015], uc_2895, uc_2896, uc_2897, uc_2898, uc_2899, uc_2900, 
    uc_2901, uc_2902, uc_2903, uc_2904, uc_2905, uc_2906, uc_2907, uc_2908, uc_2909, 
    uc_2910, uc_2911, uc_2912, uc_2913, uc_2914, uc_2915, uc_2916, uc_2917, uc_2918, 
    uc_2919, uc_2920, uc_2921, uc_2922, uc_2923, uc_2924, uc_2925}));
CSAlike__0_113 genblk3_0_parallelAdderStage2 (.carry ({uc_2633, uc_2634, uc_2635, 
    uc_2636, uc_2637, uc_2638, uc_2639, uc_2640, uc_2641, uc_2642, uc_2643, uc_2644, 
    uc_2645, uc_2646, uc_2647, uc_2648, uc_2649, uc_2650, uc_2651, uc_2652, uc_2653, 
    uc_2654, uc_2655, uc_2656, uc_2657, uc_2658, uc_2659, uc_2660, uc_2661, uc_2662, 
    \intermediateWiresStage2[1][33] , \intermediateWiresStage2[1][32] , \intermediateWiresStage2[1][31] , 
    \intermediateWiresStage2[1][30] , \intermediateWiresStage2[1][29] , \intermediateWiresStage2[1][28] , 
    \intermediateWiresStage2[1][27] , \intermediateWiresStage2[1][26] , \intermediateWiresStage2[1][25] , 
    \intermediateWiresStage2[1][24] , \intermediateWiresStage2[1][23] , \intermediateWiresStage2[1][22] , 
    \intermediateWiresStage2[1][21] , \intermediateWiresStage2[1][20] , \intermediateWiresStage2[1][19] , 
    \intermediateWiresStage2[1][18] , \intermediateWiresStage2[1][17] , \intermediateWiresStage2[1][16] , 
    \intermediateWiresStage2[1][15] , \intermediateWiresStage2[1][14] , \intermediateWiresStage2[1][13] , 
    \intermediateWiresStage2[1][12] , \intermediateWiresStage2[1][11] , \intermediateWiresStage2[1][10] , 
    \intermediateWiresStage2[1][9] , \intermediateWiresStage2[1][8] , \intermediateWiresStage2[1][7] , 
    \intermediateWiresStage2[1][6] , \intermediateWiresStage2[1][5] , \intermediateWiresStage2[1][4] , 
    \intermediateWiresStage2[1][3] , uc_2663, uc_2664, uc_2665}), .result ({uc_2600, 
    uc_2601, uc_2602, uc_2603, uc_2604, uc_2605, uc_2606, uc_2607, uc_2608, uc_2609, 
    uc_2610, uc_2611, uc_2612, uc_2613, uc_2614, uc_2615, uc_2616, uc_2617, uc_2618, 
    uc_2619, uc_2620, uc_2621, uc_2622, uc_2623, uc_2624, uc_2625, uc_2626, uc_2627, 
    uc_2628, uc_2629, uc_2630, \intermediateWiresStage2[0][32] , \intermediateWiresStage2[0][31] , 
    \intermediateWiresStage2[0][30] , \intermediateWiresStage2[0][29] , \intermediateWiresStage2[0][28] , 
    \intermediateWiresStage2[0][27] , \intermediateWiresStage2[0][26] , \intermediateWiresStage2[0][25] , 
    \intermediateWiresStage2[0][24] , \intermediateWiresStage2[0][23] , \intermediateWiresStage2[0][22] , 
    \intermediateWiresStage2[0][21] , \intermediateWiresStage2[0][20] , \intermediateWiresStage2[0][19] , 
    \intermediateWiresStage2[0][18] , \intermediateWiresStage2[0][17] , \intermediateWiresStage2[0][16] , 
    \intermediateWiresStage2[0][15] , \intermediateWiresStage2[0][14] , \intermediateWiresStage2[0][13] , 
    \intermediateWiresStage2[0][12] , \intermediateWiresStage2[0][11] , \intermediateWiresStage2[0][10] , 
    \intermediateWiresStage2[0][9] , \intermediateWiresStage2[0][8] , \intermediateWiresStage2[0][7] , 
    \intermediateWiresStage2[0][6] , \intermediateWiresStage2[0][5] , \intermediateWiresStage2[0][4] , 
    \intermediateWiresStage2[0][3] , Res[2], uc_2631, uc_2632}), .A ({1'b0 , uc_2666, 
    uc_2667, uc_2668, uc_2669, uc_2670, uc_2671, uc_2672, uc_2673, uc_2674, uc_2675, 
    uc_2676, uc_2677, uc_2678, uc_2679, uc_2680, uc_2681, uc_2682, uc_2683, uc_2684, 
    uc_2685, uc_2686, uc_2687, uc_2688, uc_2689, uc_2690, uc_2691, uc_2692, uc_2693, 
    uc_2694, uc_2695, normalizedWires[160], \intermediateWiresStage1[0][31] , \intermediateWiresStage1[0][30] , 
    \intermediateWiresStage1[0][29] , \intermediateWiresStage1[0][28] , \intermediateWiresStage1[0][27] , 
    \intermediateWiresStage1[0][26] , \intermediateWiresStage1[0][25] , \intermediateWiresStage1[0][24] , 
    \intermediateWiresStage1[0][23] , \intermediateWiresStage1[0][22] , \intermediateWiresStage1[0][21] , 
    \intermediateWiresStage1[0][20] , \intermediateWiresStage1[0][19] , \intermediateWiresStage1[0][18] , 
    \intermediateWiresStage1[0][17] , \intermediateWiresStage1[0][16] , \intermediateWiresStage1[0][15] , 
    \intermediateWiresStage1[0][14] , \intermediateWiresStage1[0][13] , \intermediateWiresStage1[0][12] , 
    \intermediateWiresStage1[0][11] , \intermediateWiresStage1[0][10] , \intermediateWiresStage1[0][9] , 
    \intermediateWiresStage1[0][8] , \intermediateWiresStage1[0][7] , \intermediateWiresStage1[0][6] , 
    \intermediateWiresStage1[0][5] , \intermediateWiresStage1[0][4] , \intermediateWiresStage1[0][3] , 
    \intermediateWiresStage1[0][2] , uc_2696, uc_2697}), .B ({1'b0 , uc_2698, uc_2699, 
    uc_2700, uc_2701, uc_2702, uc_2703, uc_2704, uc_2705, uc_2706, uc_2707, uc_2708, 
    uc_2709, uc_2710, uc_2711, uc_2712, uc_2713, uc_2714, uc_2715, uc_2716, uc_2717, 
    uc_2718, uc_2719, uc_2720, uc_2721, uc_2722, uc_2723, uc_2724, uc_2725, uc_2726, 
    uc_2727, \intermediateWiresStage1[1][32] , \intermediateWiresStage1[1][31] , 
    \intermediateWiresStage1[1][30] , \intermediateWiresStage1[1][29] , \intermediateWiresStage1[1][28] , 
    \intermediateWiresStage1[1][27] , \intermediateWiresStage1[1][26] , \intermediateWiresStage1[1][25] , 
    \intermediateWiresStage1[1][24] , \intermediateWiresStage1[1][23] , \intermediateWiresStage1[1][22] , 
    \intermediateWiresStage1[1][21] , \intermediateWiresStage1[1][20] , \intermediateWiresStage1[1][19] , 
    \intermediateWiresStage1[1][18] , \intermediateWiresStage1[1][17] , \intermediateWiresStage1[1][16] , 
    \intermediateWiresStage1[1][15] , \intermediateWiresStage1[1][14] , \intermediateWiresStage1[1][13] , 
    \intermediateWiresStage1[1][12] , \intermediateWiresStage1[1][11] , \intermediateWiresStage1[1][10] , 
    \intermediateWiresStage1[1][9] , \intermediateWiresStage1[1][8] , \intermediateWiresStage1[1][7] , 
    \intermediateWiresStage1[1][6] , \intermediateWiresStage1[1][5] , \intermediateWiresStage1[1][4] , 
    \intermediateWiresStage1[1][3] , \intermediateWiresStage1[1][2] , uc_2728, uc_2729})
    , .C ({1'b0 , uc_2730, uc_2731, uc_2732, uc_2733, uc_2734, uc_2735, uc_2736, 
    uc_2737, uc_2738, uc_2739, uc_2740, uc_2741, uc_2742, uc_2743, uc_2744, uc_2745, 
    uc_2746, uc_2747, uc_2748, uc_2749, uc_2750, uc_2751, uc_2752, uc_2753, uc_2754, 
    uc_2755, uc_2756, uc_2757, uc_2758, uc_2759, \intermediateWiresStage1[2][32] , 
    \intermediateWiresStage1[2][31] , \intermediateWiresStage1[2][30] , \intermediateWiresStage1[2][29] , 
    \intermediateWiresStage1[2][28] , \intermediateWiresStage1[2][27] , \intermediateWiresStage1[2][26] , 
    \intermediateWiresStage1[2][25] , \intermediateWiresStage1[2][24] , \intermediateWiresStage1[2][23] , 
    \intermediateWiresStage1[2][22] , \intermediateWiresStage1[2][21] , \intermediateWiresStage1[2][20] , 
    \intermediateWiresStage1[2][19] , \intermediateWiresStage1[2][18] , \intermediateWiresStage1[2][17] , 
    \intermediateWiresStage1[2][16] , \intermediateWiresStage1[2][15] , \intermediateWiresStage1[2][14] , 
    \intermediateWiresStage1[2][13] , \intermediateWiresStage1[2][12] , \intermediateWiresStage1[2][11] , 
    \intermediateWiresStage1[2][10] , \intermediateWiresStage1[2][9] , \intermediateWiresStage1[2][8] , 
    \intermediateWiresStage1[2][7] , \intermediateWiresStage1[2][6] , \intermediateWiresStage1[2][5] , 
    \intermediateWiresStage1[2][4] , normalizedWires[195], uc_2760, uc_2761, uc_2762}));
CSAlike__2_1765 genblk3_1_parallelAdderStage2 (.carry ({uc_2474, uc_2475, uc_2476, 
    uc_2477, uc_2478, uc_2479, uc_2480, uc_2481, uc_2482, uc_2483, uc_2484, uc_2485, 
    uc_2486, uc_2487, uc_2488, uc_2489, uc_2490, uc_2491, uc_2492, uc_2493, uc_2494, 
    uc_2495, uc_2496, uc_2497, \intermediateWiresStage2[3][39] , \intermediateWiresStage2[3][38] , 
    \intermediateWiresStage2[3][37] , \intermediateWiresStage2[3][36] , \intermediateWiresStage2[3][35] , 
    \intermediateWiresStage2[3][34] , \intermediateWiresStage2[3][33] , \intermediateWiresStage2[3][32] , 
    \intermediateWiresStage2[3][31] , \intermediateWiresStage2[3][30] , \intermediateWiresStage2[3][29] , 
    \intermediateWiresStage2[3][28] , \intermediateWiresStage2[3][27] , \intermediateWiresStage2[3][26] , 
    \intermediateWiresStage2[3][25] , \intermediateWiresStage2[3][24] , \intermediateWiresStage2[3][23] , 
    \intermediateWiresStage2[3][22] , \intermediateWiresStage2[3][21] , \intermediateWiresStage2[3][20] , 
    \intermediateWiresStage2[3][19] , \intermediateWiresStage2[3][18] , \intermediateWiresStage2[3][17] , 
    \intermediateWiresStage2[3][16] , \intermediateWiresStage2[3][15] , \intermediateWiresStage2[3][14] , 
    \intermediateWiresStage2[3][13] , \intermediateWiresStage2[3][12] , \intermediateWiresStage2[3][11] , 
    \intermediateWiresStage2[3][10] , \intermediateWiresStage2[3][9] , \intermediateWiresStage2[3][8] , 
    \intermediateWiresStage2[3][7] , uc_2498, uc_2499, uc_2500, uc_2501, uc_2502, 
    uc_2503, uc_2504}), .result ({uc_2443, uc_2444, uc_2445, uc_2446, uc_2447, uc_2448, 
    uc_2449, uc_2450, uc_2451, uc_2452, uc_2453, uc_2454, uc_2455, uc_2456, uc_2457, 
    uc_2458, uc_2459, uc_2460, uc_2461, uc_2462, uc_2463, uc_2464, uc_2465, uc_2466, 
    uc_2467, \intermediateWiresStage2[2][38] , \intermediateWiresStage2[2][37] , 
    \intermediateWiresStage2[2][36] , \intermediateWiresStage2[2][35] , \intermediateWiresStage2[2][34] , 
    \intermediateWiresStage2[2][33] , \intermediateWiresStage2[2][32] , \intermediateWiresStage2[2][31] , 
    \intermediateWiresStage2[2][30] , \intermediateWiresStage2[2][29] , \intermediateWiresStage2[2][28] , 
    \intermediateWiresStage2[2][27] , \intermediateWiresStage2[2][26] , \intermediateWiresStage2[2][25] , 
    \intermediateWiresStage2[2][24] , \intermediateWiresStage2[2][23] , \intermediateWiresStage2[2][22] , 
    \intermediateWiresStage2[2][21] , \intermediateWiresStage2[2][20] , \intermediateWiresStage2[2][19] , 
    \intermediateWiresStage2[2][18] , \intermediateWiresStage2[2][17] , \intermediateWiresStage2[2][16] , 
    \intermediateWiresStage2[2][15] , \intermediateWiresStage2[2][14] , \intermediateWiresStage2[2][13] , 
    \intermediateWiresStage2[2][12] , \intermediateWiresStage2[2][11] , \intermediateWiresStage2[2][10] , 
    \intermediateWiresStage2[2][9] , \intermediateWiresStage2[2][8] , \intermediateWiresStage2[2][7] , 
    \intermediateWiresStage2[2][6] , uc_2468, uc_2469, uc_2470, uc_2471, uc_2472, 
    uc_2473}), .A ({1'b0 , uc_2505, uc_2506, uc_2507, uc_2508, uc_2509, uc_2510, 
    uc_2511, uc_2512, uc_2513, uc_2514, uc_2515, uc_2516, uc_2517, uc_2518, uc_2519, 
    uc_2520, uc_2521, uc_2522, uc_2523, uc_2524, uc_2525, uc_2526, uc_2527, uc_2528, 
    uc_2529, uc_2530, uc_2531, \intermediateWiresStage1[3][35] , \intermediateWiresStage1[3][34] , 
    \intermediateWiresStage1[3][33] , \intermediateWiresStage1[3][32] , \intermediateWiresStage1[3][31] , 
    \intermediateWiresStage1[3][30] , \intermediateWiresStage1[3][29] , \intermediateWiresStage1[3][28] , 
    \intermediateWiresStage1[3][27] , \intermediateWiresStage1[3][26] , \intermediateWiresStage1[3][25] , 
    \intermediateWiresStage1[3][24] , \intermediateWiresStage1[3][23] , \intermediateWiresStage1[3][22] , 
    \intermediateWiresStage1[3][21] , \intermediateWiresStage1[3][20] , \intermediateWiresStage1[3][19] , 
    \intermediateWiresStage1[3][18] , \intermediateWiresStage1[3][17] , \intermediateWiresStage1[3][16] , 
    \intermediateWiresStage1[3][15] , \intermediateWiresStage1[3][14] , \intermediateWiresStage1[3][13] , 
    \intermediateWiresStage1[3][12] , \intermediateWiresStage1[3][11] , \intermediateWiresStage1[3][10] , 
    \intermediateWiresStage1[3][9] , \intermediateWiresStage1[3][8] , \intermediateWiresStage1[3][7] , 
    \intermediateWiresStage1[3][6] , uc_2532, uc_2533, uc_2534, uc_2535, uc_2536, 
    uc_2537}), .B ({1'b0 , uc_2538, uc_2539, uc_2540, uc_2541, uc_2542, uc_2543, 
    uc_2544, uc_2545, uc_2546, uc_2547, uc_2548, uc_2549, uc_2550, uc_2551, uc_2552, 
    uc_2553, uc_2554, uc_2555, uc_2556, uc_2557, uc_2558, uc_2559, uc_2560, uc_2561, 
    normalizedWires[550], \intermediateWiresStage1[4][37] , \intermediateWiresStage1[4][36] , 
    \intermediateWiresStage1[4][35] , \intermediateWiresStage1[4][34] , \intermediateWiresStage1[4][33] , 
    \intermediateWiresStage1[4][32] , \intermediateWiresStage1[4][31] , \intermediateWiresStage1[4][30] , 
    \intermediateWiresStage1[4][29] , \intermediateWiresStage1[4][28] , \intermediateWiresStage1[4][27] , 
    \intermediateWiresStage1[4][26] , \intermediateWiresStage1[4][25] , \intermediateWiresStage1[4][24] , 
    \intermediateWiresStage1[4][23] , \intermediateWiresStage1[4][22] , \intermediateWiresStage1[4][21] , 
    \intermediateWiresStage1[4][20] , \intermediateWiresStage1[4][19] , \intermediateWiresStage1[4][18] , 
    \intermediateWiresStage1[4][17] , \intermediateWiresStage1[4][16] , \intermediateWiresStage1[4][15] , 
    \intermediateWiresStage1[4][14] , \intermediateWiresStage1[4][13] , \intermediateWiresStage1[4][12] , 
    \intermediateWiresStage1[4][11] , \intermediateWiresStage1[4][10] , \intermediateWiresStage1[4][9] , 
    \intermediateWiresStage1[4][8] , \intermediateWiresStage1[4][7] , normalizedWires[390], 
    uc_2562, uc_2563, uc_2564, uc_2565, uc_2566, uc_2567}), .C ({1'b0 , uc_2568, 
    uc_2569, uc_2570, uc_2571, uc_2572, uc_2573, uc_2574, uc_2575, uc_2576, uc_2577, 
    uc_2578, uc_2579, uc_2580, uc_2581, uc_2582, uc_2583, uc_2584, uc_2585, uc_2586, 
    uc_2587, uc_2588, uc_2589, uc_2590, uc_2591, \intermediateWiresStage1[5][38] , 
    \intermediateWiresStage1[5][37] , \intermediateWiresStage1[5][36] , \intermediateWiresStage1[5][35] , 
    \intermediateWiresStage1[5][34] , \intermediateWiresStage1[5][33] , \intermediateWiresStage1[5][32] , 
    \intermediateWiresStage1[5][31] , \intermediateWiresStage1[5][30] , \intermediateWiresStage1[5][29] , 
    \intermediateWiresStage1[5][28] , \intermediateWiresStage1[5][27] , \intermediateWiresStage1[5][26] , 
    \intermediateWiresStage1[5][25] , \intermediateWiresStage1[5][24] , \intermediateWiresStage1[5][23] , 
    \intermediateWiresStage1[5][22] , \intermediateWiresStage1[5][21] , \intermediateWiresStage1[5][20] , 
    \intermediateWiresStage1[5][19] , \intermediateWiresStage1[5][18] , \intermediateWiresStage1[5][17] , 
    \intermediateWiresStage1[5][16] , \intermediateWiresStage1[5][15] , \intermediateWiresStage1[5][14] , 
    \intermediateWiresStage1[5][13] , \intermediateWiresStage1[5][12] , \intermediateWiresStage1[5][11] , 
    \intermediateWiresStage1[5][10] , \intermediateWiresStage1[5][9] , \intermediateWiresStage1[5][8] , 
    uc_2592, uc_2593, uc_2594, uc_2595, uc_2596, uc_2597, uc_2598, uc_2599}));
CSAlike__2_1512 genblk3_2_parallelAdderStage2 (.carry ({uc_2313, uc_2314, uc_2315, 
    uc_2316, uc_2317, uc_2318, uc_2319, uc_2320, uc_2321, uc_2322, uc_2323, uc_2324, 
    uc_2325, uc_2326, uc_2327, uc_2328, uc_2329, uc_2330, uc_2331, uc_2332, uc_2333, 
    \intermediateWiresStage2[5][42] , \intermediateWiresStage2[5][41] , \intermediateWiresStage2[5][40] , 
    \intermediateWiresStage2[5][39] , \intermediateWiresStage2[5][38] , \intermediateWiresStage2[5][37] , 
    \intermediateWiresStage2[5][36] , \intermediateWiresStage2[5][35] , \intermediateWiresStage2[5][34] , 
    \intermediateWiresStage2[5][33] , \intermediateWiresStage2[5][32] , \intermediateWiresStage2[5][31] , 
    \intermediateWiresStage2[5][30] , \intermediateWiresStage2[5][29] , \intermediateWiresStage2[5][28] , 
    \intermediateWiresStage2[5][27] , \intermediateWiresStage2[5][26] , \intermediateWiresStage2[5][25] , 
    \intermediateWiresStage2[5][24] , \intermediateWiresStage2[5][23] , \intermediateWiresStage2[5][22] , 
    \intermediateWiresStage2[5][21] , \intermediateWiresStage2[5][20] , \intermediateWiresStage2[5][19] , 
    \intermediateWiresStage2[5][18] , \intermediateWiresStage2[5][17] , \intermediateWiresStage2[5][16] , 
    \intermediateWiresStage2[5][15] , \intermediateWiresStage2[5][14] , \intermediateWiresStage2[5][13] , 
    \intermediateWiresStage2[5][12] , uc_2334, uc_2335, uc_2336, uc_2337, uc_2338, 
    uc_2339, uc_2340, uc_2341, uc_2342, uc_2343, uc_2344, uc_2345}), .result ({uc_2280, 
    uc_2281, uc_2282, uc_2283, uc_2284, uc_2285, uc_2286, uc_2287, uc_2288, uc_2289, 
    uc_2290, uc_2291, uc_2292, uc_2293, uc_2294, uc_2295, uc_2296, uc_2297, uc_2298, 
    uc_2299, uc_2300, uc_2301, \intermediateWiresStage2[4][41] , \intermediateWiresStage2[4][40] , 
    \intermediateWiresStage2[4][39] , \intermediateWiresStage2[4][38] , \intermediateWiresStage2[4][37] , 
    \intermediateWiresStage2[4][36] , \intermediateWiresStage2[4][35] , \intermediateWiresStage2[4][34] , 
    \intermediateWiresStage2[4][33] , \intermediateWiresStage2[4][32] , \intermediateWiresStage2[4][31] , 
    \intermediateWiresStage2[4][30] , \intermediateWiresStage2[4][29] , \intermediateWiresStage2[4][28] , 
    \intermediateWiresStage2[4][27] , \intermediateWiresStage2[4][26] , \intermediateWiresStage2[4][25] , 
    \intermediateWiresStage2[4][24] , \intermediateWiresStage2[4][23] , \intermediateWiresStage2[4][22] , 
    \intermediateWiresStage2[4][21] , \intermediateWiresStage2[4][20] , \intermediateWiresStage2[4][19] , 
    \intermediateWiresStage2[4][18] , \intermediateWiresStage2[4][17] , \intermediateWiresStage2[4][16] , 
    \intermediateWiresStage2[4][15] , \intermediateWiresStage2[4][14] , \intermediateWiresStage2[4][13] , 
    \intermediateWiresStage2[4][12] , \intermediateWiresStage2[4][11] , uc_2302, 
    uc_2303, uc_2304, uc_2305, uc_2306, uc_2307, uc_2308, uc_2309, uc_2310, uc_2311, 
    uc_2312}), .A ({1'b0 , uc_2346, uc_2347, uc_2348, uc_2349, uc_2350, uc_2351, 
    uc_2352, uc_2353, uc_2354, uc_2355, uc_2356, uc_2357, uc_2358, uc_2359, uc_2360, 
    uc_2361, uc_2362, uc_2363, uc_2364, uc_2365, uc_2366, normalizedWires[745], \intermediateWiresStage1[6][40] , 
    \intermediateWiresStage1[6][39] , \intermediateWiresStage1[6][38] , \intermediateWiresStage1[6][37] , 
    \intermediateWiresStage1[6][36] , \intermediateWiresStage1[6][35] , \intermediateWiresStage1[6][34] , 
    \intermediateWiresStage1[6][33] , \intermediateWiresStage1[6][32] , \intermediateWiresStage1[6][31] , 
    \intermediateWiresStage1[6][30] , \intermediateWiresStage1[6][29] , \intermediateWiresStage1[6][28] , 
    \intermediateWiresStage1[6][27] , \intermediateWiresStage1[6][26] , \intermediateWiresStage1[6][25] , 
    \intermediateWiresStage1[6][24] , \intermediateWiresStage1[6][23] , \intermediateWiresStage1[6][22] , 
    \intermediateWiresStage1[6][21] , \intermediateWiresStage1[6][20] , \intermediateWiresStage1[6][19] , 
    \intermediateWiresStage1[6][18] , \intermediateWiresStage1[6][17] , \intermediateWiresStage1[6][16] , 
    \intermediateWiresStage1[6][15] , \intermediateWiresStage1[6][14] , \intermediateWiresStage1[6][13] , 
    \intermediateWiresStage1[6][12] , \intermediateWiresStage1[6][11] , uc_2367, 
    uc_2368, uc_2369, uc_2370, uc_2371, uc_2372, uc_2373, uc_2374, uc_2375, uc_2376, 
    uc_2377}), .B ({1'b0 , uc_2378, uc_2379, uc_2380, uc_2381, uc_2382, uc_2383, 
    uc_2384, uc_2385, uc_2386, uc_2387, uc_2388, uc_2389, uc_2390, uc_2391, uc_2392, 
    uc_2393, uc_2394, uc_2395, uc_2396, uc_2397, uc_2398, \intermediateWiresStage1[7][41] , 
    \intermediateWiresStage1[7][40] , \intermediateWiresStage1[7][39] , \intermediateWiresStage1[7][38] , 
    \intermediateWiresStage1[7][37] , \intermediateWiresStage1[7][36] , \intermediateWiresStage1[7][35] , 
    \intermediateWiresStage1[7][34] , \intermediateWiresStage1[7][33] , \intermediateWiresStage1[7][32] , 
    \intermediateWiresStage1[7][31] , \intermediateWiresStage1[7][30] , \intermediateWiresStage1[7][29] , 
    \intermediateWiresStage1[7][28] , \intermediateWiresStage1[7][27] , \intermediateWiresStage1[7][26] , 
    \intermediateWiresStage1[7][25] , \intermediateWiresStage1[7][24] , \intermediateWiresStage1[7][23] , 
    \intermediateWiresStage1[7][22] , \intermediateWiresStage1[7][21] , \intermediateWiresStage1[7][20] , 
    \intermediateWiresStage1[7][19] , \intermediateWiresStage1[7][18] , \intermediateWiresStage1[7][17] , 
    \intermediateWiresStage1[7][16] , \intermediateWiresStage1[7][15] , \intermediateWiresStage1[7][14] , 
    \intermediateWiresStage1[7][13] , \intermediateWiresStage1[7][12] , \intermediateWiresStage1[7][11] , 
    uc_2399, uc_2400, uc_2401, uc_2402, uc_2403, uc_2404, uc_2405, uc_2406, uc_2407, 
    uc_2408, uc_2409}), .C ({1'b0 , uc_2410, uc_2411, uc_2412, uc_2413, uc_2414, 
    uc_2415, uc_2416, uc_2417, uc_2418, uc_2419, uc_2420, uc_2421, uc_2422, uc_2423, 
    uc_2424, uc_2425, uc_2426, uc_2427, uc_2428, uc_2429, uc_2430, \intermediateWiresStage1[8][41] , 
    \intermediateWiresStage1[8][40] , \intermediateWiresStage1[8][39] , \intermediateWiresStage1[8][38] , 
    \intermediateWiresStage1[8][37] , \intermediateWiresStage1[8][36] , \intermediateWiresStage1[8][35] , 
    \intermediateWiresStage1[8][34] , \intermediateWiresStage1[8][33] , \intermediateWiresStage1[8][32] , 
    \intermediateWiresStage1[8][31] , \intermediateWiresStage1[8][30] , \intermediateWiresStage1[8][29] , 
    \intermediateWiresStage1[8][28] , \intermediateWiresStage1[8][27] , \intermediateWiresStage1[8][26] , 
    \intermediateWiresStage1[8][25] , \intermediateWiresStage1[8][24] , \intermediateWiresStage1[8][23] , 
    \intermediateWiresStage1[8][22] , \intermediateWiresStage1[8][21] , \intermediateWiresStage1[8][20] , 
    \intermediateWiresStage1[8][19] , \intermediateWiresStage1[8][18] , \intermediateWiresStage1[8][17] , 
    \intermediateWiresStage1[8][16] , \intermediateWiresStage1[8][15] , \intermediateWiresStage1[8][14] , 
    \intermediateWiresStage1[8][13] , normalizedWires[780], uc_2431, uc_2432, uc_2433, 
    uc_2434, uc_2435, uc_2436, uc_2437, uc_2438, uc_2439, uc_2440, uc_2441, uc_2442}));
CSAlike__2_1259 genblk3_3_parallelAdderStage2 (.carry ({uc_2154, uc_2155, uc_2156, 
    uc_2157, uc_2158, uc_2159, uc_2160, uc_2161, uc_2162, uc_2163, uc_2164, uc_2165, 
    uc_2166, uc_2167, uc_2168, \intermediateWiresStage2[7][48] , \intermediateWiresStage2[7][47] , 
    \intermediateWiresStage2[7][46] , \intermediateWiresStage2[7][45] , \intermediateWiresStage2[7][44] , 
    \intermediateWiresStage2[7][43] , \intermediateWiresStage2[7][42] , \intermediateWiresStage2[7][41] , 
    \intermediateWiresStage2[7][40] , \intermediateWiresStage2[7][39] , \intermediateWiresStage2[7][38] , 
    \intermediateWiresStage2[7][37] , \intermediateWiresStage2[7][36] , \intermediateWiresStage2[7][35] , 
    \intermediateWiresStage2[7][34] , \intermediateWiresStage2[7][33] , \intermediateWiresStage2[7][32] , 
    \intermediateWiresStage2[7][31] , \intermediateWiresStage2[7][30] , \intermediateWiresStage2[7][29] , 
    \intermediateWiresStage2[7][28] , \intermediateWiresStage2[7][27] , \intermediateWiresStage2[7][26] , 
    \intermediateWiresStage2[7][25] , \intermediateWiresStage2[7][24] , \intermediateWiresStage2[7][23] , 
    \intermediateWiresStage2[7][22] , \intermediateWiresStage2[7][21] , \intermediateWiresStage2[7][20] , 
    \intermediateWiresStage2[7][19] , \intermediateWiresStage2[7][18] , \intermediateWiresStage2[7][17] , 
    \intermediateWiresStage2[7][16] , uc_2169, uc_2170, uc_2171, uc_2172, uc_2173, 
    uc_2174, uc_2175, uc_2176, uc_2177, uc_2178, uc_2179, uc_2180, uc_2181, uc_2182, 
    uc_2183, uc_2184}), .result ({uc_2123, uc_2124, uc_2125, uc_2126, uc_2127, uc_2128, 
    uc_2129, uc_2130, uc_2131, uc_2132, uc_2133, uc_2134, uc_2135, uc_2136, uc_2137, 
    uc_2138, \intermediateWiresStage2[6][47] , \intermediateWiresStage2[6][46] , 
    \intermediateWiresStage2[6][45] , \intermediateWiresStage2[6][44] , \intermediateWiresStage2[6][43] , 
    \intermediateWiresStage2[6][42] , \intermediateWiresStage2[6][41] , \intermediateWiresStage2[6][40] , 
    \intermediateWiresStage2[6][39] , \intermediateWiresStage2[6][38] , \intermediateWiresStage2[6][37] , 
    \intermediateWiresStage2[6][36] , \intermediateWiresStage2[6][35] , \intermediateWiresStage2[6][34] , 
    \intermediateWiresStage2[6][33] , \intermediateWiresStage2[6][32] , \intermediateWiresStage2[6][31] , 
    \intermediateWiresStage2[6][30] , \intermediateWiresStage2[6][29] , \intermediateWiresStage2[6][28] , 
    \intermediateWiresStage2[6][27] , \intermediateWiresStage2[6][26] , \intermediateWiresStage2[6][25] , 
    \intermediateWiresStage2[6][24] , \intermediateWiresStage2[6][23] , \intermediateWiresStage2[6][22] , 
    \intermediateWiresStage2[6][21] , \intermediateWiresStage2[6][20] , \intermediateWiresStage2[6][19] , 
    \intermediateWiresStage2[6][18] , \intermediateWiresStage2[6][17] , \intermediateWiresStage2[6][16] , 
    \intermediateWiresStage2[6][15] , uc_2139, uc_2140, uc_2141, uc_2142, uc_2143, 
    uc_2144, uc_2145, uc_2146, uc_2147, uc_2148, uc_2149, uc_2150, uc_2151, uc_2152, 
    uc_2153}), .A ({1'b0 , uc_2185, uc_2186, uc_2187, uc_2188, uc_2189, uc_2190, 
    uc_2191, uc_2192, uc_2193, uc_2194, uc_2195, uc_2196, uc_2197, uc_2198, uc_2199, 
    uc_2200, uc_2201, uc_2202, \intermediateWiresStage1[9][44] , \intermediateWiresStage1[9][43] , 
    \intermediateWiresStage1[9][42] , \intermediateWiresStage1[9][41] , \intermediateWiresStage1[9][40] , 
    \intermediateWiresStage1[9][39] , \intermediateWiresStage1[9][38] , \intermediateWiresStage1[9][37] , 
    \intermediateWiresStage1[9][36] , \intermediateWiresStage1[9][35] , \intermediateWiresStage1[9][34] , 
    \intermediateWiresStage1[9][33] , \intermediateWiresStage1[9][32] , \intermediateWiresStage1[9][31] , 
    \intermediateWiresStage1[9][30] , \intermediateWiresStage1[9][29] , \intermediateWiresStage1[9][28] , 
    \intermediateWiresStage1[9][27] , \intermediateWiresStage1[9][26] , \intermediateWiresStage1[9][25] , 
    \intermediateWiresStage1[9][24] , \intermediateWiresStage1[9][23] , \intermediateWiresStage1[9][22] , 
    \intermediateWiresStage1[9][21] , \intermediateWiresStage1[9][20] , \intermediateWiresStage1[9][19] , 
    \intermediateWiresStage1[9][18] , \intermediateWiresStage1[9][17] , \intermediateWiresStage1[9][16] , 
    \intermediateWiresStage1[9][15] , uc_2203, uc_2204, uc_2205, uc_2206, uc_2207, 
    uc_2208, uc_2209, uc_2210, uc_2211, uc_2212, uc_2213, uc_2214, uc_2215, uc_2216, 
    uc_2217}), .B ({1'b0 , uc_2218, uc_2219, uc_2220, uc_2221, uc_2222, uc_2223, 
    uc_2224, uc_2225, uc_2226, uc_2227, uc_2228, uc_2229, uc_2230, uc_2231, uc_2232, 
    normalizedWires[1135], \intermediateWiresStage1[10][46] , \intermediateWiresStage1[10][45] , 
    \intermediateWiresStage1[10][44] , \intermediateWiresStage1[10][43] , \intermediateWiresStage1[10][42] , 
    \intermediateWiresStage1[10][41] , \intermediateWiresStage1[10][40] , \intermediateWiresStage1[10][39] , 
    \intermediateWiresStage1[10][38] , \intermediateWiresStage1[10][37] , \intermediateWiresStage1[10][36] , 
    \intermediateWiresStage1[10][35] , \intermediateWiresStage1[10][34] , \intermediateWiresStage1[10][33] , 
    \intermediateWiresStage1[10][32] , \intermediateWiresStage1[10][31] , \intermediateWiresStage1[10][30] , 
    \intermediateWiresStage1[10][29] , \intermediateWiresStage1[10][28] , \intermediateWiresStage1[10][27] , 
    \intermediateWiresStage1[10][26] , \intermediateWiresStage1[10][25] , \intermediateWiresStage1[10][24] , 
    \intermediateWiresStage1[10][23] , \intermediateWiresStage1[10][22] , \intermediateWiresStage1[10][21] , 
    \intermediateWiresStage1[10][20] , \intermediateWiresStage1[10][19] , \intermediateWiresStage1[10][18] , 
    \intermediateWiresStage1[10][17] , \intermediateWiresStage1[10][16] , normalizedWires[975], 
    uc_2233, uc_2234, uc_2235, uc_2236, uc_2237, uc_2238, uc_2239, uc_2240, uc_2241, 
    uc_2242, uc_2243, uc_2244, uc_2245, uc_2246, uc_2247}), .C ({1'b0 , uc_2248, 
    uc_2249, uc_2250, uc_2251, uc_2252, uc_2253, uc_2254, uc_2255, uc_2256, uc_2257, 
    uc_2258, uc_2259, uc_2260, uc_2261, uc_2262, \intermediateWiresStage1[11][47] , 
    \intermediateWiresStage1[11][46] , \intermediateWiresStage1[11][45] , \intermediateWiresStage1[11][44] , 
    \intermediateWiresStage1[11][43] , \intermediateWiresStage1[11][42] , \intermediateWiresStage1[11][41] , 
    \intermediateWiresStage1[11][40] , \intermediateWiresStage1[11][39] , \intermediateWiresStage1[11][38] , 
    \intermediateWiresStage1[11][37] , \intermediateWiresStage1[11][36] , \intermediateWiresStage1[11][35] , 
    \intermediateWiresStage1[11][34] , \intermediateWiresStage1[11][33] , \intermediateWiresStage1[11][32] , 
    \intermediateWiresStage1[11][31] , \intermediateWiresStage1[11][30] , \intermediateWiresStage1[11][29] , 
    \intermediateWiresStage1[11][28] , \intermediateWiresStage1[11][27] , \intermediateWiresStage1[11][26] , 
    \intermediateWiresStage1[11][25] , \intermediateWiresStage1[11][24] , \intermediateWiresStage1[11][23] , 
    \intermediateWiresStage1[11][22] , \intermediateWiresStage1[11][21] , \intermediateWiresStage1[11][20] , 
    \intermediateWiresStage1[11][19] , \intermediateWiresStage1[11][18] , \intermediateWiresStage1[11][17] , 
    uc_2263, uc_2264, uc_2265, uc_2266, uc_2267, uc_2268, uc_2269, uc_2270, uc_2271, 
    uc_2272, uc_2273, uc_2274, uc_2275, uc_2276, uc_2277, uc_2278, uc_2279}));
CSAlike__2_1006 genblk3_4_parallelAdderStage2 (.carry ({uc_1993, uc_1994, uc_1995, 
    uc_1996, uc_1997, uc_1998, uc_1999, uc_2000, uc_2001, uc_2002, uc_2003, uc_2004, 
    \intermediateWiresStage2[9][51] , \intermediateWiresStage2[9][50] , \intermediateWiresStage2[9][49] , 
    \intermediateWiresStage2[9][48] , \intermediateWiresStage2[9][47] , \intermediateWiresStage2[9][46] , 
    \intermediateWiresStage2[9][45] , \intermediateWiresStage2[9][44] , \intermediateWiresStage2[9][43] , 
    \intermediateWiresStage2[9][42] , \intermediateWiresStage2[9][41] , \intermediateWiresStage2[9][40] , 
    \intermediateWiresStage2[9][39] , \intermediateWiresStage2[9][38] , \intermediateWiresStage2[9][37] , 
    \intermediateWiresStage2[9][36] , \intermediateWiresStage2[9][35] , \intermediateWiresStage2[9][34] , 
    \intermediateWiresStage2[9][33] , \intermediateWiresStage2[9][32] , \intermediateWiresStage2[9][31] , 
    \intermediateWiresStage2[9][30] , \intermediateWiresStage2[9][29] , \intermediateWiresStage2[9][28] , 
    \intermediateWiresStage2[9][27] , \intermediateWiresStage2[9][26] , \intermediateWiresStage2[9][25] , 
    \intermediateWiresStage2[9][24] , \intermediateWiresStage2[9][23] , \intermediateWiresStage2[9][22] , 
    \intermediateWiresStage2[9][21] , uc_2005, uc_2006, uc_2007, uc_2008, uc_2009, 
    uc_2010, uc_2011, uc_2012, uc_2013, uc_2014, uc_2015, uc_2016, uc_2017, uc_2018, 
    uc_2019, uc_2020, uc_2021, uc_2022, uc_2023, uc_2024, uc_2025}), .result ({uc_1960, 
    uc_1961, uc_1962, uc_1963, uc_1964, uc_1965, uc_1966, uc_1967, uc_1968, uc_1969, 
    uc_1970, uc_1971, uc_1972, \intermediateWiresStage2[8][50] , \intermediateWiresStage2[8][49] , 
    \intermediateWiresStage2[8][48] , \intermediateWiresStage2[8][47] , \intermediateWiresStage2[8][46] , 
    \intermediateWiresStage2[8][45] , \intermediateWiresStage2[8][44] , \intermediateWiresStage2[8][43] , 
    \intermediateWiresStage2[8][42] , \intermediateWiresStage2[8][41] , \intermediateWiresStage2[8][40] , 
    \intermediateWiresStage2[8][39] , \intermediateWiresStage2[8][38] , \intermediateWiresStage2[8][37] , 
    \intermediateWiresStage2[8][36] , \intermediateWiresStage2[8][35] , \intermediateWiresStage2[8][34] , 
    \intermediateWiresStage2[8][33] , \intermediateWiresStage2[8][32] , \intermediateWiresStage2[8][31] , 
    \intermediateWiresStage2[8][30] , \intermediateWiresStage2[8][29] , \intermediateWiresStage2[8][28] , 
    \intermediateWiresStage2[8][27] , \intermediateWiresStage2[8][26] , \intermediateWiresStage2[8][25] , 
    \intermediateWiresStage2[8][24] , \intermediateWiresStage2[8][23] , \intermediateWiresStage2[8][22] , 
    \intermediateWiresStage2[8][21] , \intermediateWiresStage2[8][20] , uc_1973, 
    uc_1974, uc_1975, uc_1976, uc_1977, uc_1978, uc_1979, uc_1980, uc_1981, uc_1982, 
    uc_1983, uc_1984, uc_1985, uc_1986, uc_1987, uc_1988, uc_1989, uc_1990, uc_1991, 
    uc_1992}), .A ({1'b0 , uc_2026, uc_2027, uc_2028, uc_2029, uc_2030, uc_2031, 
    uc_2032, uc_2033, uc_2034, uc_2035, uc_2036, uc_2037, normalizedWires[1330], 
    \intermediateWiresStage1[12][49] , \intermediateWiresStage1[12][48] , \intermediateWiresStage1[12][47] , 
    \intermediateWiresStage1[12][46] , \intermediateWiresStage1[12][45] , \intermediateWiresStage1[12][44] , 
    \intermediateWiresStage1[12][43] , \intermediateWiresStage1[12][42] , \intermediateWiresStage1[12][41] , 
    \intermediateWiresStage1[12][40] , \intermediateWiresStage1[12][39] , \intermediateWiresStage1[12][38] , 
    \intermediateWiresStage1[12][37] , \intermediateWiresStage1[12][36] , \intermediateWiresStage1[12][35] , 
    \intermediateWiresStage1[12][34] , \intermediateWiresStage1[12][33] , \intermediateWiresStage1[12][32] , 
    \intermediateWiresStage1[12][31] , \intermediateWiresStage1[12][30] , \intermediateWiresStage1[12][29] , 
    \intermediateWiresStage1[12][28] , \intermediateWiresStage1[12][27] , \intermediateWiresStage1[12][26] , 
    \intermediateWiresStage1[12][25] , \intermediateWiresStage1[12][24] , \intermediateWiresStage1[12][23] , 
    \intermediateWiresStage1[12][22] , \intermediateWiresStage1[12][21] , \intermediateWiresStage1[12][20] , 
    uc_2038, uc_2039, uc_2040, uc_2041, uc_2042, uc_2043, uc_2044, uc_2045, uc_2046, 
    uc_2047, uc_2048, uc_2049, uc_2050, uc_2051, uc_2052, uc_2053, uc_2054, uc_2055, 
    uc_2056, uc_2057}), .B ({1'b0 , uc_2058, uc_2059, uc_2060, uc_2061, uc_2062, 
    uc_2063, uc_2064, uc_2065, uc_2066, uc_2067, uc_2068, uc_2069, \intermediateWiresStage1[13][50] , 
    \intermediateWiresStage1[13][49] , \intermediateWiresStage1[13][48] , \intermediateWiresStage1[13][47] , 
    \intermediateWiresStage1[13][46] , \intermediateWiresStage1[13][45] , \intermediateWiresStage1[13][44] , 
    \intermediateWiresStage1[13][43] , \intermediateWiresStage1[13][42] , \intermediateWiresStage1[13][41] , 
    \intermediateWiresStage1[13][40] , \intermediateWiresStage1[13][39] , \intermediateWiresStage1[13][38] , 
    \intermediateWiresStage1[13][37] , \intermediateWiresStage1[13][36] , \intermediateWiresStage1[13][35] , 
    \intermediateWiresStage1[13][34] , \intermediateWiresStage1[13][33] , \intermediateWiresStage1[13][32] , 
    \intermediateWiresStage1[13][31] , \intermediateWiresStage1[13][30] , \intermediateWiresStage1[13][29] , 
    \intermediateWiresStage1[13][28] , \intermediateWiresStage1[13][27] , \intermediateWiresStage1[13][26] , 
    \intermediateWiresStage1[13][25] , \intermediateWiresStage1[13][24] , \intermediateWiresStage1[13][23] , 
    \intermediateWiresStage1[13][22] , \intermediateWiresStage1[13][21] , \intermediateWiresStage1[13][20] , 
    uc_2070, uc_2071, uc_2072, uc_2073, uc_2074, uc_2075, uc_2076, uc_2077, uc_2078, 
    uc_2079, uc_2080, uc_2081, uc_2082, uc_2083, uc_2084, uc_2085, uc_2086, uc_2087, 
    uc_2088, uc_2089}), .C ({1'b0 , uc_2090, uc_2091, uc_2092, uc_2093, uc_2094, 
    uc_2095, uc_2096, uc_2097, uc_2098, uc_2099, uc_2100, uc_2101, \intermediateWiresStage1[14][50] , 
    \intermediateWiresStage1[14][49] , \intermediateWiresStage1[14][48] , \intermediateWiresStage1[14][47] , 
    \intermediateWiresStage1[14][46] , \intermediateWiresStage1[14][45] , \intermediateWiresStage1[14][44] , 
    \intermediateWiresStage1[14][43] , \intermediateWiresStage1[14][42] , \intermediateWiresStage1[14][41] , 
    \intermediateWiresStage1[14][40] , \intermediateWiresStage1[14][39] , \intermediateWiresStage1[14][38] , 
    \intermediateWiresStage1[14][37] , \intermediateWiresStage1[14][36] , \intermediateWiresStage1[14][35] , 
    \intermediateWiresStage1[14][34] , \intermediateWiresStage1[14][33] , \intermediateWiresStage1[14][32] , 
    \intermediateWiresStage1[14][31] , \intermediateWiresStage1[14][30] , \intermediateWiresStage1[14][29] , 
    \intermediateWiresStage1[14][28] , \intermediateWiresStage1[14][27] , \intermediateWiresStage1[14][26] , 
    \intermediateWiresStage1[14][25] , \intermediateWiresStage1[14][24] , \intermediateWiresStage1[14][23] , 
    \intermediateWiresStage1[14][22] , normalizedWires[1365], uc_2102, uc_2103, uc_2104, 
    uc_2105, uc_2106, uc_2107, uc_2108, uc_2109, uc_2110, uc_2111, uc_2112, uc_2113, 
    uc_2114, uc_2115, uc_2116, uc_2117, uc_2118, uc_2119, uc_2120, uc_2121, uc_2122}));
CSAlike__2_753 genblk3_5_parallelAdderStage2 (.carry ({uc_1834, uc_1835, uc_1836, 
    uc_1837, uc_1838, uc_1839, \intermediateWiresStage2[11][57] , \intermediateWiresStage2[11][56] , 
    \intermediateWiresStage2[11][55] , \intermediateWiresStage2[11][54] , \intermediateWiresStage2[11][53] , 
    \intermediateWiresStage2[11][52] , \intermediateWiresStage2[11][51] , \intermediateWiresStage2[11][50] , 
    \intermediateWiresStage2[11][49] , \intermediateWiresStage2[11][48] , \intermediateWiresStage2[11][47] , 
    \intermediateWiresStage2[11][46] , \intermediateWiresStage2[11][45] , \intermediateWiresStage2[11][44] , 
    \intermediateWiresStage2[11][43] , \intermediateWiresStage2[11][42] , \intermediateWiresStage2[11][41] , 
    \intermediateWiresStage2[11][40] , \intermediateWiresStage2[11][39] , \intermediateWiresStage2[11][38] , 
    \intermediateWiresStage2[11][37] , \intermediateWiresStage2[11][36] , \intermediateWiresStage2[11][35] , 
    \intermediateWiresStage2[11][34] , \intermediateWiresStage2[11][33] , \intermediateWiresStage2[11][32] , 
    \intermediateWiresStage2[11][31] , \intermediateWiresStage2[11][30] , \intermediateWiresStage2[11][29] , 
    \intermediateWiresStage2[11][28] , \intermediateWiresStage2[11][27] , \intermediateWiresStage2[11][26] , 
    \intermediateWiresStage2[11][25] , uc_1840, uc_1841, uc_1842, uc_1843, uc_1844, 
    uc_1845, uc_1846, uc_1847, uc_1848, uc_1849, uc_1850, uc_1851, uc_1852, uc_1853, 
    uc_1854, uc_1855, uc_1856, uc_1857, uc_1858, uc_1859, uc_1860, uc_1861, uc_1862, 
    uc_1863, uc_1864}), .result ({uc_1803, uc_1804, uc_1805, uc_1806, uc_1807, uc_1808, 
    uc_1809, \intermediateWiresStage2[10][56] , \intermediateWiresStage2[10][55] , 
    \intermediateWiresStage2[10][54] , \intermediateWiresStage2[10][53] , \intermediateWiresStage2[10][52] , 
    \intermediateWiresStage2[10][51] , \intermediateWiresStage2[10][50] , \intermediateWiresStage2[10][49] , 
    \intermediateWiresStage2[10][48] , \intermediateWiresStage2[10][47] , \intermediateWiresStage2[10][46] , 
    \intermediateWiresStage2[10][45] , \intermediateWiresStage2[10][44] , \intermediateWiresStage2[10][43] , 
    \intermediateWiresStage2[10][42] , \intermediateWiresStage2[10][41] , \intermediateWiresStage2[10][40] , 
    \intermediateWiresStage2[10][39] , \intermediateWiresStage2[10][38] , \intermediateWiresStage2[10][37] , 
    \intermediateWiresStage2[10][36] , \intermediateWiresStage2[10][35] , \intermediateWiresStage2[10][34] , 
    \intermediateWiresStage2[10][33] , \intermediateWiresStage2[10][32] , \intermediateWiresStage2[10][31] , 
    \intermediateWiresStage2[10][30] , \intermediateWiresStage2[10][29] , \intermediateWiresStage2[10][28] , 
    \intermediateWiresStage2[10][27] , \intermediateWiresStage2[10][26] , \intermediateWiresStage2[10][25] , 
    \intermediateWiresStage2[10][24] , uc_1810, uc_1811, uc_1812, uc_1813, uc_1814, 
    uc_1815, uc_1816, uc_1817, uc_1818, uc_1819, uc_1820, uc_1821, uc_1822, uc_1823, 
    uc_1824, uc_1825, uc_1826, uc_1827, uc_1828, uc_1829, uc_1830, uc_1831, uc_1832, 
    uc_1833}), .A ({1'b0 , uc_1865, uc_1866, uc_1867, uc_1868, uc_1869, uc_1870, 
    uc_1871, uc_1872, uc_1873, \intermediateWiresStage1[15][53] , \intermediateWiresStage1[15][52] , 
    \intermediateWiresStage1[15][51] , \intermediateWiresStage1[15][50] , \intermediateWiresStage1[15][49] , 
    \intermediateWiresStage1[15][48] , \intermediateWiresStage1[15][47] , \intermediateWiresStage1[15][46] , 
    \intermediateWiresStage1[15][45] , \intermediateWiresStage1[15][44] , \intermediateWiresStage1[15][43] , 
    \intermediateWiresStage1[15][42] , \intermediateWiresStage1[15][41] , \intermediateWiresStage1[15][40] , 
    \intermediateWiresStage1[15][39] , \intermediateWiresStage1[15][38] , \intermediateWiresStage1[15][37] , 
    \intermediateWiresStage1[15][36] , \intermediateWiresStage1[15][35] , \intermediateWiresStage1[15][34] , 
    \intermediateWiresStage1[15][33] , \intermediateWiresStage1[15][32] , \intermediateWiresStage1[15][31] , 
    \intermediateWiresStage1[15][30] , \intermediateWiresStage1[15][29] , \intermediateWiresStage1[15][28] , 
    \intermediateWiresStage1[15][27] , \intermediateWiresStage1[15][26] , \intermediateWiresStage1[15][25] , 
    \intermediateWiresStage1[15][24] , uc_1874, uc_1875, uc_1876, uc_1877, uc_1878, 
    uc_1879, uc_1880, uc_1881, uc_1882, uc_1883, uc_1884, uc_1885, uc_1886, uc_1887, 
    uc_1888, uc_1889, uc_1890, uc_1891, uc_1892, uc_1893, uc_1894, uc_1895, uc_1896, 
    uc_1897}), .B ({1'b0 , uc_1898, uc_1899, uc_1900, uc_1901, uc_1902, uc_1903, 
    normalizedWires[1720], \intermediateWiresStage1[16][55] , \intermediateWiresStage1[16][54] , 
    \intermediateWiresStage1[16][53] , \intermediateWiresStage1[16][52] , \intermediateWiresStage1[16][51] , 
    \intermediateWiresStage1[16][50] , \intermediateWiresStage1[16][49] , \intermediateWiresStage1[16][48] , 
    \intermediateWiresStage1[16][47] , \intermediateWiresStage1[16][46] , \intermediateWiresStage1[16][45] , 
    \intermediateWiresStage1[16][44] , \intermediateWiresStage1[16][43] , \intermediateWiresStage1[16][42] , 
    \intermediateWiresStage1[16][41] , \intermediateWiresStage1[16][40] , \intermediateWiresStage1[16][39] , 
    \intermediateWiresStage1[16][38] , \intermediateWiresStage1[16][37] , \intermediateWiresStage1[16][36] , 
    \intermediateWiresStage1[16][35] , \intermediateWiresStage1[16][34] , \intermediateWiresStage1[16][33] , 
    \intermediateWiresStage1[16][32] , \intermediateWiresStage1[16][31] , \intermediateWiresStage1[16][30] , 
    \intermediateWiresStage1[16][29] , \intermediateWiresStage1[16][28] , \intermediateWiresStage1[16][27] , 
    \intermediateWiresStage1[16][26] , \intermediateWiresStage1[16][25] , normalizedWires[1560], 
    uc_1904, uc_1905, uc_1906, uc_1907, uc_1908, uc_1909, uc_1910, uc_1911, uc_1912, 
    uc_1913, uc_1914, uc_1915, uc_1916, uc_1917, uc_1918, uc_1919, uc_1920, uc_1921, 
    uc_1922, uc_1923, uc_1924, uc_1925, uc_1926, uc_1927}), .C ({1'b0 , uc_1928, 
    uc_1929, uc_1930, uc_1931, uc_1932, uc_1933, \intermediateWiresStage1[17][56] , 
    \intermediateWiresStage1[17][55] , \intermediateWiresStage1[17][54] , \intermediateWiresStage1[17][53] , 
    \intermediateWiresStage1[17][52] , \intermediateWiresStage1[17][51] , \intermediateWiresStage1[17][50] , 
    \intermediateWiresStage1[17][49] , \intermediateWiresStage1[17][48] , \intermediateWiresStage1[17][47] , 
    \intermediateWiresStage1[17][46] , \intermediateWiresStage1[17][45] , \intermediateWiresStage1[17][44] , 
    \intermediateWiresStage1[17][43] , \intermediateWiresStage1[17][42] , \intermediateWiresStage1[17][41] , 
    \intermediateWiresStage1[17][40] , \intermediateWiresStage1[17][39] , \intermediateWiresStage1[17][38] , 
    \intermediateWiresStage1[17][37] , \intermediateWiresStage1[17][36] , \intermediateWiresStage1[17][35] , 
    \intermediateWiresStage1[17][34] , \intermediateWiresStage1[17][33] , \intermediateWiresStage1[17][32] , 
    \intermediateWiresStage1[17][31] , \intermediateWiresStage1[17][30] , \intermediateWiresStage1[17][29] , 
    \intermediateWiresStage1[17][28] , \intermediateWiresStage1[17][27] , \intermediateWiresStage1[17][26] , 
    uc_1934, uc_1935, uc_1936, uc_1937, uc_1938, uc_1939, uc_1940, uc_1941, uc_1942, 
    uc_1943, uc_1944, uc_1945, uc_1946, uc_1947, uc_1948, uc_1949, uc_1950, uc_1951, 
    uc_1952, uc_1953, uc_1954, uc_1955, uc_1956, uc_1957, uc_1958, uc_1959}));
CSAlike__2_500 genblk3_6_parallelAdderStage2 (.carry ({uc_1673, uc_1674, uc_1675, 
    \intermediateWiresStage2[13][60] , \intermediateWiresStage2[13][59] , \intermediateWiresStage2[13][58] , 
    \intermediateWiresStage2[13][57] , \intermediateWiresStage2[13][56] , \intermediateWiresStage2[13][55] , 
    \intermediateWiresStage2[13][54] , \intermediateWiresStage2[13][53] , \intermediateWiresStage2[13][52] , 
    \intermediateWiresStage2[13][51] , \intermediateWiresStage2[13][50] , \intermediateWiresStage2[13][49] , 
    \intermediateWiresStage2[13][48] , \intermediateWiresStage2[13][47] , \intermediateWiresStage2[13][46] , 
    \intermediateWiresStage2[13][45] , \intermediateWiresStage2[13][44] , \intermediateWiresStage2[13][43] , 
    \intermediateWiresStage2[13][42] , \intermediateWiresStage2[13][41] , \intermediateWiresStage2[13][40] , 
    \intermediateWiresStage2[13][39] , \intermediateWiresStage2[13][38] , \intermediateWiresStage2[13][37] , 
    \intermediateWiresStage2[13][36] , \intermediateWiresStage2[13][35] , \intermediateWiresStage2[13][34] , 
    \intermediateWiresStage2[13][33] , \intermediateWiresStage2[13][32] , \intermediateWiresStage2[13][31] , 
    \intermediateWiresStage2[13][30] , uc_1676, uc_1677, uc_1678, uc_1679, uc_1680, 
    uc_1681, uc_1682, uc_1683, uc_1684, uc_1685, uc_1686, uc_1687, uc_1688, uc_1689, 
    uc_1690, uc_1691, uc_1692, uc_1693, uc_1694, uc_1695, uc_1696, uc_1697, uc_1698, 
    uc_1699, uc_1700, uc_1701, uc_1702, uc_1703, uc_1704, uc_1705}), .result ({uc_1640, 
    uc_1641, uc_1642, uc_1643, \intermediateWiresStage2[12][59] , \intermediateWiresStage2[12][58] , 
    \intermediateWiresStage2[12][57] , \intermediateWiresStage2[12][56] , \intermediateWiresStage2[12][55] , 
    \intermediateWiresStage2[12][54] , \intermediateWiresStage2[12][53] , \intermediateWiresStage2[12][52] , 
    \intermediateWiresStage2[12][51] , \intermediateWiresStage2[12][50] , \intermediateWiresStage2[12][49] , 
    \intermediateWiresStage2[12][48] , \intermediateWiresStage2[12][47] , \intermediateWiresStage2[12][46] , 
    \intermediateWiresStage2[12][45] , \intermediateWiresStage2[12][44] , \intermediateWiresStage2[12][43] , 
    \intermediateWiresStage2[12][42] , \intermediateWiresStage2[12][41] , \intermediateWiresStage2[12][40] , 
    \intermediateWiresStage2[12][39] , \intermediateWiresStage2[12][38] , \intermediateWiresStage2[12][37] , 
    \intermediateWiresStage2[12][36] , \intermediateWiresStage2[12][35] , \intermediateWiresStage2[12][34] , 
    \intermediateWiresStage2[12][33] , \intermediateWiresStage2[12][32] , \intermediateWiresStage2[12][31] , 
    \intermediateWiresStage2[12][30] , \intermediateWiresStage2[12][29] , uc_1644, 
    uc_1645, uc_1646, uc_1647, uc_1648, uc_1649, uc_1650, uc_1651, uc_1652, uc_1653, 
    uc_1654, uc_1655, uc_1656, uc_1657, uc_1658, uc_1659, uc_1660, uc_1661, uc_1662, 
    uc_1663, uc_1664, uc_1665, uc_1666, uc_1667, uc_1668, uc_1669, uc_1670, uc_1671, 
    uc_1672}), .A ({1'b0 , uc_1706, uc_1707, uc_1708, normalizedWires[1915], \intermediateWiresStage1[18][58] , 
    \intermediateWiresStage1[18][57] , \intermediateWiresStage1[18][56] , \intermediateWiresStage1[18][55] , 
    \intermediateWiresStage1[18][54] , \intermediateWiresStage1[18][53] , \intermediateWiresStage1[18][52] , 
    \intermediateWiresStage1[18][51] , \intermediateWiresStage1[18][50] , \intermediateWiresStage1[18][49] , 
    \intermediateWiresStage1[18][48] , \intermediateWiresStage1[18][47] , \intermediateWiresStage1[18][46] , 
    \intermediateWiresStage1[18][45] , \intermediateWiresStage1[18][44] , \intermediateWiresStage1[18][43] , 
    \intermediateWiresStage1[18][42] , \intermediateWiresStage1[18][41] , \intermediateWiresStage1[18][40] , 
    \intermediateWiresStage1[18][39] , \intermediateWiresStage1[18][38] , \intermediateWiresStage1[18][37] , 
    \intermediateWiresStage1[18][36] , \intermediateWiresStage1[18][35] , \intermediateWiresStage1[18][34] , 
    \intermediateWiresStage1[18][33] , \intermediateWiresStage1[18][32] , \intermediateWiresStage1[18][31] , 
    \intermediateWiresStage1[18][30] , \intermediateWiresStage1[18][29] , uc_1709, 
    uc_1710, uc_1711, uc_1712, uc_1713, uc_1714, uc_1715, uc_1716, uc_1717, uc_1718, 
    uc_1719, uc_1720, uc_1721, uc_1722, uc_1723, uc_1724, uc_1725, uc_1726, uc_1727, 
    uc_1728, uc_1729, uc_1730, uc_1731, uc_1732, uc_1733, uc_1734, uc_1735, uc_1736, 
    uc_1737}), .B ({1'b0 , uc_1738, uc_1739, uc_1740, \intermediateWiresStage1[19][59] , 
    \intermediateWiresStage1[19][58] , \intermediateWiresStage1[19][57] , \intermediateWiresStage1[19][56] , 
    \intermediateWiresStage1[19][55] , \intermediateWiresStage1[19][54] , \intermediateWiresStage1[19][53] , 
    \intermediateWiresStage1[19][52] , \intermediateWiresStage1[19][51] , \intermediateWiresStage1[19][50] , 
    \intermediateWiresStage1[19][49] , \intermediateWiresStage1[19][48] , \intermediateWiresStage1[19][47] , 
    \intermediateWiresStage1[19][46] , \intermediateWiresStage1[19][45] , \intermediateWiresStage1[19][44] , 
    \intermediateWiresStage1[19][43] , \intermediateWiresStage1[19][42] , \intermediateWiresStage1[19][41] , 
    \intermediateWiresStage1[19][40] , \intermediateWiresStage1[19][39] , \intermediateWiresStage1[19][38] , 
    \intermediateWiresStage1[19][37] , \intermediateWiresStage1[19][36] , \intermediateWiresStage1[19][35] , 
    \intermediateWiresStage1[19][34] , \intermediateWiresStage1[19][33] , \intermediateWiresStage1[19][32] , 
    \intermediateWiresStage1[19][31] , \intermediateWiresStage1[19][30] , \intermediateWiresStage1[19][29] , 
    uc_1741, uc_1742, uc_1743, uc_1744, uc_1745, uc_1746, uc_1747, uc_1748, uc_1749, 
    uc_1750, uc_1751, uc_1752, uc_1753, uc_1754, uc_1755, uc_1756, uc_1757, uc_1758, 
    uc_1759, uc_1760, uc_1761, uc_1762, uc_1763, uc_1764, uc_1765, uc_1766, uc_1767, 
    uc_1768, uc_1769}), .C ({1'b0 , uc_1770, uc_1771, uc_1772, normalizedWires[1979], 
    normalizedWires[1978], normalizedWires[1977], normalizedWires[1976], normalizedWires[1975], 
    normalizedWires[1974], normalizedWires[1973], normalizedWires[1972], normalizedWires[1971], 
    normalizedWires[1970], normalizedWires[1969], normalizedWires[1968], normalizedWires[1967], 
    normalizedWires[1966], normalizedWires[1965], normalizedWires[1964], normalizedWires[1963], 
    normalizedWires[1962], normalizedWires[1961], normalizedWires[1960], normalizedWires[1959], 
    normalizedWires[1958], normalizedWires[1957], normalizedWires[1956], normalizedWires[1955], 
    normalizedWires[1954], normalizedWires[1953], normalizedWires[1952], normalizedWires[1951], 
    normalizedWires[1950], uc_1773, uc_1774, uc_1775, uc_1776, uc_1777, uc_1778, 
    uc_1779, uc_1780, uc_1781, uc_1782, uc_1783, uc_1784, uc_1785, uc_1786, uc_1787, 
    uc_1788, uc_1789, uc_1790, uc_1791, uc_1792, uc_1793, uc_1794, uc_1795, uc_1796, 
    uc_1797, uc_1798, uc_1799, uc_1800, uc_1801, uc_1802}));
CSAlike__0_108 genblk2_0_parallelAdderStage1 (.carry ({uc_1509, uc_1510, uc_1511, 
    uc_1512, uc_1513, uc_1514, uc_1515, uc_1516, uc_1517, uc_1518, uc_1519, uc_1520, 
    uc_1521, uc_1522, uc_1523, uc_1524, uc_1525, uc_1526, uc_1527, uc_1528, uc_1529, 
    uc_1530, uc_1531, uc_1532, uc_1533, uc_1534, uc_1535, uc_1536, uc_1537, uc_1538, 
    uc_1539, \intermediateWiresStage1[1][32] , \intermediateWiresStage1[1][31] , 
    \intermediateWiresStage1[1][30] , \intermediateWiresStage1[1][29] , \intermediateWiresStage1[1][28] , 
    \intermediateWiresStage1[1][27] , \intermediateWiresStage1[1][26] , \intermediateWiresStage1[1][25] , 
    \intermediateWiresStage1[1][24] , \intermediateWiresStage1[1][23] , \intermediateWiresStage1[1][22] , 
    \intermediateWiresStage1[1][21] , \intermediateWiresStage1[1][20] , \intermediateWiresStage1[1][19] , 
    \intermediateWiresStage1[1][18] , \intermediateWiresStage1[1][17] , \intermediateWiresStage1[1][16] , 
    \intermediateWiresStage1[1][15] , \intermediateWiresStage1[1][14] , \intermediateWiresStage1[1][13] , 
    \intermediateWiresStage1[1][12] , \intermediateWiresStage1[1][11] , \intermediateWiresStage1[1][10] , 
    \intermediateWiresStage1[1][9] , \intermediateWiresStage1[1][8] , \intermediateWiresStage1[1][7] , 
    \intermediateWiresStage1[1][6] , \intermediateWiresStage1[1][5] , \intermediateWiresStage1[1][4] , 
    \intermediateWiresStage1[1][3] , \intermediateWiresStage1[1][2] , uc_1540, uc_1541})
    , .result ({uc_1476, uc_1477, uc_1478, uc_1479, uc_1480, uc_1481, uc_1482, uc_1483, 
    uc_1484, uc_1485, uc_1486, uc_1487, uc_1488, uc_1489, uc_1490, uc_1491, uc_1492, 
    uc_1493, uc_1494, uc_1495, uc_1496, uc_1497, uc_1498, uc_1499, uc_1500, uc_1501, 
    uc_1502, uc_1503, uc_1504, uc_1505, uc_1506, uc_1507, \intermediateWiresStage1[0][31] , 
    \intermediateWiresStage1[0][30] , \intermediateWiresStage1[0][29] , \intermediateWiresStage1[0][28] , 
    \intermediateWiresStage1[0][27] , \intermediateWiresStage1[0][26] , \intermediateWiresStage1[0][25] , 
    \intermediateWiresStage1[0][24] , \intermediateWiresStage1[0][23] , \intermediateWiresStage1[0][22] , 
    \intermediateWiresStage1[0][21] , \intermediateWiresStage1[0][20] , \intermediateWiresStage1[0][19] , 
    \intermediateWiresStage1[0][18] , \intermediateWiresStage1[0][17] , \intermediateWiresStage1[0][16] , 
    \intermediateWiresStage1[0][15] , \intermediateWiresStage1[0][14] , \intermediateWiresStage1[0][13] , 
    \intermediateWiresStage1[0][12] , \intermediateWiresStage1[0][11] , \intermediateWiresStage1[0][10] , 
    \intermediateWiresStage1[0][9] , \intermediateWiresStage1[0][8] , \intermediateWiresStage1[0][7] , 
    \intermediateWiresStage1[0][6] , \intermediateWiresStage1[0][5] , \intermediateWiresStage1[0][4] , 
    \intermediateWiresStage1[0][3] , \intermediateWiresStage1[0][2] , Res[1], uc_1508})
    , .A ({1'b0 , uc_1542, uc_1543, uc_1544, uc_1545, uc_1546, uc_1547, uc_1548, 
    uc_1549, uc_1550, uc_1551, uc_1552, uc_1553, uc_1554, uc_1555, uc_1556, uc_1557, 
    uc_1558, uc_1559, uc_1560, uc_1561, uc_1562, uc_1563, uc_1564, uc_1565, uc_1566, 
    uc_1567, uc_1568, uc_1569, uc_1570, uc_1571, uc_1572, uc_1573, normalizedWires[30], 
    normalizedWires[29], normalizedWires[28], normalizedWires[27], normalizedWires[26], 
    normalizedWires[25], normalizedWires[24], normalizedWires[23], normalizedWires[22], 
    normalizedWires[21], normalizedWires[20], normalizedWires[19], normalizedWires[18], 
    normalizedWires[17], normalizedWires[16], normalizedWires[15], normalizedWires[14], 
    normalizedWires[13], normalizedWires[12], normalizedWires[11], normalizedWires[10], 
    normalizedWires[9], normalizedWires[8], normalizedWires[7], normalizedWires[6], 
    normalizedWires[5], normalizedWires[4], normalizedWires[3], normalizedWires[2], 
    normalizedWires[1], uc_1574}), .B ({1'b0 , uc_1575, uc_1576, uc_1577, uc_1578, 
    uc_1579, uc_1580, uc_1581, uc_1582, uc_1583, uc_1584, uc_1585, uc_1586, uc_1587, 
    uc_1588, uc_1589, uc_1590, uc_1591, uc_1592, uc_1593, uc_1594, uc_1595, uc_1596, 
    uc_1597, uc_1598, uc_1599, uc_1600, uc_1601, uc_1602, uc_1603, uc_1604, uc_1605, 
    normalizedWires[95], normalizedWires[94], normalizedWires[93], normalizedWires[92], 
    normalizedWires[91], normalizedWires[90], normalizedWires[89], normalizedWires[88], 
    normalizedWires[87], normalizedWires[86], normalizedWires[85], normalizedWires[84], 
    normalizedWires[83], normalizedWires[82], normalizedWires[81], normalizedWires[80], 
    normalizedWires[79], normalizedWires[78], normalizedWires[77], normalizedWires[76], 
    normalizedWires[75], normalizedWires[74], normalizedWires[73], normalizedWires[72], 
    normalizedWires[71], normalizedWires[70], normalizedWires[69], normalizedWires[68], 
    normalizedWires[67], normalizedWires[66], normalizedWires[65], uc_1606}), .C ({
    1'b0 , uc_1607, uc_1608, uc_1609, uc_1610, uc_1611, uc_1612, uc_1613, uc_1614, 
    uc_1615, uc_1616, uc_1617, uc_1618, uc_1619, uc_1620, uc_1621, uc_1622, uc_1623, 
    uc_1624, uc_1625, uc_1626, uc_1627, uc_1628, uc_1629, uc_1630, uc_1631, uc_1632, 
    uc_1633, uc_1634, uc_1635, uc_1636, uc_1637, normalizedWires[159], normalizedWires[158], 
    normalizedWires[157], normalizedWires[156], normalizedWires[155], normalizedWires[154], 
    normalizedWires[153], normalizedWires[152], normalizedWires[151], normalizedWires[150], 
    normalizedWires[149], normalizedWires[148], normalizedWires[147], normalizedWires[146], 
    normalizedWires[145], normalizedWires[144], normalizedWires[143], normalizedWires[142], 
    normalizedWires[141], normalizedWires[140], normalizedWires[139], normalizedWires[138], 
    normalizedWires[137], normalizedWires[136], normalizedWires[135], normalizedWires[134], 
    normalizedWires[133], normalizedWires[132], normalizedWires[131], normalizedWires[130], 
    uc_1638, uc_1639}));
CSAlike__1_2524 genblk2_1_parallelAdderStage1 (.carry ({uc_1345, uc_1346, uc_1347, 
    uc_1348, uc_1349, uc_1350, uc_1351, uc_1352, uc_1353, uc_1354, uc_1355, uc_1356, 
    uc_1357, uc_1358, uc_1359, uc_1360, uc_1361, uc_1362, uc_1363, uc_1364, uc_1365, 
    uc_1366, uc_1367, uc_1368, uc_1369, uc_1370, uc_1371, uc_1372, \intermediateWiresStage1[3][35] , 
    \intermediateWiresStage1[3][34] , \intermediateWiresStage1[3][33] , \intermediateWiresStage1[3][32] , 
    \intermediateWiresStage1[3][31] , \intermediateWiresStage1[3][30] , \intermediateWiresStage1[3][29] , 
    \intermediateWiresStage1[3][28] , \intermediateWiresStage1[3][27] , \intermediateWiresStage1[3][26] , 
    \intermediateWiresStage1[3][25] , \intermediateWiresStage1[3][24] , \intermediateWiresStage1[3][23] , 
    \intermediateWiresStage1[3][22] , \intermediateWiresStage1[3][21] , \intermediateWiresStage1[3][20] , 
    \intermediateWiresStage1[3][19] , \intermediateWiresStage1[3][18] , \intermediateWiresStage1[3][17] , 
    \intermediateWiresStage1[3][16] , \intermediateWiresStage1[3][15] , \intermediateWiresStage1[3][14] , 
    \intermediateWiresStage1[3][13] , \intermediateWiresStage1[3][12] , \intermediateWiresStage1[3][11] , 
    \intermediateWiresStage1[3][10] , \intermediateWiresStage1[3][9] , \intermediateWiresStage1[3][8] , 
    \intermediateWiresStage1[3][7] , \intermediateWiresStage1[3][6] , \intermediateWiresStage1[3][5] , 
    uc_1373, uc_1374, uc_1375, uc_1376, uc_1377}), .result ({uc_1312, uc_1313, uc_1314, 
    uc_1315, uc_1316, uc_1317, uc_1318, uc_1319, uc_1320, uc_1321, uc_1322, uc_1323, 
    uc_1324, uc_1325, uc_1326, uc_1327, uc_1328, uc_1329, uc_1330, uc_1331, uc_1332, 
    uc_1333, uc_1334, uc_1335, uc_1336, uc_1337, uc_1338, uc_1339, uc_1340, \intermediateWiresStage1[2][34] , 
    \intermediateWiresStage1[2][33] , \intermediateWiresStage1[2][32] , \intermediateWiresStage1[2][31] , 
    \intermediateWiresStage1[2][30] , \intermediateWiresStage1[2][29] , \intermediateWiresStage1[2][28] , 
    \intermediateWiresStage1[2][27] , \intermediateWiresStage1[2][26] , \intermediateWiresStage1[2][25] , 
    \intermediateWiresStage1[2][24] , \intermediateWiresStage1[2][23] , \intermediateWiresStage1[2][22] , 
    \intermediateWiresStage1[2][21] , \intermediateWiresStage1[2][20] , \intermediateWiresStage1[2][19] , 
    \intermediateWiresStage1[2][18] , \intermediateWiresStage1[2][17] , \intermediateWiresStage1[2][16] , 
    \intermediateWiresStage1[2][15] , \intermediateWiresStage1[2][14] , \intermediateWiresStage1[2][13] , 
    \intermediateWiresStage1[2][12] , \intermediateWiresStage1[2][11] , \intermediateWiresStage1[2][10] , 
    \intermediateWiresStage1[2][9] , \intermediateWiresStage1[2][8] , \intermediateWiresStage1[2][7] , 
    \intermediateWiresStage1[2][6] , \intermediateWiresStage1[2][5] , \intermediateWiresStage1[2][4] , 
    uc_1341, uc_1342, uc_1343, uc_1344}), .A ({1'b0 , uc_1378, uc_1379, uc_1380, 
    uc_1381, uc_1382, uc_1383, uc_1384, uc_1385, uc_1386, uc_1387, uc_1388, uc_1389, 
    uc_1390, uc_1391, uc_1392, uc_1393, uc_1394, uc_1395, uc_1396, uc_1397, uc_1398, 
    uc_1399, uc_1400, uc_1401, uc_1402, uc_1403, uc_1404, uc_1405, uc_1406, normalizedWires[225], 
    normalizedWires[224], normalizedWires[223], normalizedWires[222], normalizedWires[221], 
    normalizedWires[220], normalizedWires[219], normalizedWires[218], normalizedWires[217], 
    normalizedWires[216], normalizedWires[215], normalizedWires[214], normalizedWires[213], 
    normalizedWires[212], normalizedWires[211], normalizedWires[210], normalizedWires[209], 
    normalizedWires[208], normalizedWires[207], normalizedWires[206], normalizedWires[205], 
    normalizedWires[204], normalizedWires[203], normalizedWires[202], normalizedWires[201], 
    normalizedWires[200], normalizedWires[199], normalizedWires[198], normalizedWires[197], 
    normalizedWires[196], uc_1407, uc_1408, uc_1409, uc_1410}), .B ({1'b0 , uc_1411, 
    uc_1412, uc_1413, uc_1414, uc_1415, uc_1416, uc_1417, uc_1418, uc_1419, uc_1420, 
    uc_1421, uc_1422, uc_1423, uc_1424, uc_1425, uc_1426, uc_1427, uc_1428, uc_1429, 
    uc_1430, uc_1431, uc_1432, uc_1433, uc_1434, uc_1435, uc_1436, uc_1437, uc_1438, 
    normalizedWires[290], normalizedWires[289], normalizedWires[288], normalizedWires[287], 
    normalizedWires[286], normalizedWires[285], normalizedWires[284], normalizedWires[283], 
    normalizedWires[282], normalizedWires[281], normalizedWires[280], normalizedWires[279], 
    normalizedWires[278], normalizedWires[277], normalizedWires[276], normalizedWires[275], 
    normalizedWires[274], normalizedWires[273], normalizedWires[272], normalizedWires[271], 
    normalizedWires[270], normalizedWires[269], normalizedWires[268], normalizedWires[267], 
    normalizedWires[266], normalizedWires[265], normalizedWires[264], normalizedWires[263], 
    normalizedWires[262], normalizedWires[261], normalizedWires[260], uc_1439, uc_1440, 
    uc_1441, uc_1442}), .C ({1'b0 , uc_1443, uc_1444, uc_1445, uc_1446, uc_1447, 
    uc_1448, uc_1449, uc_1450, uc_1451, uc_1452, uc_1453, uc_1454, uc_1455, uc_1456, 
    uc_1457, uc_1458, uc_1459, uc_1460, uc_1461, uc_1462, uc_1463, uc_1464, uc_1465, 
    uc_1466, uc_1467, uc_1468, uc_1469, uc_1470, normalizedWires[354], normalizedWires[353], 
    normalizedWires[352], normalizedWires[351], normalizedWires[350], normalizedWires[349], 
    normalizedWires[348], normalizedWires[347], normalizedWires[346], normalizedWires[345], 
    normalizedWires[344], normalizedWires[343], normalizedWires[342], normalizedWires[341], 
    normalizedWires[340], normalizedWires[339], normalizedWires[338], normalizedWires[337], 
    normalizedWires[336], normalizedWires[335], normalizedWires[334], normalizedWires[333], 
    normalizedWires[332], normalizedWires[331], normalizedWires[330], normalizedWires[329], 
    normalizedWires[328], normalizedWires[327], normalizedWires[326], normalizedWires[325], 
    uc_1471, uc_1472, uc_1473, uc_1474, uc_1475}));
CSAlike__1_2271 genblk2_2_parallelAdderStage1 (.carry ({uc_1181, uc_1182, uc_1183, 
    uc_1184, uc_1185, uc_1186, uc_1187, uc_1188, uc_1189, uc_1190, uc_1191, uc_1192, 
    uc_1193, uc_1194, uc_1195, uc_1196, uc_1197, uc_1198, uc_1199, uc_1200, uc_1201, 
    uc_1202, uc_1203, uc_1204, uc_1205, \intermediateWiresStage1[5][38] , \intermediateWiresStage1[5][37] , 
    \intermediateWiresStage1[5][36] , \intermediateWiresStage1[5][35] , \intermediateWiresStage1[5][34] , 
    \intermediateWiresStage1[5][33] , \intermediateWiresStage1[5][32] , \intermediateWiresStage1[5][31] , 
    \intermediateWiresStage1[5][30] , \intermediateWiresStage1[5][29] , \intermediateWiresStage1[5][28] , 
    \intermediateWiresStage1[5][27] , \intermediateWiresStage1[5][26] , \intermediateWiresStage1[5][25] , 
    \intermediateWiresStage1[5][24] , \intermediateWiresStage1[5][23] , \intermediateWiresStage1[5][22] , 
    \intermediateWiresStage1[5][21] , \intermediateWiresStage1[5][20] , \intermediateWiresStage1[5][19] , 
    \intermediateWiresStage1[5][18] , \intermediateWiresStage1[5][17] , \intermediateWiresStage1[5][16] , 
    \intermediateWiresStage1[5][15] , \intermediateWiresStage1[5][14] , \intermediateWiresStage1[5][13] , 
    \intermediateWiresStage1[5][12] , \intermediateWiresStage1[5][11] , \intermediateWiresStage1[5][10] , 
    \intermediateWiresStage1[5][9] , \intermediateWiresStage1[5][8] , uc_1206, uc_1207, 
    uc_1208, uc_1209, uc_1210, uc_1211, uc_1212, uc_1213}), .result ({uc_1148, uc_1149, 
    uc_1150, uc_1151, uc_1152, uc_1153, uc_1154, uc_1155, uc_1156, uc_1157, uc_1158, 
    uc_1159, uc_1160, uc_1161, uc_1162, uc_1163, uc_1164, uc_1165, uc_1166, uc_1167, 
    uc_1168, uc_1169, uc_1170, uc_1171, uc_1172, uc_1173, \intermediateWiresStage1[4][37] , 
    \intermediateWiresStage1[4][36] , \intermediateWiresStage1[4][35] , \intermediateWiresStage1[4][34] , 
    \intermediateWiresStage1[4][33] , \intermediateWiresStage1[4][32] , \intermediateWiresStage1[4][31] , 
    \intermediateWiresStage1[4][30] , \intermediateWiresStage1[4][29] , \intermediateWiresStage1[4][28] , 
    \intermediateWiresStage1[4][27] , \intermediateWiresStage1[4][26] , \intermediateWiresStage1[4][25] , 
    \intermediateWiresStage1[4][24] , \intermediateWiresStage1[4][23] , \intermediateWiresStage1[4][22] , 
    \intermediateWiresStage1[4][21] , \intermediateWiresStage1[4][20] , \intermediateWiresStage1[4][19] , 
    \intermediateWiresStage1[4][18] , \intermediateWiresStage1[4][17] , \intermediateWiresStage1[4][16] , 
    \intermediateWiresStage1[4][15] , \intermediateWiresStage1[4][14] , \intermediateWiresStage1[4][13] , 
    \intermediateWiresStage1[4][12] , \intermediateWiresStage1[4][11] , \intermediateWiresStage1[4][10] , 
    \intermediateWiresStage1[4][9] , \intermediateWiresStage1[4][8] , \intermediateWiresStage1[4][7] , 
    uc_1174, uc_1175, uc_1176, uc_1177, uc_1178, uc_1179, uc_1180}), .A ({1'b0 , 
    uc_1214, uc_1215, uc_1216, uc_1217, uc_1218, uc_1219, uc_1220, uc_1221, uc_1222, 
    uc_1223, uc_1224, uc_1225, uc_1226, uc_1227, uc_1228, uc_1229, uc_1230, uc_1231, 
    uc_1232, uc_1233, uc_1234, uc_1235, uc_1236, uc_1237, uc_1238, uc_1239, normalizedWires[420], 
    normalizedWires[419], normalizedWires[418], normalizedWires[417], normalizedWires[416], 
    normalizedWires[415], normalizedWires[414], normalizedWires[413], normalizedWires[412], 
    normalizedWires[411], normalizedWires[410], normalizedWires[409], normalizedWires[408], 
    normalizedWires[407], normalizedWires[406], normalizedWires[405], normalizedWires[404], 
    normalizedWires[403], normalizedWires[402], normalizedWires[401], normalizedWires[400], 
    normalizedWires[399], normalizedWires[398], normalizedWires[397], normalizedWires[396], 
    normalizedWires[395], normalizedWires[394], normalizedWires[393], normalizedWires[392], 
    normalizedWires[391], uc_1240, uc_1241, uc_1242, uc_1243, uc_1244, uc_1245, uc_1246})
    , .B ({1'b0 , uc_1247, uc_1248, uc_1249, uc_1250, uc_1251, uc_1252, uc_1253, 
    uc_1254, uc_1255, uc_1256, uc_1257, uc_1258, uc_1259, uc_1260, uc_1261, uc_1262, 
    uc_1263, uc_1264, uc_1265, uc_1266, uc_1267, uc_1268, uc_1269, uc_1270, uc_1271, 
    normalizedWires[485], normalizedWires[484], normalizedWires[483], normalizedWires[482], 
    normalizedWires[481], normalizedWires[480], normalizedWires[479], normalizedWires[478], 
    normalizedWires[477], normalizedWires[476], normalizedWires[475], normalizedWires[474], 
    normalizedWires[473], normalizedWires[472], normalizedWires[471], normalizedWires[470], 
    normalizedWires[469], normalizedWires[468], normalizedWires[467], normalizedWires[466], 
    normalizedWires[465], normalizedWires[464], normalizedWires[463], normalizedWires[462], 
    normalizedWires[461], normalizedWires[460], normalizedWires[459], normalizedWires[458], 
    normalizedWires[457], normalizedWires[456], normalizedWires[455], uc_1272, uc_1273, 
    uc_1274, uc_1275, uc_1276, uc_1277, uc_1278}), .C ({1'b0 , uc_1279, uc_1280, 
    uc_1281, uc_1282, uc_1283, uc_1284, uc_1285, uc_1286, uc_1287, uc_1288, uc_1289, 
    uc_1290, uc_1291, uc_1292, uc_1293, uc_1294, uc_1295, uc_1296, uc_1297, uc_1298, 
    uc_1299, uc_1300, uc_1301, uc_1302, uc_1303, normalizedWires[549], normalizedWires[548], 
    normalizedWires[547], normalizedWires[546], normalizedWires[545], normalizedWires[544], 
    normalizedWires[543], normalizedWires[542], normalizedWires[541], normalizedWires[540], 
    normalizedWires[539], normalizedWires[538], normalizedWires[537], normalizedWires[536], 
    normalizedWires[535], normalizedWires[534], normalizedWires[533], normalizedWires[532], 
    normalizedWires[531], normalizedWires[530], normalizedWires[529], normalizedWires[528], 
    normalizedWires[527], normalizedWires[526], normalizedWires[525], normalizedWires[524], 
    normalizedWires[523], normalizedWires[522], normalizedWires[521], normalizedWires[520], 
    uc_1304, uc_1305, uc_1306, uc_1307, uc_1308, uc_1309, uc_1310, uc_1311}));
CSAlike__1_2018 genblk2_3_parallelAdderStage1 (.carry ({uc_1017, uc_1018, uc_1019, 
    uc_1020, uc_1021, uc_1022, uc_1023, uc_1024, uc_1025, uc_1026, uc_1027, uc_1028, 
    uc_1029, uc_1030, uc_1031, uc_1032, uc_1033, uc_1034, uc_1035, uc_1036, uc_1037, 
    uc_1038, \intermediateWiresStage1[7][41] , \intermediateWiresStage1[7][40] , 
    \intermediateWiresStage1[7][39] , \intermediateWiresStage1[7][38] , \intermediateWiresStage1[7][37] , 
    \intermediateWiresStage1[7][36] , \intermediateWiresStage1[7][35] , \intermediateWiresStage1[7][34] , 
    \intermediateWiresStage1[7][33] , \intermediateWiresStage1[7][32] , \intermediateWiresStage1[7][31] , 
    \intermediateWiresStage1[7][30] , \intermediateWiresStage1[7][29] , \intermediateWiresStage1[7][28] , 
    \intermediateWiresStage1[7][27] , \intermediateWiresStage1[7][26] , \intermediateWiresStage1[7][25] , 
    \intermediateWiresStage1[7][24] , \intermediateWiresStage1[7][23] , \intermediateWiresStage1[7][22] , 
    \intermediateWiresStage1[7][21] , \intermediateWiresStage1[7][20] , \intermediateWiresStage1[7][19] , 
    \intermediateWiresStage1[7][18] , \intermediateWiresStage1[7][17] , \intermediateWiresStage1[7][16] , 
    \intermediateWiresStage1[7][15] , \intermediateWiresStage1[7][14] , \intermediateWiresStage1[7][13] , 
    \intermediateWiresStage1[7][12] , \intermediateWiresStage1[7][11] , uc_1039, 
    uc_1040, uc_1041, uc_1042, uc_1043, uc_1044, uc_1045, uc_1046, uc_1047, uc_1048, 
    uc_1049}), .result ({uc_984, uc_985, uc_986, uc_987, uc_988, uc_989, uc_990, 
    uc_991, uc_992, uc_993, uc_994, uc_995, uc_996, uc_997, uc_998, uc_999, uc_1000, 
    uc_1001, uc_1002, uc_1003, uc_1004, uc_1005, uc_1006, \intermediateWiresStage1[6][40] , 
    \intermediateWiresStage1[6][39] , \intermediateWiresStage1[6][38] , \intermediateWiresStage1[6][37] , 
    \intermediateWiresStage1[6][36] , \intermediateWiresStage1[6][35] , \intermediateWiresStage1[6][34] , 
    \intermediateWiresStage1[6][33] , \intermediateWiresStage1[6][32] , \intermediateWiresStage1[6][31] , 
    \intermediateWiresStage1[6][30] , \intermediateWiresStage1[6][29] , \intermediateWiresStage1[6][28] , 
    \intermediateWiresStage1[6][27] , \intermediateWiresStage1[6][26] , \intermediateWiresStage1[6][25] , 
    \intermediateWiresStage1[6][24] , \intermediateWiresStage1[6][23] , \intermediateWiresStage1[6][22] , 
    \intermediateWiresStage1[6][21] , \intermediateWiresStage1[6][20] , \intermediateWiresStage1[6][19] , 
    \intermediateWiresStage1[6][18] , \intermediateWiresStage1[6][17] , \intermediateWiresStage1[6][16] , 
    \intermediateWiresStage1[6][15] , \intermediateWiresStage1[6][14] , \intermediateWiresStage1[6][13] , 
    \intermediateWiresStage1[6][12] , \intermediateWiresStage1[6][11] , \intermediateWiresStage1[6][10] , 
    uc_1007, uc_1008, uc_1009, uc_1010, uc_1011, uc_1012, uc_1013, uc_1014, uc_1015, 
    uc_1016}), .A ({1'b0 , uc_1050, uc_1051, uc_1052, uc_1053, uc_1054, uc_1055, 
    uc_1056, uc_1057, uc_1058, uc_1059, uc_1060, uc_1061, uc_1062, uc_1063, uc_1064, 
    uc_1065, uc_1066, uc_1067, uc_1068, uc_1069, uc_1070, uc_1071, uc_1072, normalizedWires[615], 
    normalizedWires[614], normalizedWires[613], normalizedWires[612], normalizedWires[611], 
    normalizedWires[610], normalizedWires[609], normalizedWires[608], normalizedWires[607], 
    normalizedWires[606], normalizedWires[605], normalizedWires[604], normalizedWires[603], 
    normalizedWires[602], normalizedWires[601], normalizedWires[600], normalizedWires[599], 
    normalizedWires[598], normalizedWires[597], normalizedWires[596], normalizedWires[595], 
    normalizedWires[594], normalizedWires[593], normalizedWires[592], normalizedWires[591], 
    normalizedWires[590], normalizedWires[589], normalizedWires[588], normalizedWires[587], 
    normalizedWires[586], uc_1073, uc_1074, uc_1075, uc_1076, uc_1077, uc_1078, uc_1079, 
    uc_1080, uc_1081, uc_1082}), .B ({1'b0 , uc_1083, uc_1084, uc_1085, uc_1086, 
    uc_1087, uc_1088, uc_1089, uc_1090, uc_1091, uc_1092, uc_1093, uc_1094, uc_1095, 
    uc_1096, uc_1097, uc_1098, uc_1099, uc_1100, uc_1101, uc_1102, uc_1103, uc_1104, 
    normalizedWires[680], normalizedWires[679], normalizedWires[678], normalizedWires[677], 
    normalizedWires[676], normalizedWires[675], normalizedWires[674], normalizedWires[673], 
    normalizedWires[672], normalizedWires[671], normalizedWires[670], normalizedWires[669], 
    normalizedWires[668], normalizedWires[667], normalizedWires[666], normalizedWires[665], 
    normalizedWires[664], normalizedWires[663], normalizedWires[662], normalizedWires[661], 
    normalizedWires[660], normalizedWires[659], normalizedWires[658], normalizedWires[657], 
    normalizedWires[656], normalizedWires[655], normalizedWires[654], normalizedWires[653], 
    normalizedWires[652], normalizedWires[651], normalizedWires[650], uc_1105, uc_1106, 
    uc_1107, uc_1108, uc_1109, uc_1110, uc_1111, uc_1112, uc_1113, uc_1114}), .C ({
    1'b0 , uc_1115, uc_1116, uc_1117, uc_1118, uc_1119, uc_1120, uc_1121, uc_1122, 
    uc_1123, uc_1124, uc_1125, uc_1126, uc_1127, uc_1128, uc_1129, uc_1130, uc_1131, 
    uc_1132, uc_1133, uc_1134, uc_1135, uc_1136, normalizedWires[744], normalizedWires[743], 
    normalizedWires[742], normalizedWires[741], normalizedWires[740], normalizedWires[739], 
    normalizedWires[738], normalizedWires[737], normalizedWires[736], normalizedWires[735], 
    normalizedWires[734], normalizedWires[733], normalizedWires[732], normalizedWires[731], 
    normalizedWires[730], normalizedWires[729], normalizedWires[728], normalizedWires[727], 
    normalizedWires[726], normalizedWires[725], normalizedWires[724], normalizedWires[723], 
    normalizedWires[722], normalizedWires[721], normalizedWires[720], normalizedWires[719], 
    normalizedWires[718], normalizedWires[717], normalizedWires[716], normalizedWires[715], 
    uc_1137, uc_1138, uc_1139, uc_1140, uc_1141, uc_1142, uc_1143, uc_1144, uc_1145, 
    uc_1146, uc_1147}));
CSAlike__1_1765 genblk2_4_parallelAdderStage1 (.carry ({uc_853, uc_854, uc_855, uc_856, 
    uc_857, uc_858, uc_859, uc_860, uc_861, uc_862, uc_863, uc_864, uc_865, uc_866, 
    uc_867, uc_868, uc_869, uc_870, uc_871, \intermediateWiresStage1[9][44] , \intermediateWiresStage1[9][43] , 
    \intermediateWiresStage1[9][42] , \intermediateWiresStage1[9][41] , \intermediateWiresStage1[9][40] , 
    \intermediateWiresStage1[9][39] , \intermediateWiresStage1[9][38] , \intermediateWiresStage1[9][37] , 
    \intermediateWiresStage1[9][36] , \intermediateWiresStage1[9][35] , \intermediateWiresStage1[9][34] , 
    \intermediateWiresStage1[9][33] , \intermediateWiresStage1[9][32] , \intermediateWiresStage1[9][31] , 
    \intermediateWiresStage1[9][30] , \intermediateWiresStage1[9][29] , \intermediateWiresStage1[9][28] , 
    \intermediateWiresStage1[9][27] , \intermediateWiresStage1[9][26] , \intermediateWiresStage1[9][25] , 
    \intermediateWiresStage1[9][24] , \intermediateWiresStage1[9][23] , \intermediateWiresStage1[9][22] , 
    \intermediateWiresStage1[9][21] , \intermediateWiresStage1[9][20] , \intermediateWiresStage1[9][19] , 
    \intermediateWiresStage1[9][18] , \intermediateWiresStage1[9][17] , \intermediateWiresStage1[9][16] , 
    \intermediateWiresStage1[9][15] , \intermediateWiresStage1[9][14] , uc_872, uc_873, 
    uc_874, uc_875, uc_876, uc_877, uc_878, uc_879, uc_880, uc_881, uc_882, uc_883, 
    uc_884, uc_885}), .result ({uc_820, uc_821, uc_822, uc_823, uc_824, uc_825, uc_826, 
    uc_827, uc_828, uc_829, uc_830, uc_831, uc_832, uc_833, uc_834, uc_835, uc_836, 
    uc_837, uc_838, uc_839, \intermediateWiresStage1[8][43] , \intermediateWiresStage1[8][42] , 
    \intermediateWiresStage1[8][41] , \intermediateWiresStage1[8][40] , \intermediateWiresStage1[8][39] , 
    \intermediateWiresStage1[8][38] , \intermediateWiresStage1[8][37] , \intermediateWiresStage1[8][36] , 
    \intermediateWiresStage1[8][35] , \intermediateWiresStage1[8][34] , \intermediateWiresStage1[8][33] , 
    \intermediateWiresStage1[8][32] , \intermediateWiresStage1[8][31] , \intermediateWiresStage1[8][30] , 
    \intermediateWiresStage1[8][29] , \intermediateWiresStage1[8][28] , \intermediateWiresStage1[8][27] , 
    \intermediateWiresStage1[8][26] , \intermediateWiresStage1[8][25] , \intermediateWiresStage1[8][24] , 
    \intermediateWiresStage1[8][23] , \intermediateWiresStage1[8][22] , \intermediateWiresStage1[8][21] , 
    \intermediateWiresStage1[8][20] , \intermediateWiresStage1[8][19] , \intermediateWiresStage1[8][18] , 
    \intermediateWiresStage1[8][17] , \intermediateWiresStage1[8][16] , \intermediateWiresStage1[8][15] , 
    \intermediateWiresStage1[8][14] , \intermediateWiresStage1[8][13] , uc_840, uc_841, 
    uc_842, uc_843, uc_844, uc_845, uc_846, uc_847, uc_848, uc_849, uc_850, uc_851, 
    uc_852}), .A ({1'b0 , uc_886, uc_887, uc_888, uc_889, uc_890, uc_891, uc_892, 
    uc_893, uc_894, uc_895, uc_896, uc_897, uc_898, uc_899, uc_900, uc_901, uc_902, 
    uc_903, uc_904, uc_905, normalizedWires[810], normalizedWires[809], normalizedWires[808], 
    normalizedWires[807], normalizedWires[806], normalizedWires[805], normalizedWires[804], 
    normalizedWires[803], normalizedWires[802], normalizedWires[801], normalizedWires[800], 
    normalizedWires[799], normalizedWires[798], normalizedWires[797], normalizedWires[796], 
    normalizedWires[795], normalizedWires[794], normalizedWires[793], normalizedWires[792], 
    normalizedWires[791], normalizedWires[790], normalizedWires[789], normalizedWires[788], 
    normalizedWires[787], normalizedWires[786], normalizedWires[785], normalizedWires[784], 
    normalizedWires[783], normalizedWires[782], normalizedWires[781], uc_906, uc_907, 
    uc_908, uc_909, uc_910, uc_911, uc_912, uc_913, uc_914, uc_915, uc_916, uc_917, 
    uc_918}), .B ({1'b0 , uc_919, uc_920, uc_921, uc_922, uc_923, uc_924, uc_925, 
    uc_926, uc_927, uc_928, uc_929, uc_930, uc_931, uc_932, uc_933, uc_934, uc_935, 
    uc_936, uc_937, normalizedWires[875], normalizedWires[874], normalizedWires[873], 
    normalizedWires[872], normalizedWires[871], normalizedWires[870], normalizedWires[869], 
    normalizedWires[868], normalizedWires[867], normalizedWires[866], normalizedWires[865], 
    normalizedWires[864], normalizedWires[863], normalizedWires[862], normalizedWires[861], 
    normalizedWires[860], normalizedWires[859], normalizedWires[858], normalizedWires[857], 
    normalizedWires[856], normalizedWires[855], normalizedWires[854], normalizedWires[853], 
    normalizedWires[852], normalizedWires[851], normalizedWires[850], normalizedWires[849], 
    normalizedWires[848], normalizedWires[847], normalizedWires[846], normalizedWires[845], 
    uc_938, uc_939, uc_940, uc_941, uc_942, uc_943, uc_944, uc_945, uc_946, uc_947, 
    uc_948, uc_949, uc_950}), .C ({1'b0 , uc_951, uc_952, uc_953, uc_954, uc_955, 
    uc_956, uc_957, uc_958, uc_959, uc_960, uc_961, uc_962, uc_963, uc_964, uc_965, 
    uc_966, uc_967, uc_968, uc_969, normalizedWires[939], normalizedWires[938], normalizedWires[937], 
    normalizedWires[936], normalizedWires[935], normalizedWires[934], normalizedWires[933], 
    normalizedWires[932], normalizedWires[931], normalizedWires[930], normalizedWires[929], 
    normalizedWires[928], normalizedWires[927], normalizedWires[926], normalizedWires[925], 
    normalizedWires[924], normalizedWires[923], normalizedWires[922], normalizedWires[921], 
    normalizedWires[920], normalizedWires[919], normalizedWires[918], normalizedWires[917], 
    normalizedWires[916], normalizedWires[915], normalizedWires[914], normalizedWires[913], 
    normalizedWires[912], normalizedWires[911], normalizedWires[910], uc_970, uc_971, 
    uc_972, uc_973, uc_974, uc_975, uc_976, uc_977, uc_978, uc_979, uc_980, uc_981, 
    uc_982, uc_983}));
CSAlike__1_1512 genblk2_5_parallelAdderStage1 (.carry ({uc_689, uc_690, uc_691, uc_692, 
    uc_693, uc_694, uc_695, uc_696, uc_697, uc_698, uc_699, uc_700, uc_701, uc_702, 
    uc_703, uc_704, \intermediateWiresStage1[11][47] , \intermediateWiresStage1[11][46] , 
    \intermediateWiresStage1[11][45] , \intermediateWiresStage1[11][44] , \intermediateWiresStage1[11][43] , 
    \intermediateWiresStage1[11][42] , \intermediateWiresStage1[11][41] , \intermediateWiresStage1[11][40] , 
    \intermediateWiresStage1[11][39] , \intermediateWiresStage1[11][38] , \intermediateWiresStage1[11][37] , 
    \intermediateWiresStage1[11][36] , \intermediateWiresStage1[11][35] , \intermediateWiresStage1[11][34] , 
    \intermediateWiresStage1[11][33] , \intermediateWiresStage1[11][32] , \intermediateWiresStage1[11][31] , 
    \intermediateWiresStage1[11][30] , \intermediateWiresStage1[11][29] , \intermediateWiresStage1[11][28] , 
    \intermediateWiresStage1[11][27] , \intermediateWiresStage1[11][26] , \intermediateWiresStage1[11][25] , 
    \intermediateWiresStage1[11][24] , \intermediateWiresStage1[11][23] , \intermediateWiresStage1[11][22] , 
    \intermediateWiresStage1[11][21] , \intermediateWiresStage1[11][20] , \intermediateWiresStage1[11][19] , 
    \intermediateWiresStage1[11][18] , \intermediateWiresStage1[11][17] , uc_705, 
    uc_706, uc_707, uc_708, uc_709, uc_710, uc_711, uc_712, uc_713, uc_714, uc_715, 
    uc_716, uc_717, uc_718, uc_719, uc_720, uc_721}), .result ({uc_656, uc_657, uc_658, 
    uc_659, uc_660, uc_661, uc_662, uc_663, uc_664, uc_665, uc_666, uc_667, uc_668, 
    uc_669, uc_670, uc_671, uc_672, \intermediateWiresStage1[10][46] , \intermediateWiresStage1[10][45] , 
    \intermediateWiresStage1[10][44] , \intermediateWiresStage1[10][43] , \intermediateWiresStage1[10][42] , 
    \intermediateWiresStage1[10][41] , \intermediateWiresStage1[10][40] , \intermediateWiresStage1[10][39] , 
    \intermediateWiresStage1[10][38] , \intermediateWiresStage1[10][37] , \intermediateWiresStage1[10][36] , 
    \intermediateWiresStage1[10][35] , \intermediateWiresStage1[10][34] , \intermediateWiresStage1[10][33] , 
    \intermediateWiresStage1[10][32] , \intermediateWiresStage1[10][31] , \intermediateWiresStage1[10][30] , 
    \intermediateWiresStage1[10][29] , \intermediateWiresStage1[10][28] , \intermediateWiresStage1[10][27] , 
    \intermediateWiresStage1[10][26] , \intermediateWiresStage1[10][25] , \intermediateWiresStage1[10][24] , 
    \intermediateWiresStage1[10][23] , \intermediateWiresStage1[10][22] , \intermediateWiresStage1[10][21] , 
    \intermediateWiresStage1[10][20] , \intermediateWiresStage1[10][19] , \intermediateWiresStage1[10][18] , 
    \intermediateWiresStage1[10][17] , \intermediateWiresStage1[10][16] , uc_673, 
    uc_674, uc_675, uc_676, uc_677, uc_678, uc_679, uc_680, uc_681, uc_682, uc_683, 
    uc_684, uc_685, uc_686, uc_687, uc_688}), .A ({1'b0 , uc_722, uc_723, uc_724, 
    uc_725, uc_726, uc_727, uc_728, uc_729, uc_730, uc_731, uc_732, uc_733, uc_734, 
    uc_735, uc_736, uc_737, uc_738, normalizedWires[1005], normalizedWires[1004], 
    normalizedWires[1003], normalizedWires[1002], normalizedWires[1001], normalizedWires[1000], 
    normalizedWires[999], normalizedWires[998], normalizedWires[997], normalizedWires[996], 
    normalizedWires[995], normalizedWires[994], normalizedWires[993], normalizedWires[992], 
    normalizedWires[991], normalizedWires[990], normalizedWires[989], normalizedWires[988], 
    normalizedWires[987], normalizedWires[986], normalizedWires[985], normalizedWires[984], 
    normalizedWires[983], normalizedWires[982], normalizedWires[981], normalizedWires[980], 
    normalizedWires[979], normalizedWires[978], normalizedWires[977], normalizedWires[976], 
    uc_739, uc_740, uc_741, uc_742, uc_743, uc_744, uc_745, uc_746, uc_747, uc_748, 
    uc_749, uc_750, uc_751, uc_752, uc_753, uc_754}), .B ({1'b0 , uc_755, uc_756, 
    uc_757, uc_758, uc_759, uc_760, uc_761, uc_762, uc_763, uc_764, uc_765, uc_766, 
    uc_767, uc_768, uc_769, uc_770, normalizedWires[1070], normalizedWires[1069], 
    normalizedWires[1068], normalizedWires[1067], normalizedWires[1066], normalizedWires[1065], 
    normalizedWires[1064], normalizedWires[1063], normalizedWires[1062], normalizedWires[1061], 
    normalizedWires[1060], normalizedWires[1059], normalizedWires[1058], normalizedWires[1057], 
    normalizedWires[1056], normalizedWires[1055], normalizedWires[1054], normalizedWires[1053], 
    normalizedWires[1052], normalizedWires[1051], normalizedWires[1050], normalizedWires[1049], 
    normalizedWires[1048], normalizedWires[1047], normalizedWires[1046], normalizedWires[1045], 
    normalizedWires[1044], normalizedWires[1043], normalizedWires[1042], normalizedWires[1041], 
    normalizedWires[1040], uc_771, uc_772, uc_773, uc_774, uc_775, uc_776, uc_777, 
    uc_778, uc_779, uc_780, uc_781, uc_782, uc_783, uc_784, uc_785, uc_786}), .C ({
    1'b0 , uc_787, uc_788, uc_789, uc_790, uc_791, uc_792, uc_793, uc_794, uc_795, 
    uc_796, uc_797, uc_798, uc_799, uc_800, uc_801, uc_802, normalizedWires[1134], 
    normalizedWires[1133], normalizedWires[1132], normalizedWires[1131], normalizedWires[1130], 
    normalizedWires[1129], normalizedWires[1128], normalizedWires[1127], normalizedWires[1126], 
    normalizedWires[1125], normalizedWires[1124], normalizedWires[1123], normalizedWires[1122], 
    normalizedWires[1121], normalizedWires[1120], normalizedWires[1119], normalizedWires[1118], 
    normalizedWires[1117], normalizedWires[1116], normalizedWires[1115], normalizedWires[1114], 
    normalizedWires[1113], normalizedWires[1112], normalizedWires[1111], normalizedWires[1110], 
    normalizedWires[1109], normalizedWires[1108], normalizedWires[1107], normalizedWires[1106], 
    normalizedWires[1105], uc_803, uc_804, uc_805, uc_806, uc_807, uc_808, uc_809, 
    uc_810, uc_811, uc_812, uc_813, uc_814, uc_815, uc_816, uc_817, uc_818, uc_819}));
CSAlike__1_1259 genblk2_6_parallelAdderStage1 (.carry ({uc_525, uc_526, uc_527, uc_528, 
    uc_529, uc_530, uc_531, uc_532, uc_533, uc_534, uc_535, uc_536, uc_537, \intermediateWiresStage1[13][50] , 
    \intermediateWiresStage1[13][49] , \intermediateWiresStage1[13][48] , \intermediateWiresStage1[13][47] , 
    \intermediateWiresStage1[13][46] , \intermediateWiresStage1[13][45] , \intermediateWiresStage1[13][44] , 
    \intermediateWiresStage1[13][43] , \intermediateWiresStage1[13][42] , \intermediateWiresStage1[13][41] , 
    \intermediateWiresStage1[13][40] , \intermediateWiresStage1[13][39] , \intermediateWiresStage1[13][38] , 
    \intermediateWiresStage1[13][37] , \intermediateWiresStage1[13][36] , \intermediateWiresStage1[13][35] , 
    \intermediateWiresStage1[13][34] , \intermediateWiresStage1[13][33] , \intermediateWiresStage1[13][32] , 
    \intermediateWiresStage1[13][31] , \intermediateWiresStage1[13][30] , \intermediateWiresStage1[13][29] , 
    \intermediateWiresStage1[13][28] , \intermediateWiresStage1[13][27] , \intermediateWiresStage1[13][26] , 
    \intermediateWiresStage1[13][25] , \intermediateWiresStage1[13][24] , \intermediateWiresStage1[13][23] , 
    \intermediateWiresStage1[13][22] , \intermediateWiresStage1[13][21] , \intermediateWiresStage1[13][20] , 
    uc_538, uc_539, uc_540, uc_541, uc_542, uc_543, uc_544, uc_545, uc_546, uc_547, 
    uc_548, uc_549, uc_550, uc_551, uc_552, uc_553, uc_554, uc_555, uc_556, uc_557})
    , .result ({uc_492, uc_493, uc_494, uc_495, uc_496, uc_497, uc_498, uc_499, uc_500, 
    uc_501, uc_502, uc_503, uc_504, uc_505, \intermediateWiresStage1[12][49] , \intermediateWiresStage1[12][48] , 
    \intermediateWiresStage1[12][47] , \intermediateWiresStage1[12][46] , \intermediateWiresStage1[12][45] , 
    \intermediateWiresStage1[12][44] , \intermediateWiresStage1[12][43] , \intermediateWiresStage1[12][42] , 
    \intermediateWiresStage1[12][41] , \intermediateWiresStage1[12][40] , \intermediateWiresStage1[12][39] , 
    \intermediateWiresStage1[12][38] , \intermediateWiresStage1[12][37] , \intermediateWiresStage1[12][36] , 
    \intermediateWiresStage1[12][35] , \intermediateWiresStage1[12][34] , \intermediateWiresStage1[12][33] , 
    \intermediateWiresStage1[12][32] , \intermediateWiresStage1[12][31] , \intermediateWiresStage1[12][30] , 
    \intermediateWiresStage1[12][29] , \intermediateWiresStage1[12][28] , \intermediateWiresStage1[12][27] , 
    \intermediateWiresStage1[12][26] , \intermediateWiresStage1[12][25] , \intermediateWiresStage1[12][24] , 
    \intermediateWiresStage1[12][23] , \intermediateWiresStage1[12][22] , \intermediateWiresStage1[12][21] , 
    \intermediateWiresStage1[12][20] , \intermediateWiresStage1[12][19] , uc_506, 
    uc_507, uc_508, uc_509, uc_510, uc_511, uc_512, uc_513, uc_514, uc_515, uc_516, 
    uc_517, uc_518, uc_519, uc_520, uc_521, uc_522, uc_523, uc_524}), .A ({1'b0 , 
    uc_558, uc_559, uc_560, uc_561, uc_562, uc_563, uc_564, uc_565, uc_566, uc_567, 
    uc_568, uc_569, uc_570, uc_571, normalizedWires[1200], normalizedWires[1199], 
    normalizedWires[1198], normalizedWires[1197], normalizedWires[1196], normalizedWires[1195], 
    normalizedWires[1194], normalizedWires[1193], normalizedWires[1192], normalizedWires[1191], 
    normalizedWires[1190], normalizedWires[1189], normalizedWires[1188], normalizedWires[1187], 
    normalizedWires[1186], normalizedWires[1185], normalizedWires[1184], normalizedWires[1183], 
    normalizedWires[1182], normalizedWires[1181], normalizedWires[1180], normalizedWires[1179], 
    normalizedWires[1178], normalizedWires[1177], normalizedWires[1176], normalizedWires[1175], 
    normalizedWires[1174], normalizedWires[1173], normalizedWires[1172], normalizedWires[1171], 
    uc_572, uc_573, uc_574, uc_575, uc_576, uc_577, uc_578, uc_579, uc_580, uc_581, 
    uc_582, uc_583, uc_584, uc_585, uc_586, uc_587, uc_588, uc_589, uc_590}), .B ({
    1'b0 , uc_591, uc_592, uc_593, uc_594, uc_595, uc_596, uc_597, uc_598, uc_599, 
    uc_600, uc_601, uc_602, uc_603, normalizedWires[1265], normalizedWires[1264], 
    normalizedWires[1263], normalizedWires[1262], normalizedWires[1261], normalizedWires[1260], 
    normalizedWires[1259], normalizedWires[1258], normalizedWires[1257], normalizedWires[1256], 
    normalizedWires[1255], normalizedWires[1254], normalizedWires[1253], normalizedWires[1252], 
    normalizedWires[1251], normalizedWires[1250], normalizedWires[1249], normalizedWires[1248], 
    normalizedWires[1247], normalizedWires[1246], normalizedWires[1245], normalizedWires[1244], 
    normalizedWires[1243], normalizedWires[1242], normalizedWires[1241], normalizedWires[1240], 
    normalizedWires[1239], normalizedWires[1238], normalizedWires[1237], normalizedWires[1236], 
    normalizedWires[1235], uc_604, uc_605, uc_606, uc_607, uc_608, uc_609, uc_610, 
    uc_611, uc_612, uc_613, uc_614, uc_615, uc_616, uc_617, uc_618, uc_619, uc_620, 
    uc_621, uc_622}), .C ({1'b0 , uc_623, uc_624, uc_625, uc_626, uc_627, uc_628, 
    uc_629, uc_630, uc_631, uc_632, uc_633, uc_634, uc_635, normalizedWires[1329], 
    normalizedWires[1328], normalizedWires[1327], normalizedWires[1326], normalizedWires[1325], 
    normalizedWires[1324], normalizedWires[1323], normalizedWires[1322], normalizedWires[1321], 
    normalizedWires[1320], normalizedWires[1319], normalizedWires[1318], normalizedWires[1317], 
    normalizedWires[1316], normalizedWires[1315], normalizedWires[1314], normalizedWires[1313], 
    normalizedWires[1312], normalizedWires[1311], normalizedWires[1310], normalizedWires[1309], 
    normalizedWires[1308], normalizedWires[1307], normalizedWires[1306], normalizedWires[1305], 
    normalizedWires[1304], normalizedWires[1303], normalizedWires[1302], normalizedWires[1301], 
    normalizedWires[1300], uc_636, uc_637, uc_638, uc_639, uc_640, uc_641, uc_642, 
    uc_643, uc_644, uc_645, uc_646, uc_647, uc_648, uc_649, uc_650, uc_651, uc_652, 
    uc_653, uc_654, uc_655}));
CSAlike__1_1006 genblk2_7_parallelAdderStage1 (.carry ({uc_361, uc_362, uc_363, uc_364, 
    uc_365, uc_366, uc_367, uc_368, uc_369, uc_370, \intermediateWiresStage1[15][53] , 
    \intermediateWiresStage1[15][52] , \intermediateWiresStage1[15][51] , \intermediateWiresStage1[15][50] , 
    \intermediateWiresStage1[15][49] , \intermediateWiresStage1[15][48] , \intermediateWiresStage1[15][47] , 
    \intermediateWiresStage1[15][46] , \intermediateWiresStage1[15][45] , \intermediateWiresStage1[15][44] , 
    \intermediateWiresStage1[15][43] , \intermediateWiresStage1[15][42] , \intermediateWiresStage1[15][41] , 
    \intermediateWiresStage1[15][40] , \intermediateWiresStage1[15][39] , \intermediateWiresStage1[15][38] , 
    \intermediateWiresStage1[15][37] , \intermediateWiresStage1[15][36] , \intermediateWiresStage1[15][35] , 
    \intermediateWiresStage1[15][34] , \intermediateWiresStage1[15][33] , \intermediateWiresStage1[15][32] , 
    \intermediateWiresStage1[15][31] , \intermediateWiresStage1[15][30] , \intermediateWiresStage1[15][29] , 
    \intermediateWiresStage1[15][28] , \intermediateWiresStage1[15][27] , \intermediateWiresStage1[15][26] , 
    \intermediateWiresStage1[15][25] , \intermediateWiresStage1[15][24] , \intermediateWiresStage1[15][23] , 
    uc_371, uc_372, uc_373, uc_374, uc_375, uc_376, uc_377, uc_378, uc_379, uc_380, 
    uc_381, uc_382, uc_383, uc_384, uc_385, uc_386, uc_387, uc_388, uc_389, uc_390, 
    uc_391, uc_392, uc_393}), .result ({uc_328, uc_329, uc_330, uc_331, uc_332, uc_333, 
    uc_334, uc_335, uc_336, uc_337, uc_338, \intermediateWiresStage1[14][52] , \intermediateWiresStage1[14][51] , 
    \intermediateWiresStage1[14][50] , \intermediateWiresStage1[14][49] , \intermediateWiresStage1[14][48] , 
    \intermediateWiresStage1[14][47] , \intermediateWiresStage1[14][46] , \intermediateWiresStage1[14][45] , 
    \intermediateWiresStage1[14][44] , \intermediateWiresStage1[14][43] , \intermediateWiresStage1[14][42] , 
    \intermediateWiresStage1[14][41] , \intermediateWiresStage1[14][40] , \intermediateWiresStage1[14][39] , 
    \intermediateWiresStage1[14][38] , \intermediateWiresStage1[14][37] , \intermediateWiresStage1[14][36] , 
    \intermediateWiresStage1[14][35] , \intermediateWiresStage1[14][34] , \intermediateWiresStage1[14][33] , 
    \intermediateWiresStage1[14][32] , \intermediateWiresStage1[14][31] , \intermediateWiresStage1[14][30] , 
    \intermediateWiresStage1[14][29] , \intermediateWiresStage1[14][28] , \intermediateWiresStage1[14][27] , 
    \intermediateWiresStage1[14][26] , \intermediateWiresStage1[14][25] , \intermediateWiresStage1[14][24] , 
    \intermediateWiresStage1[14][23] , \intermediateWiresStage1[14][22] , uc_339, 
    uc_340, uc_341, uc_342, uc_343, uc_344, uc_345, uc_346, uc_347, uc_348, uc_349, 
    uc_350, uc_351, uc_352, uc_353, uc_354, uc_355, uc_356, uc_357, uc_358, uc_359, 
    uc_360}), .A ({1'b0 , uc_394, uc_395, uc_396, uc_397, uc_398, uc_399, uc_400, 
    uc_401, uc_402, uc_403, uc_404, normalizedWires[1395], normalizedWires[1394], 
    normalizedWires[1393], normalizedWires[1392], normalizedWires[1391], normalizedWires[1390], 
    normalizedWires[1389], normalizedWires[1388], normalizedWires[1387], normalizedWires[1386], 
    normalizedWires[1385], normalizedWires[1384], normalizedWires[1383], normalizedWires[1382], 
    normalizedWires[1381], normalizedWires[1380], normalizedWires[1379], normalizedWires[1378], 
    normalizedWires[1377], normalizedWires[1376], normalizedWires[1375], normalizedWires[1374], 
    normalizedWires[1373], normalizedWires[1372], normalizedWires[1371], normalizedWires[1370], 
    normalizedWires[1369], normalizedWires[1368], normalizedWires[1367], normalizedWires[1366], 
    uc_405, uc_406, uc_407, uc_408, uc_409, uc_410, uc_411, uc_412, uc_413, uc_414, 
    uc_415, uc_416, uc_417, uc_418, uc_419, uc_420, uc_421, uc_422, uc_423, uc_424, 
    uc_425, uc_426}), .B ({1'b0 , uc_427, uc_428, uc_429, uc_430, uc_431, uc_432, 
    uc_433, uc_434, uc_435, uc_436, normalizedWires[1460], normalizedWires[1459], 
    normalizedWires[1458], normalizedWires[1457], normalizedWires[1456], normalizedWires[1455], 
    normalizedWires[1454], normalizedWires[1453], normalizedWires[1452], normalizedWires[1451], 
    normalizedWires[1450], normalizedWires[1449], normalizedWires[1448], normalizedWires[1447], 
    normalizedWires[1446], normalizedWires[1445], normalizedWires[1444], normalizedWires[1443], 
    normalizedWires[1442], normalizedWires[1441], normalizedWires[1440], normalizedWires[1439], 
    normalizedWires[1438], normalizedWires[1437], normalizedWires[1436], normalizedWires[1435], 
    normalizedWires[1434], normalizedWires[1433], normalizedWires[1432], normalizedWires[1431], 
    normalizedWires[1430], uc_437, uc_438, uc_439, uc_440, uc_441, uc_442, uc_443, 
    uc_444, uc_445, uc_446, uc_447, uc_448, uc_449, uc_450, uc_451, uc_452, uc_453, 
    uc_454, uc_455, uc_456, uc_457, uc_458}), .C ({1'b0 , uc_459, uc_460, uc_461, 
    uc_462, uc_463, uc_464, uc_465, uc_466, uc_467, uc_468, normalizedWires[1524], 
    normalizedWires[1523], normalizedWires[1522], normalizedWires[1521], normalizedWires[1520], 
    normalizedWires[1519], normalizedWires[1518], normalizedWires[1517], normalizedWires[1516], 
    normalizedWires[1515], normalizedWires[1514], normalizedWires[1513], normalizedWires[1512], 
    normalizedWires[1511], normalizedWires[1510], normalizedWires[1509], normalizedWires[1508], 
    normalizedWires[1507], normalizedWires[1506], normalizedWires[1505], normalizedWires[1504], 
    normalizedWires[1503], normalizedWires[1502], normalizedWires[1501], normalizedWires[1500], 
    normalizedWires[1499], normalizedWires[1498], normalizedWires[1497], normalizedWires[1496], 
    normalizedWires[1495], uc_469, uc_470, uc_471, uc_472, uc_473, uc_474, uc_475, 
    uc_476, uc_477, uc_478, uc_479, uc_480, uc_481, uc_482, uc_483, uc_484, uc_485, 
    uc_486, uc_487, uc_488, uc_489, uc_490, uc_491}));
CSAlike__1_753 genblk2_8_parallelAdderStage1 (.carry ({uc_197, uc_198, uc_199, uc_200, 
    uc_201, uc_202, uc_203, \intermediateWiresStage1[17][56] , \intermediateWiresStage1[17][55] , 
    \intermediateWiresStage1[17][54] , \intermediateWiresStage1[17][53] , \intermediateWiresStage1[17][52] , 
    \intermediateWiresStage1[17][51] , \intermediateWiresStage1[17][50] , \intermediateWiresStage1[17][49] , 
    \intermediateWiresStage1[17][48] , \intermediateWiresStage1[17][47] , \intermediateWiresStage1[17][46] , 
    \intermediateWiresStage1[17][45] , \intermediateWiresStage1[17][44] , \intermediateWiresStage1[17][43] , 
    \intermediateWiresStage1[17][42] , \intermediateWiresStage1[17][41] , \intermediateWiresStage1[17][40] , 
    \intermediateWiresStage1[17][39] , \intermediateWiresStage1[17][38] , \intermediateWiresStage1[17][37] , 
    \intermediateWiresStage1[17][36] , \intermediateWiresStage1[17][35] , \intermediateWiresStage1[17][34] , 
    \intermediateWiresStage1[17][33] , \intermediateWiresStage1[17][32] , \intermediateWiresStage1[17][31] , 
    \intermediateWiresStage1[17][30] , \intermediateWiresStage1[17][29] , \intermediateWiresStage1[17][28] , 
    \intermediateWiresStage1[17][27] , \intermediateWiresStage1[17][26] , uc_204, 
    uc_205, uc_206, uc_207, uc_208, uc_209, uc_210, uc_211, uc_212, uc_213, uc_214, 
    uc_215, uc_216, uc_217, uc_218, uc_219, uc_220, uc_221, uc_222, uc_223, uc_224, 
    uc_225, uc_226, uc_227, uc_228, uc_229}), .result ({uc_164, uc_165, uc_166, uc_167, 
    uc_168, uc_169, uc_170, uc_171, \intermediateWiresStage1[16][55] , \intermediateWiresStage1[16][54] , 
    \intermediateWiresStage1[16][53] , \intermediateWiresStage1[16][52] , \intermediateWiresStage1[16][51] , 
    \intermediateWiresStage1[16][50] , \intermediateWiresStage1[16][49] , \intermediateWiresStage1[16][48] , 
    \intermediateWiresStage1[16][47] , \intermediateWiresStage1[16][46] , \intermediateWiresStage1[16][45] , 
    \intermediateWiresStage1[16][44] , \intermediateWiresStage1[16][43] , \intermediateWiresStage1[16][42] , 
    \intermediateWiresStage1[16][41] , \intermediateWiresStage1[16][40] , \intermediateWiresStage1[16][39] , 
    \intermediateWiresStage1[16][38] , \intermediateWiresStage1[16][37] , \intermediateWiresStage1[16][36] , 
    \intermediateWiresStage1[16][35] , \intermediateWiresStage1[16][34] , \intermediateWiresStage1[16][33] , 
    \intermediateWiresStage1[16][32] , \intermediateWiresStage1[16][31] , \intermediateWiresStage1[16][30] , 
    \intermediateWiresStage1[16][29] , \intermediateWiresStage1[16][28] , \intermediateWiresStage1[16][27] , 
    \intermediateWiresStage1[16][26] , \intermediateWiresStage1[16][25] , uc_172, 
    uc_173, uc_174, uc_175, uc_176, uc_177, uc_178, uc_179, uc_180, uc_181, uc_182, 
    uc_183, uc_184, uc_185, uc_186, uc_187, uc_188, uc_189, uc_190, uc_191, uc_192, 
    uc_193, uc_194, uc_195, uc_196}), .A ({1'b0 , uc_230, uc_231, uc_232, uc_233, 
    uc_234, uc_235, uc_236, uc_237, normalizedWires[1590], normalizedWires[1589], 
    normalizedWires[1588], normalizedWires[1587], normalizedWires[1586], normalizedWires[1585], 
    normalizedWires[1584], normalizedWires[1583], normalizedWires[1582], normalizedWires[1581], 
    normalizedWires[1580], normalizedWires[1579], normalizedWires[1578], normalizedWires[1577], 
    normalizedWires[1576], normalizedWires[1575], normalizedWires[1574], normalizedWires[1573], 
    normalizedWires[1572], normalizedWires[1571], normalizedWires[1570], normalizedWires[1569], 
    normalizedWires[1568], normalizedWires[1567], normalizedWires[1566], normalizedWires[1565], 
    normalizedWires[1564], normalizedWires[1563], normalizedWires[1562], normalizedWires[1561], 
    uc_238, uc_239, uc_240, uc_241, uc_242, uc_243, uc_244, uc_245, uc_246, uc_247, 
    uc_248, uc_249, uc_250, uc_251, uc_252, uc_253, uc_254, uc_255, uc_256, uc_257, 
    uc_258, uc_259, uc_260, uc_261, uc_262}), .B ({1'b0 , uc_263, uc_264, uc_265, 
    uc_266, uc_267, uc_268, uc_269, normalizedWires[1655], normalizedWires[1654], 
    normalizedWires[1653], normalizedWires[1652], normalizedWires[1651], normalizedWires[1650], 
    normalizedWires[1649], normalizedWires[1648], normalizedWires[1647], normalizedWires[1646], 
    normalizedWires[1645], normalizedWires[1644], normalizedWires[1643], normalizedWires[1642], 
    normalizedWires[1641], normalizedWires[1640], normalizedWires[1639], normalizedWires[1638], 
    normalizedWires[1637], normalizedWires[1636], normalizedWires[1635], normalizedWires[1634], 
    normalizedWires[1633], normalizedWires[1632], normalizedWires[1631], normalizedWires[1630], 
    normalizedWires[1629], normalizedWires[1628], normalizedWires[1627], normalizedWires[1626], 
    normalizedWires[1625], uc_270, uc_271, uc_272, uc_273, uc_274, uc_275, uc_276, 
    uc_277, uc_278, uc_279, uc_280, uc_281, uc_282, uc_283, uc_284, uc_285, uc_286, 
    uc_287, uc_288, uc_289, uc_290, uc_291, uc_292, uc_293, uc_294}), .C ({1'b0 , 
    uc_295, uc_296, uc_297, uc_298, uc_299, uc_300, uc_301, normalizedWires[1719], 
    normalizedWires[1718], normalizedWires[1717], normalizedWires[1716], normalizedWires[1715], 
    normalizedWires[1714], normalizedWires[1713], normalizedWires[1712], normalizedWires[1711], 
    normalizedWires[1710], normalizedWires[1709], normalizedWires[1708], normalizedWires[1707], 
    normalizedWires[1706], normalizedWires[1705], normalizedWires[1704], normalizedWires[1703], 
    normalizedWires[1702], normalizedWires[1701], normalizedWires[1700], normalizedWires[1699], 
    normalizedWires[1698], normalizedWires[1697], normalizedWires[1696], normalizedWires[1695], 
    normalizedWires[1694], normalizedWires[1693], normalizedWires[1692], normalizedWires[1691], 
    normalizedWires[1690], uc_302, uc_303, uc_304, uc_305, uc_306, uc_307, uc_308, 
    uc_309, uc_310, uc_311, uc_312, uc_313, uc_314, uc_315, uc_316, uc_317, uc_318, 
    uc_319, uc_320, uc_321, uc_322, uc_323, uc_324, uc_325, uc_326, uc_327}));
CSAlike__1_500 genblk2_9_parallelAdderStage1 (.carry ({uc_33, uc_34, uc_35, uc_36, 
    \intermediateWiresStage1[19][59] , \intermediateWiresStage1[19][58] , \intermediateWiresStage1[19][57] , 
    \intermediateWiresStage1[19][56] , \intermediateWiresStage1[19][55] , \intermediateWiresStage1[19][54] , 
    \intermediateWiresStage1[19][53] , \intermediateWiresStage1[19][52] , \intermediateWiresStage1[19][51] , 
    \intermediateWiresStage1[19][50] , \intermediateWiresStage1[19][49] , \intermediateWiresStage1[19][48] , 
    \intermediateWiresStage1[19][47] , \intermediateWiresStage1[19][46] , \intermediateWiresStage1[19][45] , 
    \intermediateWiresStage1[19][44] , \intermediateWiresStage1[19][43] , \intermediateWiresStage1[19][42] , 
    \intermediateWiresStage1[19][41] , \intermediateWiresStage1[19][40] , \intermediateWiresStage1[19][39] , 
    \intermediateWiresStage1[19][38] , \intermediateWiresStage1[19][37] , \intermediateWiresStage1[19][36] , 
    \intermediateWiresStage1[19][35] , \intermediateWiresStage1[19][34] , \intermediateWiresStage1[19][33] , 
    \intermediateWiresStage1[19][32] , \intermediateWiresStage1[19][31] , \intermediateWiresStage1[19][30] , 
    \intermediateWiresStage1[19][29] , uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, 
    uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49, uc_50, uc_51, uc_52, uc_53, 
    uc_54, uc_55, uc_56, uc_57, uc_58, uc_59, uc_60, uc_61, uc_62, uc_63, uc_64, 
    uc_65}), .result ({uc_0, uc_1, uc_2, uc_3, uc_4, \intermediateWiresStage1[18][58] , 
    \intermediateWiresStage1[18][57] , \intermediateWiresStage1[18][56] , \intermediateWiresStage1[18][55] , 
    \intermediateWiresStage1[18][54] , \intermediateWiresStage1[18][53] , \intermediateWiresStage1[18][52] , 
    \intermediateWiresStage1[18][51] , \intermediateWiresStage1[18][50] , \intermediateWiresStage1[18][49] , 
    \intermediateWiresStage1[18][48] , \intermediateWiresStage1[18][47] , \intermediateWiresStage1[18][46] , 
    \intermediateWiresStage1[18][45] , \intermediateWiresStage1[18][44] , \intermediateWiresStage1[18][43] , 
    \intermediateWiresStage1[18][42] , \intermediateWiresStage1[18][41] , \intermediateWiresStage1[18][40] , 
    \intermediateWiresStage1[18][39] , \intermediateWiresStage1[18][38] , \intermediateWiresStage1[18][37] , 
    \intermediateWiresStage1[18][36] , \intermediateWiresStage1[18][35] , \intermediateWiresStage1[18][34] , 
    \intermediateWiresStage1[18][33] , \intermediateWiresStage1[18][32] , \intermediateWiresStage1[18][31] , 
    \intermediateWiresStage1[18][30] , \intermediateWiresStage1[18][29] , \intermediateWiresStage1[18][28] , 
    uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, 
    uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, 
    uc_28, uc_29, uc_30, uc_31, uc_32}), .A ({1'b0 , uc_66, uc_67, uc_68, uc_69, 
    uc_70, normalizedWires[1785], normalizedWires[1784], normalizedWires[1783], normalizedWires[1782], 
    normalizedWires[1781], normalizedWires[1780], normalizedWires[1779], normalizedWires[1778], 
    normalizedWires[1777], normalizedWires[1776], normalizedWires[1775], normalizedWires[1774], 
    normalizedWires[1773], normalizedWires[1772], normalizedWires[1771], normalizedWires[1770], 
    normalizedWires[1769], normalizedWires[1768], normalizedWires[1767], normalizedWires[1766], 
    normalizedWires[1765], normalizedWires[1764], normalizedWires[1763], normalizedWires[1762], 
    normalizedWires[1761], normalizedWires[1760], normalizedWires[1759], normalizedWires[1758], 
    normalizedWires[1757], normalizedWires[1756], uc_71, uc_72, uc_73, uc_74, uc_75, 
    uc_76, uc_77, uc_78, uc_79, uc_80, uc_81, uc_82, uc_83, uc_84, uc_85, uc_86, 
    uc_87, uc_88, uc_89, uc_90, uc_91, uc_92, uc_93, uc_94, uc_95, uc_96, uc_97, 
    uc_98}), .B ({1'b0 , uc_99, uc_100, uc_101, uc_102, normalizedWires[1850], normalizedWires[1849], 
    normalizedWires[1848], normalizedWires[1847], normalizedWires[1846], normalizedWires[1845], 
    normalizedWires[1844], normalizedWires[1843], normalizedWires[1842], normalizedWires[1841], 
    normalizedWires[1840], normalizedWires[1839], normalizedWires[1838], normalizedWires[1837], 
    normalizedWires[1836], normalizedWires[1835], normalizedWires[1834], normalizedWires[1833], 
    normalizedWires[1832], normalizedWires[1831], normalizedWires[1830], normalizedWires[1829], 
    normalizedWires[1828], normalizedWires[1827], normalizedWires[1826], normalizedWires[1825], 
    normalizedWires[1824], normalizedWires[1823], normalizedWires[1822], normalizedWires[1821], 
    normalizedWires[1820], uc_103, uc_104, uc_105, uc_106, uc_107, uc_108, uc_109, 
    uc_110, uc_111, uc_112, uc_113, uc_114, uc_115, uc_116, uc_117, uc_118, uc_119, 
    uc_120, uc_121, uc_122, uc_123, uc_124, uc_125, uc_126, uc_127, uc_128, uc_129, 
    uc_130}), .C ({1'b0 , uc_131, uc_132, uc_133, uc_134, normalizedWires[1914], 
    normalizedWires[1913], normalizedWires[1912], normalizedWires[1911], normalizedWires[1910], 
    normalizedWires[1909], normalizedWires[1908], normalizedWires[1907], normalizedWires[1906], 
    normalizedWires[1905], normalizedWires[1904], normalizedWires[1903], normalizedWires[1902], 
    normalizedWires[1901], normalizedWires[1900], normalizedWires[1899], normalizedWires[1898], 
    normalizedWires[1897], normalizedWires[1896], normalizedWires[1895], normalizedWires[1894], 
    normalizedWires[1893], normalizedWires[1892], normalizedWires[1891], normalizedWires[1890], 
    normalizedWires[1889], normalizedWires[1888], normalizedWires[1887], normalizedWires[1886], 
    normalizedWires[1885], uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, uc_141, 
    uc_142, uc_143, uc_144, uc_145, uc_146, uc_147, uc_148, uc_149, uc_150, uc_151, 
    uc_152, uc_153, uc_154, uc_155, uc_156, uc_157, uc_158, uc_159, uc_160, uc_161, 
    uc_162, uc_163}));

endmodule //addIntermedaiteWires

module multiplierTree (Res, OVF, A, B, clk, reset, enable);

output OVF;
output [63:0] Res;
input [31:0] A;
input [31:0] B;
input clk;
input enable;
input reset;
wire opt_ipo_n1380;
wire CLOCK_slo__sro_n2212;
wire CLOCK_slh_n3498;
wire \secondStage_carry[62] ;
wire \secondStage_carry[61] ;
wire \secondStage_carry[60] ;
wire \secondStage_carry[59] ;
wire \secondStage_carry[58] ;
wire \secondStage_carry[57] ;
wire \secondStage_carry[56] ;
wire \secondStage_carry[55] ;
wire \secondStage_carry[54] ;
wire \secondStage_carry[53] ;
wire \secondStage_carry[52] ;
wire \secondStage_carry[51] ;
wire \secondStage_carry[50] ;
wire \secondStage_carry[49] ;
wire \secondStage_carry[48] ;
wire \secondStage_carry[47] ;
wire \secondStage_carry[46] ;
wire \secondStage_carry[45] ;
wire \secondStage_carry[44] ;
wire \secondStage_carry[43] ;
wire \secondStage_carry[42] ;
wire \secondStage_carry[41] ;
wire \secondStage_carry[40] ;
wire \secondStage_carry[39] ;
wire \secondStage_carry[38] ;
wire \secondStage_carry[37] ;
wire \secondStage_carry[36] ;
wire \secondStage_carry[35] ;
wire \secondStage_carry[34] ;
wire \secondStage_carry[33] ;
wire \secondStage_carry[32] ;
wire \secondStage_carry[31] ;
wire \secondStage_carry[30] ;
wire \secondStage_carry[29] ;
wire \secondStage_carry[28] ;
wire \secondStage_carry[27] ;
wire \secondStage_carry[26] ;
wire \secondStage_carry[25] ;
wire \secondStage_carry[24] ;
wire \secondStage_carry[23] ;
wire \secondStage_carry[22] ;
wire \secondStage_carry[21] ;
wire \secondStage_carry[20] ;
wire \secondStage_carry[19] ;
wire \secondStage_carry[18] ;
wire \secondStage_carry[17] ;
wire \secondStage_carry[16] ;
wire \secondStage_carry[15] ;
wire \secondStage_carry[14] ;
wire \secondStage_carry[13] ;
wire \secondStage_carry[12] ;
wire \secondStage_carry[11] ;
wire \secondStage_carry[10] ;
wire \secondStage_carry[9] ;
wire \secondStage_Res[61] ;
wire \secondStage_Res[60] ;
wire \secondStage_Res[59] ;
wire \secondStage_Res[58] ;
wire \secondStage_Res[57] ;
wire \secondStage_Res[56] ;
wire \secondStage_Res[55] ;
wire \secondStage_Res[54] ;
wire \secondStage_Res[53] ;
wire \secondStage_Res[52] ;
wire \secondStage_Res[51] ;
wire \secondStage_Res[50] ;
wire \secondStage_Res[49] ;
wire \secondStage_Res[48] ;
wire \secondStage_Res[47] ;
wire \secondStage_Res[46] ;
wire \secondStage_Res[45] ;
wire \secondStage_Res[44] ;
wire \secondStage_Res[43] ;
wire \secondStage_Res[42] ;
wire \secondStage_Res[41] ;
wire \secondStage_Res[40] ;
wire \secondStage_Res[39] ;
wire \secondStage_Res[38] ;
wire \secondStage_Res[37] ;
wire \secondStage_Res[36] ;
wire \secondStage_Res[35] ;
wire \secondStage_Res[34] ;
wire \secondStage_Res[33] ;
wire \secondStage_Res[32] ;
wire \secondStage_Res[31] ;
wire \secondStage_Res[30] ;
wire \secondStage_Res[29] ;
wire \secondStage_Res[28] ;
wire \secondStage_Res[27] ;
wire \secondStage_Res[26] ;
wire \secondStage_Res[25] ;
wire \secondStage_Res[24] ;
wire \secondStage_Res[23] ;
wire \secondStage_Res[22] ;
wire \secondStage_Res[21] ;
wire \secondStage_Res[20] ;
wire \secondStage_Res[19] ;
wire \secondStage_Res[18] ;
wire \secondStage_Res[17] ;
wire \secondStage_Res[16] ;
wire \secondStage_Res[15] ;
wire \secondStage_Res[14] ;
wire \secondStage_Res[13] ;
wire \secondStage_Res[12] ;
wire \secondStage_Res[11] ;
wire \secondStage_Res[10] ;
wire \secondStage_Res[9] ;
wire \secondStage_Res[8] ;
wire \secondStage_Res[7] ;
wire \secondStage_Res[6] ;
wire \secondStage_Res[5] ;
wire \secondStage_Res[4] ;
wire \secondStage_Res[3] ;
wire \secondStage_Res[2] ;
wire \secondStage_Res[1] ;
wire n_0_316;
wire \normalizedWires[2045] ;
wire \normalizedWires[2044] ;
wire \normalizedWires[2043] ;
wire \normalizedWires[2042] ;
wire \normalizedWires[2041] ;
wire \normalizedWires[2040] ;
wire \normalizedWires[2039] ;
wire \normalizedWires[2038] ;
wire \normalizedWires[2037] ;
wire \normalizedWires[2036] ;
wire \normalizedWires[2035] ;
wire \normalizedWires[2034] ;
wire \normalizedWires[2033] ;
wire \normalizedWires[2032] ;
wire \normalizedWires[2031] ;
wire \normalizedWires[2030] ;
wire \normalizedWires[2029] ;
wire \normalizedWires[2028] ;
wire \normalizedWires[2027] ;
wire \normalizedWires[2026] ;
wire \normalizedWires[2025] ;
wire \normalizedWires[2024] ;
wire \normalizedWires[2023] ;
wire \normalizedWires[2022] ;
wire \normalizedWires[2021] ;
wire \normalizedWires[2020] ;
wire \normalizedWires[2019] ;
wire \normalizedWires[2018] ;
wire \normalizedWires[2017] ;
wire \normalizedWires[2016] ;
wire \normalizedWires[2015] ;
wire \normalizedWires[1980] ;
wire \normalizedWires[1979] ;
wire \normalizedWires[1978] ;
wire \normalizedWires[1977] ;
wire \normalizedWires[1976] ;
wire \normalizedWires[1975] ;
wire \normalizedWires[1974] ;
wire \normalizedWires[1973] ;
wire \normalizedWires[1972] ;
wire \normalizedWires[1971] ;
wire \normalizedWires[1970] ;
wire \normalizedWires[1969] ;
wire \normalizedWires[1968] ;
wire \normalizedWires[1967] ;
wire \normalizedWires[1966] ;
wire \normalizedWires[1965] ;
wire \normalizedWires[1964] ;
wire \normalizedWires[1963] ;
wire \normalizedWires[1962] ;
wire \normalizedWires[1961] ;
wire \normalizedWires[1960] ;
wire \normalizedWires[1959] ;
wire \normalizedWires[1958] ;
wire \normalizedWires[1957] ;
wire \normalizedWires[1956] ;
wire \normalizedWires[1955] ;
wire \normalizedWires[1954] ;
wire \normalizedWires[1953] ;
wire \normalizedWires[1952] ;
wire \normalizedWires[1951] ;
wire \normalizedWires[1950] ;
wire \normalizedWires[1915] ;
wire \normalizedWires[1914] ;
wire \normalizedWires[1913] ;
wire \normalizedWires[1912] ;
wire \normalizedWires[1911] ;
wire \normalizedWires[1910] ;
wire \normalizedWires[1909] ;
wire \normalizedWires[1908] ;
wire \normalizedWires[1907] ;
wire \normalizedWires[1906] ;
wire \normalizedWires[1905] ;
wire \normalizedWires[1904] ;
wire \normalizedWires[1903] ;
wire \normalizedWires[1902] ;
wire \normalizedWires[1901] ;
wire \normalizedWires[1900] ;
wire \normalizedWires[1899] ;
wire \normalizedWires[1898] ;
wire \normalizedWires[1897] ;
wire \normalizedWires[1896] ;
wire \normalizedWires[1895] ;
wire \normalizedWires[1894] ;
wire \normalizedWires[1893] ;
wire \normalizedWires[1892] ;
wire \normalizedWires[1891] ;
wire \normalizedWires[1890] ;
wire \normalizedWires[1889] ;
wire \normalizedWires[1888] ;
wire \normalizedWires[1887] ;
wire \normalizedWires[1886] ;
wire \normalizedWires[1885] ;
wire \normalizedWires[1850] ;
wire \normalizedWires[1849] ;
wire \normalizedWires[1848] ;
wire \normalizedWires[1847] ;
wire \normalizedWires[1846] ;
wire \normalizedWires[1845] ;
wire \normalizedWires[1844] ;
wire \normalizedWires[1843] ;
wire \normalizedWires[1842] ;
wire \normalizedWires[1841] ;
wire \normalizedWires[1840] ;
wire \normalizedWires[1839] ;
wire \normalizedWires[1838] ;
wire \normalizedWires[1837] ;
wire \normalizedWires[1836] ;
wire \normalizedWires[1835] ;
wire \normalizedWires[1834] ;
wire \normalizedWires[1833] ;
wire \normalizedWires[1832] ;
wire \normalizedWires[1831] ;
wire \normalizedWires[1830] ;
wire \normalizedWires[1829] ;
wire \normalizedWires[1828] ;
wire \normalizedWires[1827] ;
wire \normalizedWires[1826] ;
wire \normalizedWires[1825] ;
wire \normalizedWires[1824] ;
wire \normalizedWires[1823] ;
wire \normalizedWires[1822] ;
wire \normalizedWires[1821] ;
wire \normalizedWires[1820] ;
wire \normalizedWires[1785] ;
wire \normalizedWires[1784] ;
wire \normalizedWires[1783] ;
wire \normalizedWires[1782] ;
wire \normalizedWires[1781] ;
wire \normalizedWires[1780] ;
wire \normalizedWires[1779] ;
wire \normalizedWires[1778] ;
wire \normalizedWires[1777] ;
wire \normalizedWires[1776] ;
wire \normalizedWires[1775] ;
wire \normalizedWires[1774] ;
wire \normalizedWires[1773] ;
wire \normalizedWires[1772] ;
wire \normalizedWires[1771] ;
wire \normalizedWires[1770] ;
wire \normalizedWires[1769] ;
wire \normalizedWires[1768] ;
wire \normalizedWires[1767] ;
wire \normalizedWires[1766] ;
wire \normalizedWires[1765] ;
wire \normalizedWires[1764] ;
wire \normalizedWires[1763] ;
wire \normalizedWires[1762] ;
wire \normalizedWires[1761] ;
wire \normalizedWires[1760] ;
wire \normalizedWires[1759] ;
wire \normalizedWires[1758] ;
wire \normalizedWires[1757] ;
wire \normalizedWires[1756] ;
wire \normalizedWires[1755] ;
wire \normalizedWires[1720] ;
wire \normalizedWires[1719] ;
wire \normalizedWires[1718] ;
wire \normalizedWires[1717] ;
wire \normalizedWires[1716] ;
wire \normalizedWires[1715] ;
wire \normalizedWires[1714] ;
wire \normalizedWires[1713] ;
wire \normalizedWires[1712] ;
wire \normalizedWires[1711] ;
wire \normalizedWires[1710] ;
wire \normalizedWires[1709] ;
wire \normalizedWires[1708] ;
wire \normalizedWires[1707] ;
wire \normalizedWires[1706] ;
wire \normalizedWires[1705] ;
wire \normalizedWires[1704] ;
wire \normalizedWires[1703] ;
wire \normalizedWires[1702] ;
wire \normalizedWires[1701] ;
wire \normalizedWires[1700] ;
wire \normalizedWires[1699] ;
wire \normalizedWires[1698] ;
wire \normalizedWires[1697] ;
wire \normalizedWires[1696] ;
wire \normalizedWires[1695] ;
wire \normalizedWires[1694] ;
wire \normalizedWires[1693] ;
wire \normalizedWires[1692] ;
wire \normalizedWires[1691] ;
wire \normalizedWires[1690] ;
wire \normalizedWires[1655] ;
wire \normalizedWires[1654] ;
wire \normalizedWires[1653] ;
wire \normalizedWires[1652] ;
wire \normalizedWires[1651] ;
wire \normalizedWires[1650] ;
wire \normalizedWires[1649] ;
wire \normalizedWires[1648] ;
wire \normalizedWires[1647] ;
wire \normalizedWires[1646] ;
wire \normalizedWires[1645] ;
wire \normalizedWires[1644] ;
wire \normalizedWires[1643] ;
wire \normalizedWires[1642] ;
wire \normalizedWires[1641] ;
wire \normalizedWires[1640] ;
wire \normalizedWires[1639] ;
wire \normalizedWires[1638] ;
wire \normalizedWires[1637] ;
wire \normalizedWires[1636] ;
wire \normalizedWires[1635] ;
wire \normalizedWires[1634] ;
wire \normalizedWires[1633] ;
wire \normalizedWires[1632] ;
wire \normalizedWires[1631] ;
wire \normalizedWires[1630] ;
wire \normalizedWires[1629] ;
wire \normalizedWires[1628] ;
wire \normalizedWires[1627] ;
wire \normalizedWires[1626] ;
wire \normalizedWires[1625] ;
wire \normalizedWires[1590] ;
wire \normalizedWires[1589] ;
wire \normalizedWires[1588] ;
wire \normalizedWires[1587] ;
wire \normalizedWires[1586] ;
wire \normalizedWires[1585] ;
wire \normalizedWires[1584] ;
wire \normalizedWires[1583] ;
wire \normalizedWires[1582] ;
wire \normalizedWires[1581] ;
wire \normalizedWires[1580] ;
wire \normalizedWires[1579] ;
wire \normalizedWires[1578] ;
wire \normalizedWires[1577] ;
wire \normalizedWires[1576] ;
wire \normalizedWires[1575] ;
wire \normalizedWires[1574] ;
wire \normalizedWires[1573] ;
wire \normalizedWires[1572] ;
wire \normalizedWires[1571] ;
wire \normalizedWires[1570] ;
wire \normalizedWires[1569] ;
wire \normalizedWires[1568] ;
wire \normalizedWires[1567] ;
wire \normalizedWires[1566] ;
wire \normalizedWires[1565] ;
wire \normalizedWires[1564] ;
wire \normalizedWires[1563] ;
wire \normalizedWires[1562] ;
wire \normalizedWires[1561] ;
wire \normalizedWires[1560] ;
wire \normalizedWires[1525] ;
wire \normalizedWires[1524] ;
wire \normalizedWires[1523] ;
wire \normalizedWires[1522] ;
wire \normalizedWires[1521] ;
wire \normalizedWires[1520] ;
wire \normalizedWires[1519] ;
wire \normalizedWires[1518] ;
wire \normalizedWires[1517] ;
wire \normalizedWires[1516] ;
wire \normalizedWires[1515] ;
wire \normalizedWires[1514] ;
wire \normalizedWires[1513] ;
wire \normalizedWires[1512] ;
wire \normalizedWires[1511] ;
wire \normalizedWires[1510] ;
wire \normalizedWires[1509] ;
wire \normalizedWires[1508] ;
wire \normalizedWires[1507] ;
wire \normalizedWires[1506] ;
wire \normalizedWires[1505] ;
wire \normalizedWires[1504] ;
wire \normalizedWires[1503] ;
wire \normalizedWires[1502] ;
wire \normalizedWires[1501] ;
wire \normalizedWires[1500] ;
wire \normalizedWires[1499] ;
wire \normalizedWires[1498] ;
wire \normalizedWires[1497] ;
wire \normalizedWires[1496] ;
wire \normalizedWires[1495] ;
wire \normalizedWires[1460] ;
wire \normalizedWires[1459] ;
wire \normalizedWires[1458] ;
wire \normalizedWires[1457] ;
wire \normalizedWires[1456] ;
wire \normalizedWires[1455] ;
wire \normalizedWires[1454] ;
wire \normalizedWires[1453] ;
wire \normalizedWires[1452] ;
wire \normalizedWires[1451] ;
wire \normalizedWires[1450] ;
wire \normalizedWires[1449] ;
wire \normalizedWires[1448] ;
wire \normalizedWires[1447] ;
wire \normalizedWires[1446] ;
wire \normalizedWires[1445] ;
wire \normalizedWires[1444] ;
wire \normalizedWires[1443] ;
wire \normalizedWires[1442] ;
wire \normalizedWires[1441] ;
wire \normalizedWires[1440] ;
wire \normalizedWires[1439] ;
wire \normalizedWires[1438] ;
wire \normalizedWires[1437] ;
wire \normalizedWires[1436] ;
wire \normalizedWires[1435] ;
wire \normalizedWires[1434] ;
wire \normalizedWires[1433] ;
wire \normalizedWires[1432] ;
wire \normalizedWires[1431] ;
wire \normalizedWires[1430] ;
wire \normalizedWires[1395] ;
wire \normalizedWires[1394] ;
wire \normalizedWires[1393] ;
wire \normalizedWires[1392] ;
wire \normalizedWires[1391] ;
wire \normalizedWires[1390] ;
wire \normalizedWires[1389] ;
wire \normalizedWires[1388] ;
wire \normalizedWires[1387] ;
wire \normalizedWires[1386] ;
wire \normalizedWires[1385] ;
wire \normalizedWires[1384] ;
wire \normalizedWires[1383] ;
wire \normalizedWires[1382] ;
wire \normalizedWires[1381] ;
wire \normalizedWires[1380] ;
wire \normalizedWires[1379] ;
wire \normalizedWires[1378] ;
wire \normalizedWires[1377] ;
wire \normalizedWires[1376] ;
wire \normalizedWires[1375] ;
wire \normalizedWires[1374] ;
wire \normalizedWires[1373] ;
wire \normalizedWires[1372] ;
wire \normalizedWires[1371] ;
wire \normalizedWires[1370] ;
wire \normalizedWires[1369] ;
wire \normalizedWires[1368] ;
wire \normalizedWires[1367] ;
wire \normalizedWires[1366] ;
wire \normalizedWires[1365] ;
wire \normalizedWires[1330] ;
wire \normalizedWires[1329] ;
wire \normalizedWires[1328] ;
wire \normalizedWires[1327] ;
wire \normalizedWires[1326] ;
wire \normalizedWires[1325] ;
wire \normalizedWires[1324] ;
wire \normalizedWires[1323] ;
wire \normalizedWires[1322] ;
wire \normalizedWires[1321] ;
wire \normalizedWires[1320] ;
wire \normalizedWires[1319] ;
wire \normalizedWires[1318] ;
wire \normalizedWires[1317] ;
wire \normalizedWires[1316] ;
wire \normalizedWires[1315] ;
wire \normalizedWires[1314] ;
wire \normalizedWires[1313] ;
wire \normalizedWires[1312] ;
wire \normalizedWires[1311] ;
wire \normalizedWires[1310] ;
wire \normalizedWires[1309] ;
wire \normalizedWires[1308] ;
wire \normalizedWires[1307] ;
wire \normalizedWires[1306] ;
wire \normalizedWires[1305] ;
wire \normalizedWires[1304] ;
wire \normalizedWires[1303] ;
wire \normalizedWires[1302] ;
wire \normalizedWires[1301] ;
wire \normalizedWires[1300] ;
wire \normalizedWires[1265] ;
wire \normalizedWires[1264] ;
wire \normalizedWires[1263] ;
wire \normalizedWires[1262] ;
wire \normalizedWires[1261] ;
wire \normalizedWires[1260] ;
wire \normalizedWires[1259] ;
wire \normalizedWires[1258] ;
wire \normalizedWires[1257] ;
wire \normalizedWires[1256] ;
wire \normalizedWires[1255] ;
wire \normalizedWires[1254] ;
wire \normalizedWires[1253] ;
wire \normalizedWires[1252] ;
wire \normalizedWires[1251] ;
wire \normalizedWires[1250] ;
wire \normalizedWires[1249] ;
wire \normalizedWires[1248] ;
wire \normalizedWires[1247] ;
wire \normalizedWires[1246] ;
wire \normalizedWires[1245] ;
wire \normalizedWires[1244] ;
wire \normalizedWires[1243] ;
wire \normalizedWires[1242] ;
wire \normalizedWires[1241] ;
wire \normalizedWires[1240] ;
wire \normalizedWires[1239] ;
wire \normalizedWires[1238] ;
wire \normalizedWires[1237] ;
wire \normalizedWires[1236] ;
wire \normalizedWires[1235] ;
wire \normalizedWires[1200] ;
wire \normalizedWires[1199] ;
wire \normalizedWires[1198] ;
wire \normalizedWires[1197] ;
wire \normalizedWires[1196] ;
wire \normalizedWires[1195] ;
wire \normalizedWires[1194] ;
wire \normalizedWires[1193] ;
wire \normalizedWires[1192] ;
wire \normalizedWires[1191] ;
wire \normalizedWires[1190] ;
wire \normalizedWires[1189] ;
wire \normalizedWires[1188] ;
wire \normalizedWires[1187] ;
wire \normalizedWires[1186] ;
wire \normalizedWires[1185] ;
wire \normalizedWires[1184] ;
wire \normalizedWires[1183] ;
wire \normalizedWires[1182] ;
wire \normalizedWires[1181] ;
wire \normalizedWires[1180] ;
wire \normalizedWires[1179] ;
wire \normalizedWires[1178] ;
wire \normalizedWires[1177] ;
wire \normalizedWires[1176] ;
wire \normalizedWires[1175] ;
wire \normalizedWires[1174] ;
wire \normalizedWires[1173] ;
wire \normalizedWires[1172] ;
wire \normalizedWires[1171] ;
wire \normalizedWires[1170] ;
wire \normalizedWires[1135] ;
wire \normalizedWires[1134] ;
wire \normalizedWires[1133] ;
wire \normalizedWires[1132] ;
wire \normalizedWires[1131] ;
wire \normalizedWires[1130] ;
wire \normalizedWires[1129] ;
wire \normalizedWires[1128] ;
wire \normalizedWires[1127] ;
wire \normalizedWires[1126] ;
wire \normalizedWires[1125] ;
wire \normalizedWires[1124] ;
wire \normalizedWires[1123] ;
wire \normalizedWires[1122] ;
wire \normalizedWires[1121] ;
wire \normalizedWires[1120] ;
wire \normalizedWires[1119] ;
wire \normalizedWires[1118] ;
wire \normalizedWires[1117] ;
wire \normalizedWires[1116] ;
wire \normalizedWires[1115] ;
wire \normalizedWires[1114] ;
wire \normalizedWires[1113] ;
wire \normalizedWires[1112] ;
wire \normalizedWires[1111] ;
wire \normalizedWires[1110] ;
wire \normalizedWires[1109] ;
wire \normalizedWires[1108] ;
wire \normalizedWires[1107] ;
wire \normalizedWires[1106] ;
wire \normalizedWires[1105] ;
wire \normalizedWires[1070] ;
wire \normalizedWires[1069] ;
wire \normalizedWires[1068] ;
wire \normalizedWires[1067] ;
wire \normalizedWires[1066] ;
wire \normalizedWires[1065] ;
wire \normalizedWires[1064] ;
wire \normalizedWires[1063] ;
wire \normalizedWires[1062] ;
wire \normalizedWires[1061] ;
wire \normalizedWires[1060] ;
wire \normalizedWires[1059] ;
wire \normalizedWires[1058] ;
wire \normalizedWires[1057] ;
wire \normalizedWires[1056] ;
wire \normalizedWires[1055] ;
wire \normalizedWires[1054] ;
wire \normalizedWires[1053] ;
wire \normalizedWires[1052] ;
wire \normalizedWires[1051] ;
wire \normalizedWires[1050] ;
wire \normalizedWires[1049] ;
wire \normalizedWires[1048] ;
wire \normalizedWires[1047] ;
wire \normalizedWires[1046] ;
wire \normalizedWires[1045] ;
wire \normalizedWires[1044] ;
wire \normalizedWires[1043] ;
wire \normalizedWires[1042] ;
wire \normalizedWires[1041] ;
wire \normalizedWires[1040] ;
wire \normalizedWires[1005] ;
wire \normalizedWires[1004] ;
wire \normalizedWires[1003] ;
wire \normalizedWires[1002] ;
wire \normalizedWires[1001] ;
wire \normalizedWires[1000] ;
wire \normalizedWires[999] ;
wire \normalizedWires[998] ;
wire \normalizedWires[997] ;
wire \normalizedWires[996] ;
wire \normalizedWires[995] ;
wire \normalizedWires[994] ;
wire \normalizedWires[993] ;
wire \normalizedWires[992] ;
wire \normalizedWires[991] ;
wire \normalizedWires[990] ;
wire \normalizedWires[989] ;
wire \normalizedWires[988] ;
wire \normalizedWires[987] ;
wire \normalizedWires[986] ;
wire \normalizedWires[985] ;
wire \normalizedWires[984] ;
wire \normalizedWires[983] ;
wire \normalizedWires[982] ;
wire \normalizedWires[981] ;
wire \normalizedWires[980] ;
wire \normalizedWires[979] ;
wire \normalizedWires[978] ;
wire \normalizedWires[977] ;
wire \normalizedWires[976] ;
wire \normalizedWires[975] ;
wire \normalizedWires[940] ;
wire \normalizedWires[939] ;
wire \normalizedWires[938] ;
wire \normalizedWires[937] ;
wire \normalizedWires[936] ;
wire \normalizedWires[935] ;
wire \normalizedWires[934] ;
wire \normalizedWires[933] ;
wire \normalizedWires[932] ;
wire \normalizedWires[931] ;
wire \normalizedWires[930] ;
wire \normalizedWires[929] ;
wire \normalizedWires[928] ;
wire \normalizedWires[927] ;
wire \normalizedWires[926] ;
wire \normalizedWires[925] ;
wire \normalizedWires[924] ;
wire \normalizedWires[923] ;
wire \normalizedWires[922] ;
wire \normalizedWires[921] ;
wire \normalizedWires[920] ;
wire \normalizedWires[919] ;
wire \normalizedWires[918] ;
wire \normalizedWires[917] ;
wire \normalizedWires[916] ;
wire \normalizedWires[915] ;
wire \normalizedWires[914] ;
wire \normalizedWires[913] ;
wire \normalizedWires[912] ;
wire \normalizedWires[911] ;
wire \normalizedWires[910] ;
wire \normalizedWires[875] ;
wire \normalizedWires[874] ;
wire \normalizedWires[873] ;
wire \normalizedWires[872] ;
wire \normalizedWires[871] ;
wire \normalizedWires[870] ;
wire \normalizedWires[869] ;
wire \normalizedWires[868] ;
wire \normalizedWires[867] ;
wire \normalizedWires[866] ;
wire \normalizedWires[865] ;
wire \normalizedWires[864] ;
wire \normalizedWires[863] ;
wire \normalizedWires[862] ;
wire \normalizedWires[861] ;
wire \normalizedWires[860] ;
wire \normalizedWires[859] ;
wire \normalizedWires[858] ;
wire \normalizedWires[857] ;
wire \normalizedWires[856] ;
wire \normalizedWires[855] ;
wire \normalizedWires[854] ;
wire \normalizedWires[853] ;
wire \normalizedWires[852] ;
wire \normalizedWires[851] ;
wire \normalizedWires[850] ;
wire \normalizedWires[849] ;
wire \normalizedWires[848] ;
wire \normalizedWires[847] ;
wire \normalizedWires[846] ;
wire \normalizedWires[845] ;
wire \normalizedWires[810] ;
wire \normalizedWires[809] ;
wire \normalizedWires[808] ;
wire \normalizedWires[807] ;
wire \normalizedWires[806] ;
wire \normalizedWires[805] ;
wire \normalizedWires[804] ;
wire \normalizedWires[803] ;
wire \normalizedWires[802] ;
wire \normalizedWires[801] ;
wire \normalizedWires[800] ;
wire \normalizedWires[799] ;
wire \normalizedWires[798] ;
wire \normalizedWires[797] ;
wire \normalizedWires[796] ;
wire \normalizedWires[795] ;
wire \normalizedWires[794] ;
wire \normalizedWires[793] ;
wire \normalizedWires[792] ;
wire \normalizedWires[791] ;
wire \normalizedWires[790] ;
wire \normalizedWires[789] ;
wire \normalizedWires[788] ;
wire \normalizedWires[787] ;
wire \normalizedWires[786] ;
wire \normalizedWires[785] ;
wire \normalizedWires[784] ;
wire \normalizedWires[783] ;
wire \normalizedWires[782] ;
wire \normalizedWires[781] ;
wire \normalizedWires[780] ;
wire \normalizedWires[745] ;
wire \normalizedWires[744] ;
wire \normalizedWires[743] ;
wire \normalizedWires[742] ;
wire \normalizedWires[741] ;
wire \normalizedWires[740] ;
wire \normalizedWires[739] ;
wire \normalizedWires[738] ;
wire \normalizedWires[737] ;
wire \normalizedWires[736] ;
wire \normalizedWires[735] ;
wire \normalizedWires[734] ;
wire \normalizedWires[733] ;
wire \normalizedWires[732] ;
wire \normalizedWires[731] ;
wire \normalizedWires[730] ;
wire \normalizedWires[729] ;
wire \normalizedWires[728] ;
wire \normalizedWires[727] ;
wire \normalizedWires[726] ;
wire \normalizedWires[725] ;
wire \normalizedWires[724] ;
wire \normalizedWires[723] ;
wire \normalizedWires[722] ;
wire \normalizedWires[721] ;
wire \normalizedWires[720] ;
wire \normalizedWires[719] ;
wire \normalizedWires[718] ;
wire \normalizedWires[717] ;
wire \normalizedWires[716] ;
wire \normalizedWires[715] ;
wire \normalizedWires[680] ;
wire \normalizedWires[679] ;
wire \normalizedWires[678] ;
wire \normalizedWires[677] ;
wire \normalizedWires[676] ;
wire \normalizedWires[675] ;
wire \normalizedWires[674] ;
wire \normalizedWires[673] ;
wire \normalizedWires[672] ;
wire \normalizedWires[671] ;
wire \normalizedWires[670] ;
wire \normalizedWires[669] ;
wire \normalizedWires[668] ;
wire \normalizedWires[667] ;
wire \normalizedWires[666] ;
wire \normalizedWires[665] ;
wire \normalizedWires[664] ;
wire \normalizedWires[663] ;
wire \normalizedWires[662] ;
wire \normalizedWires[661] ;
wire \normalizedWires[660] ;
wire \normalizedWires[659] ;
wire \normalizedWires[658] ;
wire \normalizedWires[657] ;
wire \normalizedWires[656] ;
wire \normalizedWires[655] ;
wire \normalizedWires[654] ;
wire \normalizedWires[653] ;
wire \normalizedWires[652] ;
wire \normalizedWires[651] ;
wire \normalizedWires[650] ;
wire \normalizedWires[615] ;
wire \normalizedWires[614] ;
wire \normalizedWires[613] ;
wire \normalizedWires[612] ;
wire \normalizedWires[611] ;
wire \normalizedWires[610] ;
wire \normalizedWires[609] ;
wire \normalizedWires[608] ;
wire \normalizedWires[607] ;
wire \normalizedWires[606] ;
wire \normalizedWires[605] ;
wire \normalizedWires[604] ;
wire \normalizedWires[603] ;
wire \normalizedWires[602] ;
wire \normalizedWires[601] ;
wire \normalizedWires[600] ;
wire \normalizedWires[599] ;
wire \normalizedWires[598] ;
wire \normalizedWires[597] ;
wire \normalizedWires[596] ;
wire \normalizedWires[595] ;
wire \normalizedWires[594] ;
wire \normalizedWires[593] ;
wire \normalizedWires[592] ;
wire \normalizedWires[591] ;
wire \normalizedWires[590] ;
wire \normalizedWires[589] ;
wire \normalizedWires[588] ;
wire \normalizedWires[587] ;
wire \normalizedWires[586] ;
wire \normalizedWires[585] ;
wire \normalizedWires[550] ;
wire \normalizedWires[549] ;
wire \normalizedWires[548] ;
wire \normalizedWires[547] ;
wire \normalizedWires[546] ;
wire \normalizedWires[545] ;
wire \normalizedWires[544] ;
wire \normalizedWires[543] ;
wire \normalizedWires[542] ;
wire \normalizedWires[541] ;
wire \normalizedWires[540] ;
wire \normalizedWires[539] ;
wire \normalizedWires[538] ;
wire \normalizedWires[537] ;
wire \normalizedWires[536] ;
wire \normalizedWires[535] ;
wire \normalizedWires[534] ;
wire \normalizedWires[533] ;
wire \normalizedWires[532] ;
wire \normalizedWires[531] ;
wire \normalizedWires[530] ;
wire \normalizedWires[529] ;
wire \normalizedWires[528] ;
wire \normalizedWires[527] ;
wire \normalizedWires[526] ;
wire \normalizedWires[525] ;
wire \normalizedWires[524] ;
wire \normalizedWires[523] ;
wire \normalizedWires[522] ;
wire \normalizedWires[521] ;
wire \normalizedWires[520] ;
wire \normalizedWires[485] ;
wire \normalizedWires[484] ;
wire \normalizedWires[483] ;
wire \normalizedWires[482] ;
wire \normalizedWires[481] ;
wire \normalizedWires[480] ;
wire \normalizedWires[479] ;
wire \normalizedWires[478] ;
wire \normalizedWires[477] ;
wire \normalizedWires[476] ;
wire \normalizedWires[475] ;
wire \normalizedWires[474] ;
wire \normalizedWires[473] ;
wire \normalizedWires[472] ;
wire \normalizedWires[471] ;
wire \normalizedWires[470] ;
wire \normalizedWires[469] ;
wire \normalizedWires[468] ;
wire \normalizedWires[467] ;
wire \normalizedWires[466] ;
wire \normalizedWires[465] ;
wire \normalizedWires[464] ;
wire \normalizedWires[463] ;
wire \normalizedWires[462] ;
wire \normalizedWires[461] ;
wire \normalizedWires[460] ;
wire \normalizedWires[459] ;
wire \normalizedWires[458] ;
wire \normalizedWires[457] ;
wire \normalizedWires[456] ;
wire \normalizedWires[455] ;
wire \normalizedWires[420] ;
wire \normalizedWires[419] ;
wire \normalizedWires[418] ;
wire \normalizedWires[417] ;
wire \normalizedWires[416] ;
wire \normalizedWires[415] ;
wire \normalizedWires[414] ;
wire \normalizedWires[413] ;
wire \normalizedWires[412] ;
wire \normalizedWires[411] ;
wire \normalizedWires[410] ;
wire \normalizedWires[409] ;
wire \normalizedWires[408] ;
wire \normalizedWires[407] ;
wire \normalizedWires[406] ;
wire \normalizedWires[405] ;
wire \normalizedWires[404] ;
wire \normalizedWires[403] ;
wire \normalizedWires[402] ;
wire \normalizedWires[401] ;
wire \normalizedWires[400] ;
wire \normalizedWires[399] ;
wire \normalizedWires[398] ;
wire \normalizedWires[397] ;
wire \normalizedWires[396] ;
wire \normalizedWires[395] ;
wire \normalizedWires[394] ;
wire \normalizedWires[393] ;
wire \normalizedWires[392] ;
wire \normalizedWires[391] ;
wire \normalizedWires[390] ;
wire \normalizedWires[355] ;
wire \normalizedWires[354] ;
wire \normalizedWires[353] ;
wire \normalizedWires[352] ;
wire \normalizedWires[351] ;
wire \normalizedWires[350] ;
wire \normalizedWires[349] ;
wire \normalizedWires[348] ;
wire \normalizedWires[347] ;
wire \normalizedWires[346] ;
wire \normalizedWires[345] ;
wire \normalizedWires[344] ;
wire \normalizedWires[343] ;
wire \normalizedWires[342] ;
wire \normalizedWires[341] ;
wire \normalizedWires[340] ;
wire \normalizedWires[339] ;
wire \normalizedWires[338] ;
wire \normalizedWires[337] ;
wire \normalizedWires[336] ;
wire \normalizedWires[335] ;
wire \normalizedWires[334] ;
wire \normalizedWires[333] ;
wire \normalizedWires[332] ;
wire \normalizedWires[331] ;
wire \normalizedWires[330] ;
wire \normalizedWires[329] ;
wire \normalizedWires[328] ;
wire \normalizedWires[327] ;
wire \normalizedWires[326] ;
wire \normalizedWires[325] ;
wire \normalizedWires[290] ;
wire \normalizedWires[289] ;
wire \normalizedWires[288] ;
wire \normalizedWires[287] ;
wire \normalizedWires[286] ;
wire \normalizedWires[285] ;
wire \normalizedWires[284] ;
wire \normalizedWires[283] ;
wire \normalizedWires[282] ;
wire \normalizedWires[281] ;
wire \normalizedWires[280] ;
wire \normalizedWires[279] ;
wire \normalizedWires[278] ;
wire \normalizedWires[277] ;
wire \normalizedWires[276] ;
wire \normalizedWires[275] ;
wire \normalizedWires[274] ;
wire \normalizedWires[273] ;
wire \normalizedWires[272] ;
wire \normalizedWires[271] ;
wire \normalizedWires[270] ;
wire \normalizedWires[269] ;
wire \normalizedWires[268] ;
wire \normalizedWires[267] ;
wire \normalizedWires[266] ;
wire \normalizedWires[265] ;
wire \normalizedWires[264] ;
wire \normalizedWires[263] ;
wire \normalizedWires[262] ;
wire \normalizedWires[261] ;
wire \normalizedWires[260] ;
wire sph__n4212;
wire sph__n4211;
wire CLOCK_slh__n3555;
wire CLOCK_slh__n3554;
wire CLOCK_slh__n3553;
wire CLOCK_slh__n3549;
wire CLOCK_slh__n3548;
wire CLOCK_slh__n3547;
wire CLOCK_slh__n3543;
wire CLOCK_slh__n3542;
wire CLOCK_slh__n3541;
wire CLOCK_slh__n3537;
wire CLOCK_slh__n3536;
wire CLOCK_slh__n3535;
wire CLOCK_slh__n3531;
wire CLOCK_slh__n3530;
wire CLOCK_slh__n3529;
wire CLOCK_slh__n3521;
wire CLOCK_slh__n3520;
wire CLOCK_slh__n3519;
wire CLOCK_slh__n3511;
wire opt_ipo_n1428;
wire CLOCK_slh__n3510;
wire CLOCK_slh__n3509;
wire CLOCK_slo__mro_n3162;
wire CLOCK_slh__n3501;
wire CLOCK_slh__n3500;
wire CLOCK_slh__n3499;
wire opt_ipo_n1598;
wire CLOCK_slo__sro_n3372;
wire CLOCK_slo__sro_n3371;
wire CLOCK_slo__n3265;
wire CLOCK_slo__sro_n2844;
wire CLOCK_slo__sro_n2843;
wire \normalizedWires[225] ;
wire \normalizedWires[224] ;
wire \normalizedWires[223] ;
wire \normalizedWires[222] ;
wire \normalizedWires[221] ;
wire \normalizedWires[220] ;
wire \normalizedWires[219] ;
wire \normalizedWires[218] ;
wire \normalizedWires[217] ;
wire \normalizedWires[216] ;
wire \normalizedWires[215] ;
wire \normalizedWires[214] ;
wire \normalizedWires[213] ;
wire \normalizedWires[212] ;
wire \normalizedWires[211] ;
wire \normalizedWires[210] ;
wire \normalizedWires[209] ;
wire \normalizedWires[208] ;
wire \normalizedWires[207] ;
wire \normalizedWires[206] ;
wire \normalizedWires[205] ;
wire \normalizedWires[204] ;
wire \normalizedWires[203] ;
wire \normalizedWires[202] ;
wire \normalizedWires[201] ;
wire \normalizedWires[200] ;
wire \normalizedWires[199] ;
wire \normalizedWires[198] ;
wire \normalizedWires[197] ;
wire \normalizedWires[196] ;
wire \normalizedWires[195] ;
wire CLOCK_slo__sro_n2842;
wire CLOCK_slo__sro_n2795;
wire CLOCK_slo__sro_n2794;
wire CLOCK_slo__sro_n2793;
wire CLOCK_slo__sro_n2685;
wire CLOCK_slo__sro_n2684;
wire opt_ipo_n1569;
wire CLOCK_slo__sro_n2662;
wire CLOCK_slo__n2626;
wire CLOCK_slo__sro_n2425;
wire CLOCK_slo___n2653;
wire CLOCK_slo__sro_n2424;
wire opt_ipo_n1555;
wire CLOCK_slo__n2449;
wire opt_ipo_n1365;
wire opt_ipo_n1364;
wire opt_ipo_n1363;
wire CLOCK_slo__sro_n2299;
wire opt_ipo_n1361;
wire opt_ipo_n1551;
wire opt_ipo_n1547;
wire CLOCK_slo__sro_n3067;
wire CLOCK_sgo__sro_n1965;
wire opt_ipo_n1541;
wire opt_ipo_n1540;
wire CLOCK_slo__sro_n3066;
wire CLOCK_sgo__sro_n1964;
wire opt_ipo_n1344;
wire CLOCK_slo__sro_n3065;
wire CLOCK_slo__sro_n3068;
wire CLOCK_opt_ipo_n1683;
wire CLOCK_slo__sro_n2214;
wire CLOCK_slo__mro_n3163;
wire \normalizedWires[160] ;
wire \normalizedWires[159] ;
wire \normalizedWires[158] ;
wire \normalizedWires[157] ;
wire \normalizedWires[156] ;
wire \normalizedWires[155] ;
wire \normalizedWires[154] ;
wire \normalizedWires[153] ;
wire \normalizedWires[152] ;
wire \normalizedWires[151] ;
wire \normalizedWires[150] ;
wire \normalizedWires[149] ;
wire \normalizedWires[148] ;
wire \normalizedWires[147] ;
wire \normalizedWires[146] ;
wire \normalizedWires[145] ;
wire \normalizedWires[144] ;
wire \normalizedWires[143] ;
wire \normalizedWires[142] ;
wire \normalizedWires[141] ;
wire \normalizedWires[140] ;
wire \normalizedWires[139] ;
wire \normalizedWires[138] ;
wire \normalizedWires[137] ;
wire \normalizedWires[136] ;
wire \normalizedWires[135] ;
wire \normalizedWires[134] ;
wire \normalizedWires[133] ;
wire \normalizedWires[132] ;
wire \normalizedWires[131] ;
wire \normalizedWires[130] ;
wire slo__sro_n1189;
wire slo__sro_n1188;
wire slo__sro_n1187;
wire slo__sro_n1153;
wire slo__sro_n1152;
wire slo__sro_n1151;
wire slo__sro_n1133;
wire slo__sro_n1132;
wire slo__sro_n1131;
wire slo__sro_n1123;
wire slo__sro_n1122;
wire slo__sro_n1121;
wire slo__sro_n1082;
wire slo__sro_n1081;
wire slo__sro_n1080;
wire slo__sro_n1027;
wire slo__sro_n1026;
wire slo__sro_n1029;
wire slo__sro_n1028;
wire slo__sro_n1001;
wire slo__n980;
wire slo__n798;
wire slo__sro_n1000;
wire slo__n881;
wire slo__sro_n999;
wire slo__sro_n905;
wire CLOCK_slo__n2403;
wire slo__sro_n703;
wire slo__sro_n702;
wire slo__sro_n701;
wire slo__sro_n670;
wire slo__sro_n669;
wire slo__sro_n668;
wire slo__n619;
wire \normalizedWires[95] ;
wire \normalizedWires[94] ;
wire \normalizedWires[93] ;
wire \normalizedWires[92] ;
wire \normalizedWires[91] ;
wire \normalizedWires[90] ;
wire \normalizedWires[89] ;
wire \normalizedWires[88] ;
wire \normalizedWires[87] ;
wire \normalizedWires[86] ;
wire \normalizedWires[85] ;
wire \normalizedWires[84] ;
wire \normalizedWires[83] ;
wire \normalizedWires[82] ;
wire \normalizedWires[81] ;
wire \normalizedWires[80] ;
wire \normalizedWires[79] ;
wire \normalizedWires[78] ;
wire \normalizedWires[77] ;
wire \normalizedWires[76] ;
wire \normalizedWires[75] ;
wire \normalizedWires[74] ;
wire \normalizedWires[73] ;
wire \normalizedWires[72] ;
wire \normalizedWires[71] ;
wire \normalizedWires[70] ;
wire \normalizedWires[69] ;
wire \normalizedWires[68] ;
wire \normalizedWires[67] ;
wire \normalizedWires[66] ;
wire \normalizedWires[65] ;
wire slo__sro_n561;
wire slo__sro_n560;
wire slo__sro_n559;
wire slo__sro_n551;
wire CLOCK_slo__sro_n3369;
wire slo__sro_n549;
wire slo__sro_n541;
wire slo__sro_n540;
wire slo__sro_n539;
wire slo__sro_n538;
wire slo__mro_n474;
wire slo__sro_n516;
wire slo__sro_n515;
wire slo__sro_n514;
wire CLOCK_slo__sro_n2682;
wire slo__n453;
wire slo__sro_n423;
wire slo__sro_n422;
wire slo__sro_n421;
wire slo__sro_n408;
wire slo__mro_n394;
wire slo__mro_n393;
wire slo__mro_n392;
wire slo__sro_n384;
wire slo__sro_n383;
wire slo__sro_n382;
wire slo__sro_n381;
wire slo__sro_n366;
wire slo__sro_n365;
wire slo__sro_n364;
wire slo__xsl_n298;
wire sgo__sro_n130;
wire sgo__sro_n246;
wire sgo__sro_n145;
wire \normalizedWires[30] ;
wire \normalizedWires[29] ;
wire \normalizedWires[28] ;
wire \normalizedWires[27] ;
wire \normalizedWires[26] ;
wire \normalizedWires[25] ;
wire \normalizedWires[24] ;
wire \normalizedWires[23] ;
wire \normalizedWires[22] ;
wire \normalizedWires[21] ;
wire \normalizedWires[20] ;
wire \normalizedWires[19] ;
wire \normalizedWires[18] ;
wire \normalizedWires[17] ;
wire \normalizedWires[16] ;
wire \normalizedWires[15] ;
wire \normalizedWires[14] ;
wire \normalizedWires[13] ;
wire \normalizedWires[12] ;
wire \normalizedWires[11] ;
wire \normalizedWires[10] ;
wire \normalizedWires[9] ;
wire \normalizedWires[8] ;
wire \normalizedWires[7] ;
wire \normalizedWires[6] ;
wire \normalizedWires[5] ;
wire \normalizedWires[4] ;
wire \normalizedWires[3] ;
wire \normalizedWires[2] ;
wire \normalizedWires[1] ;
wire sgo__sro_n146;
wire \Res_imm[63] ;
wire \Res_imm[62] ;
wire \Res_imm[61] ;
wire \Res_imm[60] ;
wire \Res_imm[59] ;
wire \Res_imm[58] ;
wire \Res_imm[57] ;
wire \Res_imm[56] ;
wire \Res_imm[55] ;
wire \Res_imm[54] ;
wire \Res_imm[53] ;
wire \Res_imm[52] ;
wire \Res_imm[51] ;
wire \Res_imm[50] ;
wire \Res_imm[49] ;
wire \Res_imm[48] ;
wire \Res_imm[47] ;
wire \Res_imm[46] ;
wire \Res_imm[45] ;
wire \Res_imm[44] ;
wire \Res_imm[43] ;
wire \Res_imm[42] ;
wire \Res_imm[41] ;
wire \Res_imm[40] ;
wire \Res_imm[39] ;
wire \Res_imm[38] ;
wire \Res_imm[37] ;
wire \Res_imm[36] ;
wire \Res_imm[35] ;
wire \Res_imm[34] ;
wire \Res_imm[33] ;
wire \Res_imm[32] ;
wire \Res_imm[31] ;
wire \Res_imm[30] ;
wire \Res_imm[29] ;
wire \Res_imm[28] ;
wire \Res_imm[27] ;
wire \Res_imm[26] ;
wire \Res_imm[25] ;
wire \Res_imm[24] ;
wire \Res_imm[23] ;
wire \Res_imm[22] ;
wire \Res_imm[21] ;
wire \Res_imm[20] ;
wire \Res_imm[19] ;
wire \Res_imm[18] ;
wire \Res_imm[17] ;
wire \Res_imm[16] ;
wire \Res_imm[15] ;
wire \Res_imm[14] ;
wire \Res_imm[13] ;
wire \Res_imm[12] ;
wire \Res_imm[11] ;
wire \Res_imm[10] ;
wire \Res_imm[9] ;
wire sgo__sro_n53;
wire slo__sro_n407;
wire drc_ipo_n27;
wire sgo__n28;
wire sgo__sro_n51;
wire CLOCK_slo__mro_n2292;
wire drc_ipo_n26;
wire hfn_ipo_n25;
wire sgo__sro_n34;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire B_in;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire A_in;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_256;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_169;
wire n_0_170;
wire n_0_171;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_176;
wire n_0_177;
wire n_0_178;
wire n_0_179;
wire n_0_180;
wire n_0_181;
wire n_0_182;
wire n_0_183;
wire n_0_184;
wire n_0_249;
wire n_0_250;
wire n_0_251;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_255;
wire n_0_257;
wire n_0_258;
wire n_0_259;
wire n_0_260;
wire n_0_261;
wire n_0_262;
wire n_0_263;
wire n_0_264;
wire n_0_265;
wire n_0_266;
wire n_0_267;
wire n_0_268;
wire n_0_269;
wire n_0_270;
wire n_0_271;
wire n_0_272;
wire n_0_273;
wire n_0_274;
wire n_0_275;
wire n_0_276;
wire n_0_277;
wire n_0_278;
wire n_0_279;
wire n_0_280;
wire n_0_281;
wire n_0_283;
wire n_0_284;
wire n_0_285;
wire n_0_286;
wire n_0_287;
wire n_0_288;
wire n_0_289;
wire n_0_290;
wire n_0_291;
wire n_0_292;
wire n_0_293;
wire n_0_294;
wire n_0_295;
wire n_0_296;
wire n_0_297;
wire n_0_298;
wire n_0_299;
wire n_0_300;
wire n_0_301;
wire n_0_302;
wire n_0_303;
wire n_0_304;
wire n_0_305;
wire n_0_306;
wire n_0_307;
wire n_0_308;
wire n_0_309;
wire n_0_310;
wire n_0_311;
wire n_0_312;
wire n_0_313;
wire n_0_314;
wire \B_imm[31] ;
wire \B_imm[30] ;
wire \B_imm[29] ;
wire \B_imm[28] ;
wire \B_imm[27] ;
wire \B_imm[26] ;
wire CLOCK_slo__sro_n2301;
wire CLOCK_slo__sro_n2841;
wire \B_imm[23] ;
wire slo__sro_n534;
wire slo__sro_n1186;
wire \B_imm[20] ;
wire \B_imm[19] ;
wire \B_imm[18] ;
wire \B_imm[17] ;
wire CLOCK_slo__n2760;
wire CLOCK_slo__sro_n2796;
wire \B_imm[14] ;
wire \B_imm[13] ;
wire \B_imm[12] ;
wire \B_imm[11] ;
wire slo__sro_n513;
wire CLOCK_sgo__sro_n1959;
wire \B_imm[8] ;
wire CLOCK_slo__sro_n2298;
wire CLOCK_slo__mro_n3164;
wire \B_imm[5] ;
wire \B_imm[4] ;
wire \B_imm[3] ;
wire \B_imm[2] ;
wire \B_imm[1] ;
wire CLOCK_slo__sro_n2213;
wire \A_imm[30] ;
wire \A_imm[29] ;
wire \A_imm[28] ;
wire \A_imm[27] ;
wire slo__sro_n558;
wire slo__sro_n420;
wire CLOCK_slo___n3239;
wire \A_imm[22] ;
wire slo__sro_n700;
wire slo__n378;
wire slo__mro_n391;
wire CLOCK_slo__sro_n3370;
wire slo__sro_n1150;
wire slo__sro_n1120;
wire slo__sro_n1079;
wire CTS_n_tid0_1747;
wire CLOCK_slo__sro_n2300;
wire \A_imm[12] ;
wire \A_imm[11] ;
wire slo__sro_n667;
wire \A_imm[9] ;
wire \A_imm[8] ;
wire \A_imm[7] ;
wire \A_imm[6] ;
wire \A_imm[5] ;
wire \A_imm[4] ;
wire \A_imm[3] ;
wire \A_imm[2] ;
wire \A_imm[1] ;
wire n_0_185;
wire n_0_1_29;
wire n_0_1_30;
wire n_0_186;
wire n_0_1_31;
wire n_0_1_32;
wire n_0_187;
wire n_0_1_33;
wire n_0_1_34;
wire n_0_188;
wire n_0_1_35;
wire n_0_1_36;
wire n_0_189;
wire n_0_1_37;
wire n_0_1_38;
wire n_0_190;
wire n_0_1_39;
wire n_0_1_40;
wire n_0_191;
wire n_0_1_41;
wire n_0_1_42;
wire n_0_192;
wire n_0_1_43;
wire n_0_1_44;
wire n_0_193;
wire n_0_1_45;
wire n_0_1_46;
wire n_0_194;
wire n_0_1_47;
wire n_0_1_48;
wire n_0_195;
wire n_0_1_49;
wire n_0_1_50;
wire n_0_196;
wire n_0_1_51;
wire n_0_1_52;
wire n_0_197;
wire n_0_1_53;
wire n_0_1_54;
wire n_0_198;
wire n_0_1_55;
wire n_0_1_56;
wire n_0_199;
wire n_0_1_57;
wire n_0_1_58;
wire n_0_200;
wire n_0_1_59;
wire n_0_1_60;
wire n_0_201;
wire n_0_1_61;
wire n_0_1_62;
wire n_0_202;
wire n_0_1_63;
wire n_0_1_64;
wire n_0_203;
wire n_0_1_65;
wire n_0_1_66;
wire n_0_204;
wire n_0_1_67;
wire n_0_1_72;
wire n_0_205;
wire n_0_1_77;
wire n_0_1_78;
wire n_0_206;
wire n_0_1_79;
wire n_0_1_80;
wire n_0_207;
wire n_0_1_81;
wire n_0_1_82;
wire n_0_208;
wire n_0_1_83;
wire n_0_1_84;
wire n_0_209;
wire n_0_1_85;
wire n_0_1_86;
wire n_0_210;
wire n_0_1_87;
wire n_0_1_88;
wire n_0_211;
wire n_0_1_91;
wire n_0_1_92;
wire n_0_212;
wire n_0_1_93;
wire n_0_1_94;
wire n_0_213;
wire n_0_1_95;
wire n_0_1_96;
wire n_0_214;
wire n_0_1_97;
wire n_0_1_98;
wire n_0_215;
wire n_0_1_99;
wire n_0_1_100;
wire n_0_216;
wire n_0_1_101;
wire n_0_1_102;
wire n_0_217;
wire n_0_1_103;
wire n_0_1_104;
wire n_0_218;
wire n_0_1_105;
wire n_0_1_106;
wire n_0_219;
wire n_0_1_107;
wire n_0_1_108;
wire n_0_220;
wire n_0_1_109;
wire n_0_1_110;
wire n_0_221;
wire n_0_1_111;
wire n_0_1_112;
wire n_0_223;
wire n_0_1_113;
wire n_0_1_114;
wire n_0_224;
wire n_0_1_115;
wire n_0_1_116;
wire n_0_226;
wire n_0_1_117;
wire n_0_1_118;
wire n_0_227;
wire n_0_1_119;
wire n_0_1_120;
wire n_0_228;
wire n_0_1_121;
wire n_0_1_122;
wire n_0_229;
wire n_0_1_123;
wire n_0_1_124;
wire n_0_230;
wire n_0_1_125;
wire n_0_1_126;
wire n_0_231;
wire n_0_1_127;
wire n_0_1_128;
wire n_0_232;
wire n_0_1_129;
wire n_0_1_130;
wire n_0_233;
wire n_0_1_131;
wire n_0_1_132;
wire n_0_237;
wire n_0_1_133;
wire n_0_1_134;
wire n_0_243;
wire n_0_1_135;
wire n_0_1_136;
wire CLOCK_opt_ipo_n1670;
wire n_0_222;
wire n_0_1_138;
wire n_0_1_139;
wire n_0_234;
wire n_0_1_140;
wire n_0_1_141;
wire n_0_238;
wire n_0_1_146;
wire n_0_1_147;
wire n_0_239;
wire n_0_1_148;
wire n_0_1_149;
wire n_0_241;
wire n_0_1_152;
wire n_0_1_153;
wire sgo__sro_n35;
wire CLOCK_slo__mro_n2310;
wire n_0_246;
wire n_0_1_0;
wire n_0_1_1;
wire n_0_248;
wire n_0_1_2;
wire n_0_244;
wire n_0_1_3;
wire n_0_1_4;
wire n_0_1_24;
wire opt_ipo_n1652;
wire hfn_ipo_n23;
wire n_0_1_5;
wire n_0_1_6;
wire n_0_235;
wire n_0_1_7;
wire n_0_236;
wire n_0_1_8;
wire n_0_242;
wire n_0_1_9;
wire CLOCK_slo__sro_n2663;
wire n_0_1_10;
wire n_0_247;
wire CTS_n1731;
wire CTS_n1730;
wire n_0_315;
wire CLOCK_sgo__sro_n1963;
wire n_0_1_13;
wire hfn_ipo_n24;
wire slo__sro_n363;
wire hfn_ipo_n22;
wire CLOCK_slo__sro_n2215;
wire n_0_1_17;
wire slo__n345;
wire n_0_1_19;
wire n_0_1_20;
wire n_0_1_21;
wire n_0_1_22;
wire n_0_1_23;
wire slo__sro_n405;
wire n_0_1_26;
wire slo__sro_n406;
wire n_0_1_28;
wire n_0_1_68;
wire n_0_1_69;
wire n_0_1_70;
wire n_0_1_71;
wire n_0_1_73;
wire n_0_1_74;
wire n_0_1_75;
wire n_0_1_76;
wire n_0_1_142;
wire n_0_1_143;
wire n_0_1_144;
wire slo__sro_n535;
wire opt_ipo_n1524;
wire CLOCK_slo__sro_n2683;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire uc_28;
wire uc_29;
wire uc_30;
wire uc_31;
wire uc_32;
wire uc_33;
wire uc_34;
wire uc_35;
wire uc_36;
wire uc_37;
wire uc_38;
wire uc_39;
wire uc_40;
wire uc_41;
wire uc_42;
wire uc_43;
wire uc_44;
wire uc_45;
wire uc_46;
wire uc_47;
wire uc_48;
wire uc_49;
wire uc_50;
wire uc_51;
wire uc_52;
wire uc_53;
wire uc_54;
wire uc_55;
wire uc_56;
wire uc_57;
wire uc_58;
wire uc_59;
wire uc_60;
wire uc_61;
wire uc_62;
wire uc_63;
wire uc_64;
wire uc_65;
wire uc_66;
wire uc_67;
wire uc_68;
wire uc_69;
wire uc_70;
wire uc_71;
wire uc_72;
wire uc_73;
wire uc_74;
wire uc_75;
wire uc_76;
wire uc_77;
wire uc_78;
wire uc_79;
wire uc_80;
wire uc_81;
wire uc_82;
wire uc_83;
wire uc_84;
wire uc_85;
wire uc_86;
wire uc_87;
wire uc_88;
wire uc_89;
wire uc_90;
wire uc_91;
wire uc_92;
wire uc_93;
wire uc_94;
wire uc_95;
wire uc_96;
wire uc_97;
wire uc_98;
wire uc_99;
wire uc_100;
wire uc_101;
wire uc_102;
wire uc_103;
wire uc_104;
wire uc_105;
wire uc_106;
wire uc_107;
wire uc_108;
wire uc_109;
wire uc_110;
wire uc_111;
wire uc_112;
wire uc_113;
wire uc_114;
wire uc_115;
wire uc_116;
wire uc_117;
wire uc_118;
wire uc_119;
wire uc_120;
wire uc_121;
wire uc_122;
wire uc_123;
wire uc_124;
wire uc_125;
wire uc_126;
wire uc_127;
wire uc_128;
wire uc_129;
wire uc_130;
wire uc_131;
wire uc_132;
wire uc_133;
wire uc_134;
wire uc_135;
wire uc_136;
wire uc_137;
wire uc_138;
wire uc_139;
wire uc_140;
wire uc_141;
wire uc_142;
wire uc_143;
wire uc_144;
wire uc_145;
wire uc_146;
wire uc_147;
wire uc_148;
wire uc_149;
wire uc_150;
wire uc_151;
wire uc_152;
wire uc_153;
wire uc_154;
wire uc_155;
wire uc_156;
wire uc_157;
wire uc_158;
wire uc_159;
wire uc_160;
wire uc_161;
wire uc_162;
wire uc_163;
wire uc_164;
wire uc_165;
wire uc_166;
wire uc_167;
wire uc_168;
wire uc_169;
wire uc_170;
wire uc_171;
wire uc_172;
wire uc_173;
wire uc_174;
wire uc_175;
wire uc_176;
wire uc_177;
wire uc_178;
wire uc_179;
wire uc_180;
wire uc_181;
wire uc_182;
wire uc_183;
wire uc_184;
wire uc_185;
wire uc_186;
wire uc_187;
wire uc_188;
wire uc_189;
wire uc_190;
wire uc_191;
wire uc_192;
wire uc_193;
wire uc_194;
wire uc_195;
wire uc_196;
wire uc_197;
wire uc_198;
wire uc_199;
wire uc_200;
wire uc_201;
wire uc_202;
wire uc_203;
wire uc_204;
wire uc_205;
wire uc_206;
wire uc_207;
wire uc_208;
wire uc_209;
wire uc_210;
wire uc_211;
wire uc_212;
wire uc_213;
wire uc_214;
wire uc_215;
wire uc_216;
wire uc_217;
wire uc_218;
wire uc_219;
wire uc_220;
wire uc_221;
wire uc_222;
wire uc_223;
wire uc_224;
wire uc_225;
wire uc_226;
wire uc_227;
wire uc_228;
wire uc_229;
wire uc_230;
wire uc_231;
wire uc_232;
wire uc_233;
wire uc_234;
wire uc_235;
wire uc_236;
wire uc_237;
wire uc_238;
wire uc_239;
wire uc_240;
wire uc_241;
wire uc_242;
wire uc_243;
wire uc_244;
wire uc_245;
wire uc_246;
wire uc_247;
wire uc_248;
wire uc_249;
wire uc_250;
wire uc_251;
wire uc_252;
wire uc_253;
wire uc_254;
wire uc_255;
wire uc_256;
wire uc_257;
wire uc_258;
wire uc_259;
wire uc_260;
wire uc_261;
wire uc_262;
wire uc_263;
wire uc_264;
wire uc_265;
wire uc_266;
wire uc_267;
wire uc_268;
wire uc_269;
wire uc_270;
wire uc_271;
wire uc_272;
wire uc_273;
wire uc_274;
wire uc_275;
wire uc_276;
wire uc_277;
wire uc_278;
wire uc_279;
wire uc_280;
wire uc_281;
wire uc_282;
wire uc_283;
wire uc_284;
wire uc_285;
wire uc_286;
wire uc_287;
wire uc_288;
wire uc_289;
wire uc_290;
wire uc_291;
wire uc_292;
wire uc_293;
wire uc_294;
wire uc_295;
wire uc_296;
wire uc_297;
wire uc_298;
wire uc_299;
wire uc_300;
wire uc_301;
wire uc_302;
wire uc_303;
wire uc_304;
wire uc_305;
wire uc_306;
wire uc_307;
wire uc_308;
wire uc_309;
wire uc_310;
wire uc_311;
wire uc_312;
wire uc_313;
wire uc_314;
wire uc_315;
wire uc_316;
wire uc_317;
wire uc_318;
wire uc_319;
wire uc_320;
wire uc_321;
wire uc_322;
wire uc_323;
wire uc_324;
wire uc_325;
wire uc_326;
wire uc_327;
wire uc_328;
wire uc_329;
wire uc_330;
wire uc_331;
wire uc_332;
wire uc_333;
wire uc_334;
wire uc_335;
wire uc_336;
wire uc_337;
wire uc_338;
wire uc_339;
wire uc_340;
wire uc_341;
wire uc_342;
wire uc_343;
wire uc_344;
wire uc_345;
wire uc_346;
wire uc_347;
wire uc_348;
wire uc_349;
wire uc_350;
wire uc_351;
wire uc_352;
wire uc_353;
wire uc_354;
wire uc_355;
wire uc_356;
wire uc_357;
wire uc_358;
wire uc_359;
wire uc_360;
wire uc_361;
wire uc_362;
wire uc_363;
wire uc_364;
wire uc_365;
wire uc_366;
wire uc_367;
wire uc_368;
wire uc_369;
wire uc_370;
wire uc_371;
wire uc_372;
wire uc_373;
wire uc_374;
wire uc_375;
wire uc_376;
wire uc_377;
wire uc_378;
wire uc_379;
wire uc_380;
wire uc_381;
wire uc_382;
wire uc_383;
wire uc_384;
wire uc_385;
wire uc_386;
wire uc_387;
wire uc_388;
wire uc_389;
wire uc_390;
wire uc_391;
wire uc_392;
wire uc_393;
wire uc_394;
wire uc_395;
wire uc_396;
wire uc_397;
wire uc_398;
wire uc_399;
wire uc_400;
wire uc_401;
wire uc_402;
wire uc_403;
wire uc_404;
wire uc_405;
wire uc_406;
wire uc_407;
wire uc_408;
wire uc_409;
wire uc_410;
wire uc_411;
wire uc_412;
wire uc_413;
wire uc_414;
wire uc_415;
wire uc_416;
wire uc_417;
wire uc_418;
wire uc_419;
wire uc_420;
wire uc_421;
wire uc_422;
wire uc_423;
wire uc_424;
wire uc_425;
wire uc_426;
wire uc_427;
wire uc_428;
wire uc_429;
wire uc_430;
wire uc_431;
wire uc_432;
wire uc_433;
wire uc_434;
wire uc_435;
wire uc_436;
wire uc_437;
wire uc_438;
wire uc_439;
wire uc_440;
wire uc_441;
wire uc_442;
wire uc_443;
wire uc_444;
wire uc_445;
wire uc_446;
wire uc_447;
wire uc_448;
wire uc_449;
wire uc_450;
wire uc_451;
wire uc_452;
wire uc_453;
wire uc_454;
wire uc_455;
wire uc_456;
wire uc_457;
wire uc_458;
wire uc_459;
wire uc_460;
wire uc_461;
wire uc_462;
wire uc_463;
wire uc_464;
wire uc_465;
wire uc_466;
wire uc_467;
wire uc_468;
wire uc_469;
wire uc_470;
wire uc_471;
wire uc_472;
wire uc_473;
wire uc_474;
wire uc_475;
wire uc_476;
wire uc_477;
wire uc_478;
wire uc_479;
wire uc_480;
wire uc_481;
wire uc_482;
wire uc_483;
wire uc_484;
wire uc_485;
wire uc_486;
wire uc_487;
wire uc_488;
wire uc_489;
wire uc_490;
wire uc_491;
wire uc_492;
wire uc_493;
wire uc_494;
wire uc_495;
wire uc_496;
wire uc_497;
wire uc_498;
wire uc_499;
wire uc_500;
wire uc_501;
wire uc_502;
wire uc_503;
wire uc_504;
wire uc_505;
wire uc_506;
wire uc_507;
wire uc_508;
wire uc_509;
wire uc_510;
wire uc_511;
wire uc_512;
wire uc_513;
wire uc_514;
wire uc_515;
wire uc_516;
wire uc_517;
wire uc_518;
wire uc_519;
wire uc_520;
wire uc_521;
wire uc_522;
wire uc_523;
wire uc_524;
wire uc_525;
wire uc_526;
wire uc_527;
wire uc_528;
wire uc_529;
wire uc_530;
wire uc_531;
wire uc_532;
wire uc_533;
wire uc_534;
wire uc_535;
wire uc_536;
wire uc_537;
wire uc_538;
wire uc_539;
wire uc_540;
wire uc_541;
wire uc_542;
wire uc_543;
wire uc_544;
wire uc_545;
wire uc_546;
wire uc_547;
wire uc_548;
wire uc_549;
wire uc_550;
wire uc_551;
wire uc_552;
wire uc_553;
wire uc_554;
wire uc_555;
wire uc_556;
wire uc_557;
wire uc_558;
wire uc_559;
wire uc_560;
wire uc_561;
wire uc_562;
wire uc_563;
wire uc_564;
wire uc_565;
wire uc_566;
wire uc_567;
wire uc_568;
wire uc_569;
wire uc_570;
wire uc_571;
wire uc_572;
wire uc_573;
wire uc_574;
wire uc_575;
wire uc_576;
wire uc_577;
wire uc_578;
wire uc_579;
wire uc_580;
wire uc_581;
wire uc_582;
wire uc_583;
wire uc_584;
wire uc_585;
wire uc_586;
wire uc_587;
wire uc_588;
wire uc_589;
wire uc_590;
wire uc_591;
wire uc_592;
wire uc_593;
wire uc_594;
wire uc_595;
wire uc_596;
wire uc_597;
wire uc_598;
wire uc_599;
wire uc_600;
wire uc_601;
wire uc_602;
wire uc_603;
wire uc_604;
wire uc_605;
wire uc_606;
wire uc_607;
wire uc_608;
wire uc_609;
wire uc_610;
wire uc_611;
wire uc_612;
wire uc_613;
wire uc_614;
wire uc_615;
wire uc_616;
wire uc_617;
wire uc_618;
wire uc_619;
wire uc_620;
wire uc_621;
wire uc_622;
wire uc_623;
wire uc_624;
wire uc_625;
wire uc_626;
wire uc_627;
wire uc_628;
wire uc_629;
wire uc_630;
wire uc_631;
wire uc_632;
wire uc_633;
wire uc_634;
wire uc_635;
wire uc_636;
wire uc_637;
wire uc_638;
wire uc_639;
wire uc_640;
wire uc_641;
wire uc_642;
wire uc_643;
wire uc_644;
wire uc_645;
wire uc_646;
wire uc_647;
wire uc_648;
wire uc_649;
wire uc_650;
wire uc_651;
wire uc_652;
wire uc_653;
wire uc_654;
wire uc_655;
wire uc_656;
wire uc_657;
wire uc_658;
wire uc_659;
wire uc_660;
wire uc_661;
wire uc_662;
wire uc_663;
wire uc_664;
wire uc_665;
wire uc_666;
wire uc_667;
wire uc_668;
wire uc_669;
wire uc_670;
wire uc_671;
wire uc_672;
wire uc_673;
wire uc_674;
wire uc_675;
wire uc_676;
wire uc_677;
wire uc_678;
wire uc_679;
wire uc_680;
wire uc_681;
wire uc_682;
wire uc_683;
wire uc_684;
wire uc_685;
wire uc_686;
wire uc_687;
wire uc_688;
wire uc_689;
wire uc_690;
wire uc_691;
wire uc_692;
wire uc_693;
wire uc_694;
wire uc_695;
wire uc_696;
wire uc_697;
wire uc_698;
wire uc_699;
wire uc_700;
wire uc_701;
wire uc_702;
wire uc_703;
wire uc_704;
wire uc_705;
wire uc_706;
wire uc_707;
wire uc_708;
wire uc_709;
wire uc_710;
wire uc_711;
wire uc_712;
wire uc_713;
wire uc_714;
wire uc_715;
wire uc_716;
wire uc_717;
wire uc_718;
wire uc_719;
wire uc_720;
wire uc_721;
wire uc_722;
wire uc_723;
wire uc_724;
wire uc_725;
wire uc_726;
wire uc_727;
wire uc_728;
wire uc_729;
wire uc_730;
wire uc_731;
wire uc_732;
wire uc_733;
wire uc_734;
wire uc_735;
wire uc_736;
wire uc_737;
wire uc_738;
wire uc_739;
wire uc_740;
wire uc_741;
wire uc_742;
wire uc_743;
wire uc_744;
wire uc_745;
wire uc_746;
wire uc_747;
wire uc_748;
wire uc_749;
wire uc_750;
wire uc_751;
wire uc_752;
wire uc_753;
wire uc_754;
wire uc_755;
wire uc_756;
wire uc_757;
wire uc_758;
wire uc_759;
wire uc_760;
wire uc_761;
wire uc_762;
wire uc_763;
wire uc_764;
wire uc_765;
wire uc_766;
wire uc_767;
wire uc_768;
wire uc_769;
wire uc_770;
wire uc_771;
wire uc_772;
wire uc_773;
wire uc_774;
wire uc_775;
wire uc_776;
wire uc_777;
wire uc_778;
wire uc_779;
wire uc_780;
wire uc_781;
wire uc_782;
wire uc_783;
wire uc_784;
wire uc_785;
wire uc_786;
wire uc_787;
wire uc_788;
wire uc_789;
wire uc_790;
wire uc_791;
wire uc_792;
wire uc_793;
wire uc_794;
wire uc_795;
wire uc_796;
wire uc_797;
wire uc_798;
wire uc_799;
wire uc_800;
wire uc_801;
wire uc_802;
wire uc_803;
wire uc_804;
wire uc_805;
wire uc_806;
wire uc_807;
wire uc_808;
wire uc_809;
wire uc_810;
wire uc_811;
wire uc_812;
wire uc_813;
wire uc_814;
wire uc_815;
wire uc_816;
wire uc_817;
wire uc_818;
wire uc_819;
wire uc_820;
wire uc_821;
wire uc_822;
wire uc_823;
wire uc_824;
wire uc_825;
wire uc_826;
wire uc_827;
wire uc_828;
wire uc_829;
wire uc_830;
wire uc_831;
wire uc_832;
wire uc_833;
wire uc_834;
wire uc_835;
wire uc_836;
wire uc_837;
wire uc_838;
wire uc_839;
wire uc_840;
wire uc_841;
wire uc_842;
wire uc_843;
wire uc_844;
wire uc_845;
wire uc_846;
wire uc_847;
wire uc_848;
wire uc_849;
wire uc_850;
wire uc_851;
wire uc_852;
wire uc_853;
wire uc_854;
wire uc_855;
wire uc_856;
wire uc_857;
wire uc_858;
wire uc_859;
wire uc_860;
wire uc_861;
wire uc_862;
wire uc_863;
wire uc_864;
wire uc_865;
wire uc_866;
wire uc_867;
wire uc_868;
wire uc_869;
wire uc_870;
wire uc_871;
wire uc_872;
wire uc_873;
wire uc_874;
wire uc_875;
wire uc_876;
wire uc_877;
wire uc_878;
wire uc_879;
wire uc_880;
wire uc_881;
wire uc_882;
wire uc_883;
wire uc_884;
wire uc_885;
wire uc_886;
wire uc_887;
wire uc_888;
wire uc_889;
wire uc_890;
wire uc_891;
wire uc_892;
wire uc_893;
wire uc_894;
wire uc_895;
wire uc_896;
wire uc_897;
wire uc_898;
wire uc_899;
wire uc_900;
wire uc_901;
wire uc_902;
wire uc_903;
wire uc_904;
wire uc_905;
wire uc_906;
wire uc_907;
wire uc_908;
wire uc_909;
wire uc_910;
wire uc_911;
wire uc_912;
wire uc_913;
wire uc_914;
wire uc_915;
wire uc_916;
wire uc_917;
wire uc_918;
wire uc_919;
wire uc_920;
wire uc_921;
wire uc_922;
wire uc_923;
wire uc_924;
wire uc_925;
wire uc_926;
wire uc_927;
wire uc_928;
wire uc_929;
wire uc_930;
wire uc_931;
wire uc_932;
wire uc_933;
wire uc_934;
wire uc_935;
wire uc_936;
wire uc_937;
wire uc_938;
wire uc_939;
wire uc_940;
wire uc_941;
wire uc_942;
wire uc_943;
wire uc_944;
wire uc_945;
wire uc_946;
wire uc_947;
wire uc_948;
wire uc_949;
wire uc_950;
wire uc_951;
wire uc_952;
wire uc_953;
wire uc_954;
wire uc_955;
wire uc_956;
wire uc_957;
wire uc_958;
wire uc_959;
wire uc_960;
wire uc_961;
wire uc_962;
wire uc_963;
wire uc_964;
wire uc_965;
wire uc_966;
wire uc_967;
wire uc_968;
wire uc_969;
wire uc_970;
wire uc_971;
wire uc_972;
wire uc_973;
wire uc_974;
wire uc_975;
wire uc_976;
wire uc_977;
wire uc_978;
wire uc_979;
wire uc_980;
wire uc_981;
wire uc_982;
wire uc_983;
wire uc_984;
wire uc_985;
wire uc_986;
wire uc_987;
wire uc_988;
wire uc_989;
wire uc_990;
wire uc_991;
wire uc_992;
wire uc_993;
wire uc_994;
wire uc_995;
wire uc_996;
wire uc_997;
wire uc_998;
wire uc_999;
wire uc_1000;
wire uc_1001;
wire uc_1002;
wire uc_1003;
wire uc_1004;
wire uc_1005;
wire uc_1006;
wire uc_1007;
wire uc_1008;
wire uc_1009;
wire uc_1010;
wire uc_1011;
wire uc_1012;
wire uc_1013;
wire uc_1014;
wire uc_1015;
wire uc_1016;
wire uc_1017;
wire uc_1018;
wire uc_1019;
wire uc_1020;
wire uc_1021;
wire uc_1022;
wire uc_1023;
wire uc_1024;
wire uc_1025;
wire uc_1026;
wire uc_1027;
wire uc_1028;
wire uc_1029;
wire uc_1030;
wire uc_1031;
wire uc_1032;
wire uc_1033;
wire uc_1034;
wire uc_1035;
wire uc_1036;
wire uc_1037;
wire uc_1038;
wire uc_1039;
wire uc_1040;
wire uc_1041;
wire uc_1042;
wire uc_1043;
wire uc_1044;
wire uc_1045;
wire uc_1046;
wire uc_1047;
wire uc_1048;
wire uc_1049;
wire uc_1050;
wire uc_1051;
wire uc_1052;
wire uc_1053;
wire uc_1054;
wire uc_1055;
wire uc_1056;
wire uc_1057;
wire uc_1058;
wire uc_1059;
wire uc_1060;
wire uc_1061;
wire uc_1062;
wire uc_1063;
wire uc_1064;
wire uc_1065;
wire uc_1066;
wire uc_1067;
wire uc_1068;
wire uc_1069;
wire uc_1070;
wire uc_1071;
wire uc_1072;
wire uc_1073;
wire uc_1074;
wire uc_1075;
wire uc_1076;
wire uc_1077;
wire uc_1078;
wire uc_1079;
wire uc_1080;
wire uc_1081;
wire uc_1082;
wire uc_1083;
wire uc_1084;
wire uc_1085;
wire uc_1086;
wire uc_1087;
wire uc_1088;
wire uc_1089;
wire uc_1090;
wire uc_1091;
wire uc_1092;
wire uc_1093;
wire uc_1094;
wire uc_1095;
wire uc_1096;
wire uc_1097;
wire uc_1098;
wire uc_1099;
wire uc_1100;
wire uc_1101;
wire uc_1102;
wire uc_1103;
wire uc_1104;
wire uc_1105;
wire uc_1106;
wire uc_1107;
wire uc_1108;
wire uc_1109;
wire uc_1110;
wire uc_1111;
wire uc_1112;
wire uc_1113;
wire uc_1114;
wire uc_1115;
wire uc_1116;
wire uc_1117;
wire uc_1118;
wire uc_1119;
wire uc_1120;
wire uc_1121;
wire uc_1122;
wire uc_1123;
wire uc_1124;
wire uc_1125;
wire uc_1126;
wire uc_1127;
wire uc_1128;
wire uc_1129;
wire uc_1130;
wire uc_1131;
wire uc_1132;
wire uc_1133;
wire uc_1134;
wire uc_1135;
wire uc_1136;
wire uc_1137;
wire uc_1138;
wire uc_1139;
wire uc_1140;
wire uc_1141;
wire uc_1142;
wire uc_1143;
wire uc_1144;
wire uc_1145;
wire uc_1146;
wire uc_1147;
wire uc_1148;
wire uc_1149;
wire uc_1150;
wire uc_1151;
wire uc_1152;
wire uc_1153;
wire uc_1154;
wire uc_1155;
wire uc_1156;
wire uc_1157;
wire uc_1158;
wire uc_1159;
wire uc_1160;
wire uc_1161;
wire uc_1162;
wire uc_1163;
wire uc_1164;
wire uc_1165;
wire uc_1166;
wire uc_1167;
wire uc_1168;
wire uc_1169;
wire uc_1170;
wire uc_1171;
wire uc_1172;
wire uc_1173;
wire uc_1174;
wire uc_1175;
wire uc_1176;
wire uc_1177;
wire uc_1178;
wire uc_1179;
wire uc_1180;
wire uc_1181;
wire uc_1182;
wire uc_1183;
wire uc_1184;
wire uc_1185;
wire uc_1186;
wire uc_1187;
wire uc_1188;
wire uc_1189;
wire uc_1190;
wire uc_1191;
wire uc_1192;
wire uc_1193;
wire uc_1194;
wire uc_1195;
wire uc_1196;
wire uc_1197;
wire uc_1198;
wire uc_1199;
wire uc_1200;
wire uc_1201;
wire uc_1202;
wire uc_1203;
wire uc_1204;
wire uc_1205;
wire uc_1206;
wire uc_1207;
wire uc_1208;
wire uc_1209;
wire uc_1210;
wire uc_1211;
wire uc_1212;
wire uc_1213;
wire uc_1214;
wire uc_1215;
wire uc_1216;
wire uc_1217;
wire uc_1218;
wire uc_1219;
wire uc_1220;
wire uc_1221;
wire uc_1222;
wire uc_1223;
wire uc_1224;
wire uc_1225;
wire uc_1226;
wire uc_1227;
wire uc_1228;
wire uc_1229;
wire uc_1230;
wire uc_1231;
wire uc_1232;
wire uc_1233;
wire uc_1234;
wire uc_1235;
wire uc_1236;
wire uc_1237;
wire uc_1238;
wire uc_1239;
wire uc_1240;
wire uc_1241;
wire uc_1242;
wire uc_1243;
wire uc_1244;
wire uc_1245;
wire uc_1246;
wire uc_1247;
wire uc_1248;
wire uc_1249;
wire uc_1250;
wire uc_1251;
wire uc_1252;
wire uc_1253;
wire uc_1254;
wire uc_1255;
wire uc_1256;
wire uc_1257;
wire uc_1258;
wire uc_1259;
wire uc_1260;
wire uc_1261;
wire uc_1262;
wire uc_1263;
wire uc_1264;
wire uc_1265;
wire uc_1266;
wire uc_1267;
wire uc_1268;
wire uc_1269;
wire uc_1270;
wire uc_1271;
wire uc_1272;
wire uc_1273;
wire uc_1274;
wire uc_1275;
wire uc_1276;
wire uc_1277;
wire uc_1278;
wire uc_1279;
wire uc_1280;
wire uc_1281;
wire uc_1282;
wire uc_1283;
wire uc_1284;
wire uc_1285;
wire uc_1286;
wire uc_1287;
wire uc_1288;
wire uc_1289;
wire uc_1290;
wire uc_1291;
wire uc_1292;
wire uc_1293;
wire uc_1294;
wire uc_1295;
wire uc_1296;
wire uc_1297;
wire uc_1298;
wire uc_1299;
wire uc_1300;
wire uc_1301;
wire uc_1302;
wire uc_1303;
wire uc_1304;
wire uc_1305;
wire uc_1306;
wire uc_1307;
wire uc_1308;
wire uc_1309;
wire uc_1310;
wire uc_1311;
wire uc_1312;
wire uc_1313;
wire uc_1314;
wire uc_1315;
wire uc_1316;
wire uc_1317;
wire uc_1318;
wire uc_1319;
wire uc_1320;
wire uc_1321;
wire uc_1322;
wire uc_1323;
wire uc_1324;
wire uc_1325;
wire uc_1326;
wire uc_1327;
wire uc_1328;
wire uc_1329;
wire uc_1330;
wire uc_1331;
wire uc_1332;
wire uc_1333;
wire uc_1334;
wire uc_1335;
wire uc_1336;
wire uc_1337;
wire uc_1338;
wire uc_1339;
wire uc_1340;
wire uc_1341;
wire uc_1342;
wire uc_1343;
wire uc_1344;
wire uc_1345;
wire uc_1346;
wire uc_1347;
wire uc_1348;
wire uc_1349;
wire uc_1350;
wire uc_1351;
wire uc_1352;
wire uc_1353;
wire uc_1354;
wire uc_1355;
wire uc_1356;
wire uc_1357;
wire uc_1358;
wire uc_1359;
wire uc_1360;
wire uc_1361;
wire uc_1362;
wire uc_1363;
wire uc_1364;
wire uc_1365;
wire uc_1366;
wire uc_1367;
wire uc_1368;
wire uc_1369;
wire uc_1370;
wire uc_1371;
wire uc_1372;
wire uc_1373;
wire uc_1374;
wire uc_1375;
wire uc_1376;
wire uc_1377;
wire uc_1378;
wire uc_1379;
wire uc_1380;
wire uc_1381;
wire uc_1382;
wire uc_1383;
wire uc_1384;
wire uc_1385;
wire uc_1386;
wire uc_1387;
wire uc_1388;
wire uc_1389;
wire uc_1390;
wire uc_1391;
wire uc_1392;
wire uc_1393;
wire uc_1394;
wire uc_1395;
wire uc_1396;
wire uc_1397;
wire uc_1398;
wire uc_1399;
wire uc_1400;
wire uc_1401;
wire uc_1402;
wire uc_1403;
wire uc_1404;
wire uc_1405;
wire uc_1406;
wire uc_1407;
wire uc_1408;
wire uc_1409;
wire uc_1410;
wire uc_1411;
wire uc_1412;
wire uc_1413;
wire uc_1414;
wire uc_1415;
wire uc_1416;
wire uc_1417;
wire uc_1418;
wire uc_1419;
wire uc_1420;
wire uc_1421;
wire uc_1422;
wire uc_1423;
wire uc_1424;
wire uc_1425;
wire uc_1426;
wire uc_1427;
wire uc_1428;
wire uc_1429;
wire uc_1430;
wire uc_1431;
wire uc_1432;
wire uc_1433;
wire uc_1434;
wire uc_1435;
wire uc_1436;
wire uc_1437;
wire uc_1438;
wire uc_1439;
wire uc_1440;
wire uc_1441;
wire uc_1442;
wire uc_1443;
wire uc_1444;
wire uc_1445;
wire uc_1446;
wire uc_1447;
wire uc_1448;
wire uc_1449;
wire uc_1450;
wire uc_1451;
wire uc_1452;
wire uc_1453;
wire uc_1454;
wire uc_1455;
wire uc_1456;
wire uc_1457;
wire uc_1458;
wire uc_1459;
wire uc_1460;
wire uc_1461;
wire uc_1462;
wire uc_1463;
wire uc_1464;
wire uc_1465;
wire uc_1466;
wire uc_1467;
wire uc_1468;
wire uc_1469;
wire uc_1470;
wire uc_1471;
wire uc_1472;
wire uc_1473;
wire uc_1474;
wire uc_1475;
wire uc_1476;
wire uc_1477;
wire uc_1478;
wire uc_1479;
wire uc_1480;
wire uc_1481;
wire uc_1482;
wire uc_1483;
wire uc_1484;
wire uc_1485;
wire uc_1486;
wire uc_1487;
wire uc_1488;
wire uc_1489;
wire uc_1490;
wire uc_1491;
wire uc_1492;
wire uc_1493;
wire uc_1494;
wire uc_1495;
wire uc_1496;
wire uc_1497;
wire uc_1498;
wire uc_1499;
wire uc_1500;
wire uc_1501;
wire uc_1502;
wire uc_1503;
wire uc_1504;
wire uc_1505;
wire uc_1506;
wire uc_1507;
wire uc_1508;
wire uc_1509;
wire uc_1510;
wire uc_1511;
wire uc_1512;
wire uc_1513;
wire uc_1514;
wire uc_1515;
wire uc_1516;
wire uc_1517;
wire uc_1518;
wire uc_1519;
wire uc_1520;
wire uc_1521;
wire uc_1522;
wire uc_1523;
wire uc_1524;
wire uc_1525;
wire uc_1526;
wire uc_1527;
wire uc_1528;
wire uc_1529;
wire uc_1530;
wire uc_1531;
wire uc_1532;
wire uc_1533;
wire uc_1534;
wire uc_1535;
wire uc_1536;
wire uc_1537;
wire uc_1538;
wire uc_1539;
wire uc_1540;
wire uc_1541;
wire uc_1542;
wire uc_1543;
wire uc_1544;
wire uc_1545;
wire uc_1546;
wire uc_1547;
wire uc_1548;
wire uc_1549;
wire uc_1550;
wire uc_1551;
wire uc_1552;
wire uc_1553;
wire uc_1554;
wire uc_1555;
wire uc_1556;
wire uc_1557;
wire uc_1558;
wire uc_1559;
wire uc_1560;
wire uc_1561;
wire uc_1562;
wire uc_1563;
wire uc_1564;
wire uc_1565;
wire uc_1566;
wire uc_1567;
wire uc_1568;
wire uc_1569;
wire uc_1570;
wire uc_1571;
wire uc_1572;
wire uc_1573;
wire uc_1574;
wire uc_1575;
wire uc_1576;
wire uc_1577;
wire uc_1578;
wire uc_1579;
wire uc_1580;
wire uc_1581;
wire uc_1582;
wire uc_1583;
wire uc_1584;
wire uc_1585;
wire uc_1586;
wire uc_1587;
wire uc_1588;
wire uc_1589;
wire uc_1590;
wire uc_1591;
wire uc_1592;
wire uc_1593;
wire uc_1594;
wire uc_1595;
wire uc_1596;
wire uc_1597;
wire uc_1598;
wire uc_1599;
wire uc_1600;
wire uc_1601;
wire uc_1602;
wire uc_1603;
wire uc_1604;
wire uc_1605;
wire uc_1606;
wire uc_1607;
wire uc_1608;
wire uc_1609;
wire uc_1610;
wire uc_1611;
wire uc_1612;
wire uc_1613;
wire uc_1614;
wire uc_1615;
wire uc_1616;
wire uc_1617;
wire uc_1618;
wire uc_1619;
wire uc_1620;
wire uc_1621;
wire uc_1622;
wire uc_1623;
wire uc_1624;
wire uc_1625;
wire uc_1626;
wire uc_1627;
wire uc_1628;
wire uc_1629;
wire uc_1630;
wire uc_1631;
wire uc_1632;
wire uc_1633;
wire uc_1634;
wire uc_1635;
wire uc_1636;
wire uc_1637;
wire uc_1638;
wire uc_1639;
wire uc_1640;
wire uc_1641;
wire uc_1642;
wire uc_1643;
wire uc_1644;
wire uc_1645;
wire uc_1646;
wire uc_1647;
wire uc_1648;
wire uc_1649;
wire uc_1650;
wire uc_1651;
wire uc_1652;
wire uc_1653;
wire uc_1654;
wire uc_1655;
wire uc_1656;
wire uc_1657;
wire uc_1658;
wire uc_1659;
wire uc_1660;
wire uc_1661;
wire uc_1662;
wire uc_1663;
wire uc_1664;
wire uc_1665;
wire uc_1666;
wire uc_1667;
wire uc_1668;
wire uc_1669;
wire uc_1670;
wire uc_1671;
wire uc_1672;
wire uc_1673;
wire uc_1674;
wire uc_1675;
wire uc_1676;
wire uc_1677;
wire uc_1678;
wire uc_1679;
wire uc_1680;
wire uc_1681;
wire uc_1682;
wire uc_1683;
wire uc_1684;
wire uc_1685;
wire uc_1686;
wire uc_1687;
wire uc_1688;
wire uc_1689;
wire uc_1690;
wire uc_1691;
wire uc_1692;
wire uc_1693;
wire uc_1694;
wire uc_1695;
wire uc_1696;
wire uc_1697;
wire uc_1698;
wire uc_1699;
wire uc_1700;
wire uc_1701;
wire uc_1702;
wire uc_1703;
wire uc_1704;
wire uc_1705;
wire uc_1706;
wire uc_1707;
wire uc_1708;
wire uc_1709;
wire uc_1710;
wire uc_1711;
wire uc_1712;
wire uc_1713;
wire uc_1714;
wire uc_1715;
wire uc_1716;
wire uc_1717;
wire uc_1718;
wire uc_1719;
wire uc_1720;
wire uc_1721;
wire uc_1722;
wire uc_1723;
wire uc_1724;
wire uc_1725;
wire uc_1726;
wire uc_1727;
wire uc_1728;
wire uc_1729;
wire uc_1730;
wire uc_1731;
wire uc_1732;
wire uc_1733;
wire uc_1734;
wire uc_1735;
wire uc_1736;
wire uc_1737;
wire uc_1738;
wire uc_1739;
wire uc_1740;
wire uc_1741;
wire uc_1742;
wire uc_1743;
wire uc_1744;
wire uc_1745;
wire uc_1746;
wire uc_1747;
wire uc_1748;
wire uc_1749;
wire uc_1750;
wire uc_1751;
wire uc_1752;
wire uc_1753;
wire uc_1754;
wire uc_1755;
wire uc_1756;
wire uc_1757;
wire uc_1758;
wire uc_1759;
wire uc_1760;
wire uc_1761;
wire uc_1762;
wire uc_1763;
wire uc_1764;
wire uc_1765;
wire uc_1766;
wire uc_1767;
wire uc_1768;
wire uc_1769;
wire uc_1770;
wire uc_1771;
wire uc_1772;
wire uc_1773;
wire uc_1774;
wire uc_1775;
wire uc_1776;
wire uc_1777;
wire uc_1778;
wire uc_1779;
wire uc_1780;
wire uc_1781;
wire uc_1782;
wire uc_1783;
wire uc_1784;
wire uc_1785;
wire uc_1786;
wire uc_1787;
wire uc_1788;
wire uc_1789;
wire uc_1790;
wire uc_1791;
wire uc_1792;
wire uc_1793;
wire uc_1794;
wire uc_1795;
wire uc_1796;
wire uc_1797;
wire uc_1798;
wire uc_1799;
wire uc_1800;
wire uc_1801;
wire uc_1802;
wire uc_1803;
wire uc_1804;
wire uc_1805;
wire uc_1806;
wire uc_1807;
wire uc_1808;
wire uc_1809;
wire uc_1810;
wire uc_1811;
wire uc_1812;
wire uc_1813;
wire uc_1814;
wire uc_1815;
wire uc_1816;
wire uc_1817;
wire uc_1818;
wire uc_1819;
wire uc_1820;
wire uc_1821;
wire uc_1822;
wire uc_1823;
wire uc_1824;
wire uc_1825;
wire uc_1826;
wire uc_1827;
wire uc_1828;
wire uc_1829;
wire uc_1830;
wire uc_1831;
wire uc_1832;
wire uc_1833;
wire uc_1834;
wire uc_1835;
wire uc_1836;
wire uc_1837;
wire uc_1838;
wire uc_1839;
wire uc_1840;
wire uc_1841;
wire uc_1842;
wire uc_1843;
wire uc_1844;
wire uc_1845;
wire uc_1846;
wire uc_1847;
wire uc_1848;
wire uc_1849;
wire uc_1850;
wire uc_1851;
wire uc_1852;
wire uc_1853;
wire uc_1854;
wire uc_1855;
wire uc_1856;
wire uc_1857;
wire uc_1858;
wire uc_1859;
wire uc_1860;
wire uc_1861;
wire uc_1862;
wire uc_1863;
wire uc_1864;
wire uc_1865;
wire uc_1866;
wire uc_1867;
wire uc_1868;
wire uc_1869;
wire uc_1870;
wire uc_1871;
wire uc_1872;
wire uc_1873;
wire uc_1874;
wire uc_1875;
wire uc_1876;
wire uc_1877;
wire uc_1878;
wire uc_1879;
wire uc_1880;
wire uc_1881;
wire uc_1882;
wire uc_1883;
wire uc_1884;
wire uc_1885;
wire uc_1886;
wire uc_1887;
wire uc_1888;
wire uc_1889;
wire uc_1890;
wire uc_1891;
wire uc_1892;
wire uc_1893;
wire uc_1894;
wire uc_1895;
wire uc_1896;
wire uc_1897;
wire uc_1898;
wire uc_1899;
wire uc_1900;
wire uc_1901;
wire uc_1902;
wire uc_1903;
wire uc_1904;
wire uc_1905;
wire uc_1906;
wire uc_1907;
wire uc_1908;
wire uc_1909;
wire uc_1910;
wire uc_1911;
wire uc_1912;
wire uc_1913;
wire uc_1914;
wire uc_1915;
wire uc_1916;
wire uc_1917;
wire uc_1918;
wire uc_1919;
wire uc_1920;
wire uc_1921;
wire uc_1922;
wire uc_1923;
wire uc_1924;
wire uc_1925;
wire uc_1926;
wire uc_1927;
wire uc_1928;
wire uc_1929;
wire uc_1930;
wire uc_1931;
wire uc_1932;
wire uc_1933;
wire uc_1934;
wire uc_1935;
wire uc_1936;
wire uc_1937;
wire uc_1938;
wire uc_1939;
wire uc_1940;
wire uc_1941;
wire uc_1942;
wire uc_1943;
wire uc_1944;
wire uc_1945;
wire uc_1946;
wire uc_1947;
wire uc_1948;
wire uc_1949;
wire uc_1950;
wire uc_1951;
wire uc_1952;
wire uc_1953;
wire uc_1954;
wire uc_1955;
wire uc_1956;
wire uc_1957;
wire uc_1958;
wire uc_1959;
wire uc_1960;
wire uc_1961;
wire uc_1962;
wire uc_1963;
wire uc_1964;
wire uc_1965;
wire uc_1966;
wire uc_1967;
wire uc_1968;
wire uc_1969;
wire uc_1970;
wire uc_1971;
wire uc_1972;
wire uc_1973;
wire uc_1974;
wire uc_1975;
wire uc_1976;
wire uc_1977;
wire uc_1978;
wire uc_1979;
wire uc_1980;
wire uc_1981;
wire uc_1982;
wire uc_1983;
wire uc_1984;
wire uc_1985;
wire uc_1986;
wire uc_1987;
wire uc_1988;
wire uc_1989;
wire uc_1990;
wire uc_1991;
wire uc_1992;
wire uc_1993;
wire uc_1994;
wire uc_1995;
wire uc_1996;
wire uc_1997;
wire uc_1998;
wire uc_1999;
wire uc_2000;
wire uc_2001;
wire uc_2002;
wire uc_2003;
wire uc_2004;
wire uc_2005;
wire uc_2006;
wire uc_2007;
wire uc_2008;
wire uc_2009;
wire uc_2010;
wire uc_2011;
wire uc_2012;
wire uc_2013;
wire uc_2014;
wire uc_2015;
wire uc_2016;
wire uc_2017;
wire uc_2018;
wire uc_2019;
wire uc_2020;
wire uc_2021;
wire uc_2022;
wire uc_2023;
wire uc_2024;
wire uc_2025;
wire uc_2026;
wire uc_2027;
wire uc_2028;
wire uc_2029;
wire uc_2030;
wire uc_2031;
wire uc_2032;
wire uc_2033;
wire uc_2034;
wire uc_2035;
wire uc_2036;
wire uc_2037;
wire uc_2038;
wire uc_2039;
wire uc_2040;
wire uc_2041;
wire uc_2042;
wire uc_2043;
wire uc_2044;
wire uc_2045;
wire uc_2046;
wire uc_2047;
wire uc_2048;
wire uc_2049;
wire uc_2050;
wire uc_2051;
wire uc_2052;
wire uc_2053;
wire uc_2054;
wire uc_2055;
wire uc_2056;
wire uc_2057;
wire uc_2058;
wire uc_2059;
wire uc_2060;
wire uc_2061;
wire uc_2062;
wire uc_2063;
wire uc_2064;
wire uc_2065;
wire uc_2066;
wire uc_2067;
wire uc_2068;
wire uc_2069;
wire uc_2070;
wire uc_2071;
wire uc_2072;
wire uc_2073;
wire uc_2074;
wire uc_2075;
wire uc_2076;
wire uc_2077;
wire uc_2078;
wire uc_2079;
wire uc_2080;
wire uc_2081;
wire uc_2082;
wire uc_2083;
wire uc_2084;
wire uc_2085;
wire uc_2086;
wire uc_2087;
wire uc_2088;
wire uc_2089;
wire uc_2090;
wire uc_2091;
wire uc_2092;
wire uc_2093;
wire uc_2094;
wire uc_2095;
wire uc_2096;
wire uc_2097;
wire uc_2098;
wire uc_2099;
wire uc_2100;
wire uc_2101;
wire uc_2102;
wire uc_2103;
wire uc_2104;
wire uc_2105;
wire uc_2106;
wire uc_2107;
wire uc_2108;
wire uc_2109;
wire uc_2110;
wire uc_2111;
wire uc_2112;
wire uc_2113;
wire uc_2114;
wire uc_2115;
wire uc_2116;
wire uc_2117;
wire uc_2118;
wire uc_2119;
wire uc_2120;
wire uc_2121;
wire uc_2122;
wire uc_2123;
wire uc_2124;
wire uc_2125;
wire uc_2126;
wire uc_2127;
wire uc_2128;
wire uc_2129;
wire uc_2130;
wire uc_2131;
wire uc_2132;
wire uc_2133;
wire uc_2134;
wire uc_2135;
wire uc_2136;
wire uc_2137;
wire uc_2138;
wire uc_2139;
wire uc_2140;
wire uc_2141;
wire uc_2142;
wire uc_2143;
wire uc_2144;
wire uc_2145;
wire uc_2146;
wire uc_2147;
wire uc_2148;
wire uc_2149;
wire uc_2150;
wire uc_2151;
wire uc_2152;
wire uc_2153;
wire uc_2154;
wire uc_2155;
wire uc_2156;
wire uc_2157;
wire uc_2158;
wire uc_2159;
wire uc_2160;
wire uc_2161;


NAND2_X4 slo__sro_c506 (.ZN (slo__sro_n363), .A1 (slo__sro_n365), .A2 (slo__sro_n364));
INV_X8 opt_ipo_c1781 (.ZN (opt_ipo_n1524), .A (opt_ipo_n1551));
NAND2_X4 slo__sro_c706 (.ZN (slo__sro_n540), .A1 (n_0_140), .A2 (drc_ipo_n26));
NOR4_X2 i_0_1_288 (.ZN (n_0_1_144), .A1 (\Res_imm[47] ), .A2 (\Res_imm[41] ), .A3 (\Res_imm[42] ), .A4 (\Res_imm[44] ));
NOR4_X1 i_0_1_287 (.ZN (n_0_1_143), .A1 (\Res_imm[35] ), .A2 (\Res_imm[32] ), .A3 (\Res_imm[38] ), .A4 (\Res_imm[37] ));
NOR4_X4 i_0_1_286 (.ZN (n_0_1_142), .A1 (CLOCK_slo___n3239), .A2 (\Res_imm[56] ), .A3 (\Res_imm[62] ), .A4 (\Res_imm[61] ));
NOR4_X4 i_0_1_285 (.ZN (n_0_1_76), .A1 (\Res_imm[52] ), .A2 (\Res_imm[49] ), .A3 (\Res_imm[55] ), .A4 (\Res_imm[50] ));
NAND2_X1 CLOCK_slo__sro_c3057 (.ZN (CLOCK_slo__sro_n2683), .A1 (n_0_77), .A2 (CLOCK_slo__sro_n2685));
NOR4_X1 i_0_1_283 (.ZN (n_0_1_74), .A1 (\Res_imm[14] ), .A2 (\Res_imm[13] ), .A3 (\Res_imm[11] ), .A4 (\secondStage_Res[8] ));
NOR4_X1 i_0_1_282 (.ZN (n_0_1_73), .A1 (\secondStage_Res[2] ), .A2 (\secondStage_Res[1] )
    , .A3 (\secondStage_Res[7] ), .A4 (\secondStage_Res[4] ));
NOR4_X2 i_0_1_281 (.ZN (n_0_1_71), .A1 (CLOCK_slo___n2653), .A2 (\Res_imm[25] ), .A3 (\Res_imm[31] ), .A4 (\Res_imm[26] ));
NOR4_X1 i_0_1_280 (.ZN (n_0_1_70), .A1 (\Res_imm[19] ), .A2 (\Res_imm[16] ), .A3 (\Res_imm[22] ), .A4 (\Res_imm[21] ));
OR2_X1 sgo__sro_c332 (.ZN (sgo__sro_n246), .A1 (\Res_imm[34] ), .A2 (\Res_imm[33] ));
OAI21_X4 CLOCK_slo__mro_c2637 (.ZN (CLOCK_slo__mro_n2292), .A (slo__sro_n1131), .B1 (n_0_139), .B2 (slo__sro_n1132));
NAND2_X1 slo__sro_c505 (.ZN (slo__sro_n364), .A1 (n_0_103), .A2 (slo__sro_n366));
INV_X1 slo__sro_c545 (.ZN (slo__sro_n408), .A (drc_ipo_n26));
NAND2_X2 CLOCK_slo__sro_c2647 (.ZN (CLOCK_slo__sro_n2300), .A1 (n_0_167), .A2 (drc_ipo_n27));
NAND2_X2 sgo__sro_c202 (.ZN (n_0_1_69), .A1 (n_0_1_71), .A2 (sgo__sro_n145));
NOR4_X1 i_0_1_257 (.ZN (n_0_1_23), .A1 (\Res_imm[10] ), .A2 (\Res_imm[9] ), .A3 (\Res_imm[15] ), .A4 (\Res_imm[12] ));
NOR4_X1 i_0_1_256 (.ZN (n_0_1_22), .A1 (\secondStage_Res[3] ), .A2 (n_0_316), .A3 (\secondStage_Res[6] ), .A4 (\secondStage_Res[5] ));
INV_X1 slo__sro_c705 (.ZN (slo__sro_n541), .A (drc_ipo_n26));
NOR4_X1 i_0_1_254 (.ZN (n_0_1_20), .A1 (\Res_imm[18] ), .A2 (\Res_imm[17] ), .A3 (\Res_imm[23] ), .A4 (\Res_imm[20] ));
NAND4_X1 i_0_1_253 (.ZN (n_0_1_19), .A1 (n_0_1_20), .A2 (n_0_1_22), .A3 (n_0_1_21), .A4 (n_0_1_23));
INV_X1 slo__sro_c503 (.ZN (slo__sro_n366), .A (drc_ipo_n26));
XNOR2_X2 i_0_1_242 (.ZN (n_0_1_17), .A (drc_ipo_n26), .B (drc_ipo_n27));
NAND2_X4 slo__sro_c1290 (.ZN (slo__sro_n1081), .A1 (n_0_138), .A2 (drc_ipo_n26));
CLKBUF_X3 hfn_ipo_c22 (.Z (hfn_ipo_n22), .A (n_0_1_5));
INV_X2 sgo__sro_c38 (.ZN (sgo__sro_n35), .A (n_0_49));
BUF_X16 hfn_ipo_c24 (.Z (hfn_ipo_n24), .A (slo__n798));
XNOR2_X2 i_0_1_223 (.ZN (OVF), .A (n_0_1_13), .B (B[31]));
NAND2_X4 i_0_1_217 (.ZN (n_0_1_13), .A1 (opt_ipo_n1380), .A2 (CLOCK_opt_ipo_n1683));
OR2_X2 CLOCK_sgo__sro_c2217 (.ZN (CLOCK_sgo__sro_n1959), .A1 (\Res_imm[54] ), .A2 (\Res_imm[53] ));
MUX2_X2 i_0_1_366 (.Z (\A_imm[27] ), .A (n_0_96), .B (n_0_149), .S (drc_ipo_n26));
INV_X1 slo__sro_c725 (.ZN (slo__sro_n561), .A (drc_ipo_n26));
INV_X1 slo__sro_c563 (.ZN (slo__sro_n423), .A (drc_ipo_n27));
MUX2_X2 i_0_1_363 (.Z (slo__n378), .A (n_0_101), .B (n_0_144), .S (drc_ipo_n26));
INV_X1 slo__sro_c875 (.ZN (slo__sro_n703), .A (drc_ipo_n27));
BUF_X8 slo__c518 (.Z (\A_imm[22] ), .A (slo__n378));
AND2_X4 slo__mro_c531 (.ZN (slo__mro_n394), .A1 (n_0_1_68), .A2 (n_0_1_28));
INV_X1 slo__sro_c1350 (.ZN (slo__sro_n1153), .A (drc_ipo_n27));
INV_X1 slo__sro_c1326 (.ZN (slo__sro_n1123), .A (drc_ipo_n26));
INV_X1 slo__sro_c1289 (.ZN (slo__sro_n1082), .A (drc_ipo_n26));
INV_X1 CLOCK_slo__sro_c2538 (.ZN (CLOCK_slo__sro_n2215), .A (drc_ipo_n27));
INV_X1 slo__sro_c1336 (.ZN (slo__sro_n1133), .A (drc_ipo_n26));
MUX2_X2 i_0_1_350 (.Z (\A_imm[12] ), .A (n_0_111), .B (n_0_134), .S (drc_ipo_n26));
MUX2_X2 i_0_1_341 (.Z (\A_imm[11] ), .A (n_0_112), .B (n_0_133), .S (drc_ipo_n26));
INV_X1 slo__sro_c844 (.ZN (slo__sro_n670), .A (drc_ipo_n26));
MUX2_X2 i_0_1_339 (.Z (\A_imm[9] ), .A (n_0_114), .B (n_0_131), .S (drc_ipo_n26));
MUX2_X2 i_0_1_338 (.Z (\A_imm[8] ), .A (n_0_115), .B (n_0_130), .S (drc_ipo_n26));
MUX2_X2 i_0_1_337 (.Z (\A_imm[7] ), .A (n_0_116), .B (n_0_129), .S (drc_ipo_n26));
MUX2_X2 i_0_1_336 (.Z (\A_imm[6] ), .A (n_0_117), .B (n_0_128), .S (drc_ipo_n26));
MUX2_X2 i_0_1_330 (.Z (\A_imm[5] ), .A (n_0_118), .B (n_0_127), .S (drc_ipo_n26));
INV_X1 slo__sro_c673 (.ZN (slo__sro_n516), .A (drc_ipo_n27));
CLKBUF_X3 CTS_L1_c_tid0_2005 (.Z (CTS_n_tid0_1747), .A (clk));
INV_X1 CLOCK_slo__sro_c2646 (.ZN (CLOCK_slo__sro_n2301), .A (drc_ipo_n27));
AOI21_X4 CLOCK_slo__mro_c3590 (.ZN (CLOCK_slo__mro_n3163), .A (CLOCK_slo__mro_n3164)
    , .B1 (n_0_148), .B2 (drc_ipo_n26));
NAND2_X4 i_0_1_318 (.ZN (n_0_315), .A1 (CTS_n_tid0_1747), .A2 (hfn_ipo_n22));
INV_X4 CTS_L3_remove_c1990 (.ZN (CTS_n1730), .A (CTS_n1731));
AOI21_X1 i_0_1_316 (.ZN (CTS_n1731), .A (reset), .B1 (CLOCK_slh_n3498), .B2 (CTS_n_tid0_1747));
INV_X1 i_0_1_275 (.ZN (n_0_247), .A (n_0_1_10));
AOI22_X2 i_0_1_274 (.ZN (n_0_1_10), .A1 (opt_ipo_n1555), .A2 (opt_ipo_n1365), .B1 (n_0_61), .B2 (slo__xsl_n298));
CLKBUF_X1 CLOCK_slo___L1_c1_c3023 (.Z (\Res_imm[28] ), .A (CLOCK_slo___n2653));
AOI22_X2 i_0_1_270 (.ZN (n_0_1_9), .A1 (opt_ipo_n1555), .A2 (\Res_imm[60] ), .B1 (slo__xsl_n298), .B2 (n_0_59));
INV_X1 i_0_1_269 (.ZN (n_0_242), .A (n_0_1_8));
AOI22_X2 i_0_1_268 (.ZN (n_0_1_8), .A1 (opt_ipo_n1555), .A2 (\Res_imm[57] ), .B1 (n_0_56), .B2 (slo__xsl_n298));
INV_X1 i_0_1_267 (.ZN (n_0_236), .A (n_0_1_7));
AOI22_X1 i_0_1_265 (.ZN (n_0_1_7), .A1 (opt_ipo_n1555), .A2 (\Res_imm[51] ), .B1 (slo__xsl_n298), .B2 (n_0_50));
INV_X1 i_0_1_264 (.ZN (n_0_235), .A (n_0_1_6));
NAND2_X2 CLOCK_slo__sro_c2539 (.ZN (CLOCK_slo__sro_n2214), .A1 (n_0_159), .A2 (drc_ipo_n27));
INV_X1 i_0_1_183 (.ZN (n_0_1_5), .A (reset));
BUF_X8 hfn_ipo_c23 (.Z (hfn_ipo_n23), .A (n_0_1_5));
INV_X2 opt_ipo_c1909 (.ZN (opt_ipo_n1652), .A (slo__n980));
AOI22_X2 i_0_1_15 (.ZN (n_0_1_24), .A1 (n_0_54), .A2 (slo__xsl_n298), .B1 (opt_ipo_n1555), .B2 (\Res_imm[55] ));
INV_X1 i_0_1_360 (.ZN (n_0_1_4), .A (n_0_58));
NAND2_X2 i_0_1_359 (.ZN (n_0_1_3), .A1 (opt_ipo_n1555), .A2 (\Res_imm[59] ));
OAI21_X1 i_0_1_358 (.ZN (n_0_244), .A (n_0_1_3), .B1 (n_0_1_4), .B2 (hfn_ipo_n25));
NAND2_X1 i_0_1_150 (.ZN (n_0_1_2), .A1 (opt_ipo_n1555), .A2 (\Res_imm[63] ));
NAND2_X1 slo__sro_c707 (.ZN (slo__sro_n539), .A1 (n_0_105), .A2 (slo__sro_n541));
NAND2_X1 i_0_1_346 (.ZN (n_0_1_1), .A1 (opt_ipo_n1555), .A2 (CLOCK_opt_ipo_n1670));
NAND2_X1 i_0_1_345 (.ZN (n_0_1_0), .A1 (n_0_60), .A2 (slo__xsl_n298));
NAND2_X1 i_0_1_344 (.ZN (n_0_246), .A1 (n_0_1_0), .A2 (n_0_1_1));
OR2_X1 CLOCK_slo__sro_c3035 (.ZN (CLOCK_slo__sro_n2663), .A1 (n_0_1_17), .A2 (reset));
NAND2_X2 slo__sro_c504 (.ZN (slo__sro_n365), .A1 (n_0_142), .A2 (drc_ipo_n26));
INV_X1 i_0_1_333 (.ZN (n_0_1_153), .A (n_0_55));
NAND2_X1 i_0_1_332 (.ZN (n_0_1_152), .A1 (opt_ipo_n1555), .A2 (\Res_imm[56] ));
OAI21_X1 i_0_1_331 (.ZN (n_0_241), .A (n_0_1_152), .B1 (n_0_1_153), .B2 (hfn_ipo_n25));
INV_X1 i_0_1_327 (.ZN (n_0_1_149), .A (n_0_53));
NAND2_X2 i_0_1_326 (.ZN (n_0_1_148), .A1 (opt_ipo_n1555), .A2 (\Res_imm[54] ));
OAI21_X1 i_0_1_325 (.ZN (n_0_239), .A (n_0_1_148), .B1 (n_0_1_149), .B2 (hfn_ipo_n25));
INV_X1 i_0_1_324 (.ZN (n_0_1_147), .A (n_0_52));
NAND2_X2 i_0_1_323 (.ZN (n_0_1_146), .A1 (opt_ipo_n1555), .A2 (\Res_imm[53] ));
OAI21_X1 i_0_1_322 (.ZN (n_0_238), .A (n_0_1_146), .B1 (n_0_1_147), .B2 (hfn_ipo_n25));
INV_X1 i_0_1_315 (.ZN (n_0_1_141), .A (n_0_48));
NAND2_X2 i_0_1_314 (.ZN (n_0_1_140), .A1 (opt_ipo_n1551), .A2 (\Res_imm[49] ));
OAI21_X1 i_0_1_313 (.ZN (n_0_234), .A (n_0_1_140), .B1 (n_0_1_141), .B2 (hfn_ipo_n25));
INV_X1 i_0_1_147 (.ZN (n_0_1_139), .A (n_0_37));
NAND2_X2 i_0_1_146 (.ZN (n_0_1_138), .A1 (opt_ipo_n1555), .A2 (\Res_imm[38] ));
OAI21_X2 i_0_1_145 (.ZN (n_0_222), .A (n_0_1_138), .B1 (n_0_1_139), .B2 (hfn_ipo_n25));
BUF_X1 CLOCK_opt_ipo_c1927 (.Z (CLOCK_opt_ipo_n1670), .A (\Res_imm[61] ));
INV_X1 i_0_1_308 (.ZN (n_0_1_136), .A (n_0_57));
NAND2_X1 i_0_1_307 (.ZN (n_0_1_135), .A1 (CLOCK_slo__n3265), .A2 (\Res_imm[58] ));
OAI21_X1 i_0_1_306 (.ZN (n_0_243), .A (n_0_1_135), .B1 (n_0_1_136), .B2 (hfn_ipo_n25));
INV_X1 i_0_1_305 (.ZN (n_0_1_134), .A (\Res_imm[52] ));
INV_X1 i_0_1_304 (.ZN (n_0_1_133), .A (n_0_51));
OAI22_X1 i_0_1_303 (.ZN (n_0_237), .A1 (slo__n453), .A2 (n_0_1_134), .B1 (hfn_ipo_n25), .B2 (n_0_1_133));
INV_X1 i_0_1_302 (.ZN (n_0_1_132), .A (opt_ipo_n1361));
INV_X1 i_0_1_301 (.ZN (n_0_1_131), .A (n_0_47));
OAI22_X1 i_0_1_300 (.ZN (n_0_233), .A1 (slo__n453), .A2 (n_0_1_132), .B1 (hfn_ipo_n25), .B2 (n_0_1_131));
INV_X1 i_0_1_143 (.ZN (n_0_1_130), .A (\Res_imm[47] ));
INV_X1 i_0_1_142 (.ZN (n_0_1_129), .A (n_0_46));
OAI22_X1 i_0_1_141 (.ZN (n_0_232), .A1 (slo__n453), .A2 (n_0_1_130), .B1 (hfn_ipo_n25), .B2 (n_0_1_129));
INV_X1 i_0_1_140 (.ZN (n_0_1_128), .A (\Res_imm[46] ));
INV_X1 i_0_1_139 (.ZN (n_0_1_127), .A (n_0_45));
OAI22_X1 i_0_1_138 (.ZN (n_0_231), .A1 (slo__n453), .A2 (n_0_1_128), .B1 (hfn_ipo_n25), .B2 (n_0_1_127));
INV_X1 i_0_1_137 (.ZN (n_0_1_126), .A (\Res_imm[45] ));
INV_X1 i_0_1_136 (.ZN (n_0_1_125), .A (n_0_44));
INV_X1 slo__sro_c1198 (.ZN (slo__sro_n1001), .A (drc_ipo_n26));
INV_X1 i_0_1_134 (.ZN (n_0_1_124), .A (\Res_imm[44] ));
INV_X1 i_0_1_133 (.ZN (n_0_1_123), .A (n_0_43));
OAI22_X2 i_0_1_132 (.ZN (n_0_229), .A1 (slo__n453), .A2 (n_0_1_124), .B1 (hfn_ipo_n25), .B2 (n_0_1_123));
INV_X1 i_0_1_131 (.ZN (n_0_1_122), .A (\Res_imm[43] ));
INV_X1 i_0_1_130 (.ZN (n_0_1_121), .A (n_0_42));
OAI22_X1 i_0_1_129 (.ZN (n_0_228), .A1 (slo__n453), .A2 (n_0_1_122), .B1 (hfn_ipo_n25), .B2 (n_0_1_121));
INV_X1 i_0_1_128 (.ZN (n_0_1_120), .A (\Res_imm[42] ));
INV_X1 i_0_1_127 (.ZN (n_0_1_119), .A (n_0_41));
OAI22_X1 i_0_1_126 (.ZN (n_0_227), .A1 (slo__n453), .A2 (n_0_1_120), .B1 (hfn_ipo_n25), .B2 (n_0_1_119));
INV_X1 i_0_1_125 (.ZN (n_0_1_118), .A (\Res_imm[41] ));
INV_X1 i_0_1_124 (.ZN (n_0_1_117), .A (n_0_40));
OAI22_X1 i_0_1_123 (.ZN (n_0_226), .A1 (slo__n453), .A2 (n_0_1_118), .B1 (hfn_ipo_n25), .B2 (n_0_1_117));
INV_X1 i_0_1_122 (.ZN (n_0_1_116), .A (\Res_imm[40] ));
INV_X1 i_0_1_121 (.ZN (n_0_1_115), .A (n_0_39));
OAI22_X1 i_0_1_120 (.ZN (n_0_224), .A1 (slo__n453), .A2 (n_0_1_116), .B1 (hfn_ipo_n25), .B2 (n_0_1_115));
INV_X1 i_0_1_119 (.ZN (n_0_1_114), .A (n_0_38));
NAND2_X2 i_0_1_118 (.ZN (n_0_1_113), .A1 (opt_ipo_n1555), .A2 (\Res_imm[39] ));
OAI21_X1 i_0_1_117 (.ZN (n_0_223), .A (n_0_1_113), .B1 (n_0_1_114), .B2 (hfn_ipo_n25));
INV_X1 i_0_1_116 (.ZN (n_0_1_112), .A (\Res_imm[37] ));
INV_X1 i_0_1_115 (.ZN (n_0_1_111), .A (n_0_36));
OAI22_X1 i_0_1_114 (.ZN (n_0_221), .A1 (slo__n453), .A2 (n_0_1_112), .B1 (hfn_ipo_n25), .B2 (n_0_1_111));
INV_X1 i_0_1_113 (.ZN (n_0_1_110), .A (\Res_imm[36] ));
INV_X1 i_0_1_112 (.ZN (n_0_1_109), .A (n_0_35));
OAI22_X1 i_0_1_111 (.ZN (n_0_220), .A1 (slo__n453), .A2 (n_0_1_110), .B1 (hfn_ipo_n25), .B2 (n_0_1_109));
INV_X1 i_0_1_110 (.ZN (n_0_1_108), .A (\Res_imm[35] ));
INV_X1 i_0_1_109 (.ZN (n_0_1_107), .A (n_0_34));
OAI22_X1 i_0_1_108 (.ZN (n_0_219), .A1 (slo__n453), .A2 (n_0_1_108), .B1 (hfn_ipo_n25), .B2 (n_0_1_107));
INV_X1 i_0_1_107 (.ZN (n_0_1_106), .A (\Res_imm[34] ));
INV_X1 i_0_1_106 (.ZN (n_0_1_105), .A (n_0_33));
OAI22_X1 i_0_1_105 (.ZN (n_0_218), .A1 (slo__n453), .A2 (n_0_1_106), .B1 (hfn_ipo_n25), .B2 (n_0_1_105));
INV_X1 i_0_1_104 (.ZN (n_0_1_104), .A (\Res_imm[33] ));
INV_X1 i_0_1_103 (.ZN (n_0_1_103), .A (n_0_32));
OAI22_X1 i_0_1_102 (.ZN (n_0_217), .A1 (slo__n453), .A2 (n_0_1_104), .B1 (hfn_ipo_n25), .B2 (n_0_1_103));
INV_X1 i_0_1_101 (.ZN (n_0_1_102), .A (\Res_imm[32] ));
INV_X1 i_0_1_100 (.ZN (n_0_1_101), .A (n_0_31));
OAI22_X1 i_0_1_99 (.ZN (n_0_216), .A1 (slo__n453), .A2 (n_0_1_102), .B1 (hfn_ipo_n25), .B2 (n_0_1_101));
INV_X1 i_0_1_98 (.ZN (n_0_1_100), .A (\Res_imm[31] ));
INV_X1 i_0_1_97 (.ZN (n_0_1_99), .A (n_0_30));
OAI22_X1 i_0_1_96 (.ZN (n_0_215), .A1 (slo__n453), .A2 (n_0_1_100), .B1 (hfn_ipo_n25), .B2 (n_0_1_99));
INV_X1 i_0_1_95 (.ZN (n_0_1_98), .A (\Res_imm[30] ));
INV_X1 i_0_1_94 (.ZN (n_0_1_97), .A (n_0_29));
OAI22_X1 i_0_1_93 (.ZN (n_0_214), .A1 (slo__n453), .A2 (n_0_1_98), .B1 (hfn_ipo_n25), .B2 (n_0_1_97));
INV_X1 i_0_1_92 (.ZN (n_0_1_96), .A (\Res_imm[29] ));
INV_X1 i_0_1_91 (.ZN (n_0_1_95), .A (n_0_28));
OAI22_X1 i_0_1_90 (.ZN (n_0_213), .A1 (slo__n453), .A2 (n_0_1_96), .B1 (hfn_ipo_n25), .B2 (n_0_1_95));
INV_X1 i_0_1_89 (.ZN (n_0_1_94), .A (\Res_imm[28] ));
INV_X1 i_0_1_88 (.ZN (n_0_1_93), .A (n_0_27));
OAI22_X1 i_0_1_87 (.ZN (n_0_212), .A1 (slo__n453), .A2 (n_0_1_94), .B1 (hfn_ipo_n24), .B2 (n_0_1_93));
INV_X1 i_0_1_86 (.ZN (n_0_1_92), .A (\Res_imm[27] ));
INV_X1 i_0_1_85 (.ZN (n_0_1_91), .A (n_0_26));
OAI22_X1 i_0_1_84 (.ZN (n_0_211), .A1 (slo__n453), .A2 (n_0_1_92), .B1 (hfn_ipo_n24), .B2 (n_0_1_91));
INV_X1 i_0_1_83 (.ZN (n_0_1_88), .A (\Res_imm[26] ));
INV_X1 i_0_1_82 (.ZN (n_0_1_87), .A (n_0_25));
OAI22_X1 i_0_1_81 (.ZN (n_0_210), .A1 (slo__n453), .A2 (n_0_1_88), .B1 (hfn_ipo_n24), .B2 (n_0_1_87));
INV_X1 i_0_1_80 (.ZN (n_0_1_86), .A (\Res_imm[25] ));
INV_X1 i_0_1_79 (.ZN (n_0_1_85), .A (n_0_24));
OAI22_X1 i_0_1_78 (.ZN (n_0_209), .A1 (slo__n453), .A2 (n_0_1_86), .B1 (hfn_ipo_n24), .B2 (n_0_1_85));
INV_X1 i_0_1_77 (.ZN (n_0_1_84), .A (\Res_imm[24] ));
INV_X1 i_0_1_76 (.ZN (n_0_1_83), .A (n_0_23));
OAI22_X1 i_0_1_75 (.ZN (n_0_208), .A1 (slo__n453), .A2 (n_0_1_84), .B1 (hfn_ipo_n24), .B2 (n_0_1_83));
INV_X1 i_0_1_74 (.ZN (n_0_1_82), .A (\Res_imm[23] ));
INV_X1 i_0_1_73 (.ZN (n_0_1_81), .A (n_0_22));
OAI22_X1 i_0_1_72 (.ZN (n_0_207), .A1 (slo__n453), .A2 (n_0_1_82), .B1 (hfn_ipo_n24), .B2 (n_0_1_81));
INV_X1 i_0_1_71 (.ZN (n_0_1_80), .A (\Res_imm[22] ));
INV_X1 i_0_1_70 (.ZN (n_0_1_79), .A (n_0_21));
OAI22_X1 i_0_1_69 (.ZN (n_0_206), .A1 (slo__n453), .A2 (n_0_1_80), .B1 (hfn_ipo_n24), .B2 (n_0_1_79));
INV_X1 i_0_1_68 (.ZN (n_0_1_78), .A (\Res_imm[21] ));
INV_X1 i_0_1_67 (.ZN (n_0_1_77), .A (n_0_20));
OAI22_X1 i_0_1_66 (.ZN (n_0_205), .A1 (opt_ipo_n1524), .A2 (n_0_1_78), .B1 (hfn_ipo_n24), .B2 (n_0_1_77));
INV_X1 i_0_1_65 (.ZN (n_0_1_72), .A (\Res_imm[20] ));
INV_X1 i_0_1_64 (.ZN (n_0_1_67), .A (n_0_19));
OAI22_X1 i_0_1_63 (.ZN (n_0_204), .A1 (slo__n453), .A2 (n_0_1_72), .B1 (hfn_ipo_n24), .B2 (n_0_1_67));
INV_X1 i_0_1_62 (.ZN (n_0_1_66), .A (\Res_imm[19] ));
INV_X1 i_0_1_61 (.ZN (n_0_1_65), .A (n_0_18));
OAI22_X1 i_0_1_60 (.ZN (n_0_203), .A1 (slo__n453), .A2 (n_0_1_66), .B1 (hfn_ipo_n24), .B2 (n_0_1_65));
INV_X1 i_0_1_59 (.ZN (n_0_1_64), .A (\Res_imm[18] ));
INV_X1 i_0_1_58 (.ZN (n_0_1_63), .A (n_0_17));
OAI22_X1 i_0_1_57 (.ZN (n_0_202), .A1 (slo__n453), .A2 (n_0_1_64), .B1 (hfn_ipo_n24), .B2 (n_0_1_63));
INV_X1 i_0_1_56 (.ZN (n_0_1_62), .A (\Res_imm[17] ));
INV_X1 i_0_1_55 (.ZN (n_0_1_61), .A (n_0_16));
OAI22_X1 i_0_1_54 (.ZN (n_0_201), .A1 (slo__n453), .A2 (n_0_1_62), .B1 (hfn_ipo_n24), .B2 (n_0_1_61));
INV_X1 i_0_1_53 (.ZN (n_0_1_60), .A (\Res_imm[16] ));
INV_X1 i_0_1_52 (.ZN (n_0_1_59), .A (n_0_15));
OAI22_X1 i_0_1_51 (.ZN (n_0_200), .A1 (slo__n453), .A2 (n_0_1_60), .B1 (hfn_ipo_n24), .B2 (n_0_1_59));
INV_X1 i_0_1_50 (.ZN (n_0_1_58), .A (\Res_imm[15] ));
INV_X1 i_0_1_49 (.ZN (n_0_1_57), .A (n_0_14));
OAI22_X2 i_0_1_48 (.ZN (n_0_199), .A1 (slo__n453), .A2 (n_0_1_58), .B1 (hfn_ipo_n24), .B2 (n_0_1_57));
INV_X1 i_0_1_47 (.ZN (n_0_1_56), .A (\Res_imm[14] ));
INV_X1 i_0_1_46 (.ZN (n_0_1_55), .A (n_0_13));
OAI22_X2 i_0_1_45 (.ZN (n_0_198), .A1 (slo__n453), .A2 (n_0_1_56), .B1 (CLOCK_slo__n2626), .B2 (n_0_1_55));
INV_X1 i_0_1_44 (.ZN (n_0_1_54), .A (\Res_imm[13] ));
INV_X1 i_0_1_43 (.ZN (n_0_1_53), .A (n_0_12));
OAI22_X1 i_0_1_42 (.ZN (n_0_197), .A1 (slo__n453), .A2 (n_0_1_54), .B1 (CLOCK_slo__n2626), .B2 (n_0_1_53));
INV_X1 i_0_1_41 (.ZN (n_0_1_52), .A (\Res_imm[12] ));
INV_X1 i_0_1_40 (.ZN (n_0_1_51), .A (n_0_11));
OAI22_X1 i_0_1_39 (.ZN (n_0_196), .A1 (slo__n453), .A2 (n_0_1_52), .B1 (hfn_ipo_n24), .B2 (n_0_1_51));
INV_X1 i_0_1_38 (.ZN (n_0_1_50), .A (\Res_imm[11] ));
INV_X1 i_0_1_37 (.ZN (n_0_1_49), .A (n_0_10));
OAI22_X1 i_0_1_36 (.ZN (n_0_195), .A1 (slo__n453), .A2 (n_0_1_50), .B1 (hfn_ipo_n24), .B2 (n_0_1_49));
INV_X1 i_0_1_35 (.ZN (n_0_1_48), .A (\Res_imm[10] ));
INV_X1 i_0_1_34 (.ZN (n_0_1_47), .A (n_0_9));
OAI22_X2 i_0_1_33 (.ZN (n_0_194), .A1 (slo__n453), .A2 (n_0_1_48), .B1 (hfn_ipo_n24), .B2 (n_0_1_47));
INV_X1 i_0_1_32 (.ZN (n_0_1_46), .A (\Res_imm[9] ));
INV_X1 i_0_1_31 (.ZN (n_0_1_45), .A (n_0_8));
OAI22_X1 i_0_1_30 (.ZN (n_0_193), .A1 (slo__n453), .A2 (n_0_1_46), .B1 (hfn_ipo_n24), .B2 (n_0_1_45));
INV_X1 i_0_1_29 (.ZN (n_0_1_44), .A (\secondStage_Res[8] ));
INV_X1 i_0_1_28 (.ZN (n_0_1_43), .A (n_0_7));
OAI22_X1 i_0_1_27 (.ZN (n_0_192), .A1 (slo__n453), .A2 (n_0_1_44), .B1 (hfn_ipo_n24), .B2 (n_0_1_43));
INV_X1 i_0_1_26 (.ZN (n_0_1_42), .A (\secondStage_Res[7] ));
INV_X1 i_0_1_25 (.ZN (n_0_1_41), .A (n_0_6));
OAI22_X2 i_0_1_24 (.ZN (n_0_191), .A1 (slo__n453), .A2 (n_0_1_42), .B1 (CLOCK_slo__n2626), .B2 (n_0_1_41));
INV_X1 i_0_1_23 (.ZN (n_0_1_40), .A (\secondStage_Res[6] ));
INV_X1 i_0_1_21 (.ZN (n_0_1_39), .A (n_0_5));
OAI22_X2 i_0_1_20 (.ZN (n_0_190), .A1 (slo__n453), .A2 (n_0_1_40), .B1 (hfn_ipo_n24), .B2 (n_0_1_39));
INV_X1 i_0_1_19 (.ZN (n_0_1_38), .A (\secondStage_Res[5] ));
INV_X1 i_0_1_18 (.ZN (n_0_1_37), .A (n_0_4));
OAI22_X1 i_0_1_17 (.ZN (n_0_189), .A1 (slo__n453), .A2 (n_0_1_38), .B1 (hfn_ipo_n24), .B2 (n_0_1_37));
INV_X1 i_0_1_16 (.ZN (n_0_1_36), .A (\secondStage_Res[4] ));
INV_X1 i_0_1_14 (.ZN (n_0_1_35), .A (n_0_3));
OAI22_X1 i_0_1_13 (.ZN (n_0_188), .A1 (slo__n453), .A2 (n_0_1_36), .B1 (CLOCK_slo__n2626), .B2 (n_0_1_35));
INV_X1 i_0_1_12 (.ZN (n_0_1_34), .A (\secondStage_Res[3] ));
INV_X1 i_0_1_11 (.ZN (n_0_1_33), .A (n_0_2));
OAI22_X1 i_0_1_10 (.ZN (n_0_187), .A1 (CLOCK_slo__n2403), .A2 (n_0_1_34), .B1 (CLOCK_slo__n2449), .B2 (n_0_1_33));
INV_X1 i_0_1_9 (.ZN (n_0_1_32), .A (\secondStage_Res[2] ));
INV_X1 i_0_1_8 (.ZN (n_0_1_31), .A (n_0_1));
OAI22_X1 i_0_1_7 (.ZN (n_0_186), .A1 (slo__n453), .A2 (n_0_1_32), .B1 (hfn_ipo_n24), .B2 (n_0_1_31));
INV_X1 i_0_1_6 (.ZN (n_0_1_30), .A (\secondStage_Res[1] ));
INV_X1 i_0_1_5 (.ZN (n_0_1_29), .A (n_0_0));
OAI22_X1 i_0_1_4 (.ZN (n_0_185), .A1 (slo__n453), .A2 (n_0_1_30), .B1 (hfn_ipo_n24), .B2 (n_0_1_29));
MUX2_X2 i_0_1_2 (.Z (\B_imm[28] ), .A (n_0_65), .B (n_0_180), .S (drc_ipo_n27));
NAND2_X1 CLOCK_sgo__sro_c2230 (.ZN (CLOCK_sgo__sro_n1963), .A1 (CLOCK_sgo__sro_n1964), .A2 (CLOCK_sgo__sro_n1965));
MUX2_X2 i_0_1_278 (.Z (\A_imm[30] ), .A (n_0_93), .B (n_0_152), .S (drc_ipo_n26));
MUX2_X2 i_0_1_277 (.Z (\A_imm[29] ), .A (n_0_94), .B (n_0_151), .S (drc_ipo_n26));
MUX2_X2 i_0_1_276 (.Z (\A_imm[28] ), .A (n_0_95), .B (n_0_150), .S (drc_ipo_n26));
CLKBUF_X1 CLOCK_slo___L1_c1_c3657 (.Z (\Res_imm[59] ), .A (CLOCK_slo___n3239));
CLKBUF_X1 CLOCK_slh__c3966 (.Z (CLOCK_slh__n3499), .A (enable));
INV_X1 slo__sro_c715 (.ZN (slo__sro_n551), .A (drc_ipo_n26));
MUX2_X1 i_0_1_252 (.Z (\A_imm[4] ), .A (n_0_119), .B (opt_ipo_n1598), .S (drc_ipo_n26));
MUX2_X1 i_0_1_251 (.Z (\A_imm[3] ), .A (n_0_120), .B (n_0_125), .S (drc_ipo_n26));
MUX2_X1 i_0_1_250 (.Z (\A_imm[2] ), .A (n_0_121), .B (n_0_124), .S (drc_ipo_n26));
MUX2_X1 i_0_1_249 (.Z (\A_imm[1] ), .A (n_0_122), .B (n_0_123), .S (drc_ipo_n26));
AND2_X1 i_0_1_248 (.ZN (\B_imm[31] ), .A1 (drc_ipo_n27), .A2 (n_0_183));
MUX2_X1 i_0_1_247 (.Z (\B_imm[30] ), .A (n_0_63), .B (n_0_182), .S (drc_ipo_n27));
MUX2_X2 i_0_1_246 (.Z (\B_imm[29] ), .A (n_0_64), .B (n_0_181), .S (drc_ipo_n27));
MUX2_X2 i_0_1_244 (.Z (\B_imm[27] ), .A (n_0_66), .B (n_0_179), .S (drc_ipo_n27));
MUX2_X1 i_0_1_243 (.Z (\B_imm[26] ), .A (n_0_67), .B (n_0_178), .S (drc_ipo_n27));
INV_X1 CLOCK_slo__sro_c3217 (.ZN (CLOCK_slo__sro_n2844), .A (drc_ipo_n27));
MUX2_X1 i_0_1_240 (.Z (\B_imm[23] ), .A (n_0_70), .B (n_0_175), .S (drc_ipo_n27));
NOR2_X1 slo__sro_c697 (.ZN (slo__sro_n535), .A1 (\Res_imm[29] ), .A2 (\Res_imm[24] ));
INV_X1 slo__sro_c1401 (.ZN (slo__sro_n1189), .A (drc_ipo_n27));
MUX2_X1 i_0_1_237 (.Z (\B_imm[20] ), .A (n_0_73), .B (n_0_172), .S (drc_ipo_n27));
MUX2_X2 i_0_1_236 (.Z (\B_imm[19] ), .A (n_0_74), .B (n_0_171), .S (drc_ipo_n27));
MUX2_X2 i_0_1_235 (.Z (\B_imm[18] ), .A (n_0_75), .B (n_0_170), .S (drc_ipo_n27));
MUX2_X1 i_0_1_234 (.Z (\B_imm[17] ), .A (n_0_76), .B (n_0_169), .S (drc_ipo_n27));
BUF_X8 CLOCK_slo__c3142 (.Z (\B_imm[1] ), .A (CLOCK_slo__n2760));
NAND2_X1 CLOCK_slo__sro_c3219 (.ZN (CLOCK_slo__sro_n2842), .A1 (n_0_87), .A2 (CLOCK_slo__sro_n2844));
MUX2_X1 i_0_1_231 (.Z (\B_imm[14] ), .A (n_0_79), .B (n_0_166), .S (drc_ipo_n27));
MUX2_X2 i_0_1_230 (.Z (\B_imm[13] ), .A (n_0_80), .B (n_0_165), .S (drc_ipo_n27));
MUX2_X2 i_0_1_229 (.Z (\B_imm[12] ), .A (n_0_81), .B (n_0_164), .S (drc_ipo_n27));
MUX2_X2 i_0_1_228 (.Z (\B_imm[11] ), .A (n_0_82), .B (n_0_163), .S (drc_ipo_n27));
MUX2_X1 i_0_1_225 (.Z (\B_imm[8] ), .A (n_0_85), .B (n_0_160), .S (drc_ipo_n27));
MUX2_X1 i_0_1_222 (.Z (\B_imm[5] ), .A (n_0_88), .B (n_0_157), .S (drc_ipo_n27));
MUX2_X1 i_0_1_221 (.Z (\B_imm[4] ), .A (n_0_89), .B (n_0_156), .S (drc_ipo_n27));
MUX2_X2 i_0_1_220 (.Z (\B_imm[3] ), .A (n_0_90), .B (n_0_155), .S (drc_ipo_n27));
MUX2_X1 i_0_1_219 (.Z (\B_imm[2] ), .A (n_0_91), .B (n_0_154), .S (drc_ipo_n27));
MUX2_X1 i_0_1_218 (.Z (CLOCK_slo__n2760), .A (n_0_92), .B (n_0_153), .S (drc_ipo_n27));
AND2_X1 i_0_1_216 (.ZN (n_0_314), .A1 (hfn_ipo_n22), .A2 (B[31]));
AND2_X1 i_0_1_215 (.ZN (n_0_313), .A1 (hfn_ipo_n23), .A2 (B[30]));
AND2_X1 i_0_1_214 (.ZN (n_0_312), .A1 (hfn_ipo_n23), .A2 (B[29]));
AND2_X1 i_0_1_213 (.ZN (n_0_311), .A1 (hfn_ipo_n23), .A2 (B[28]));
AND2_X1 i_0_1_212 (.ZN (n_0_310), .A1 (hfn_ipo_n23), .A2 (B[27]));
AND2_X1 i_0_1_211 (.ZN (n_0_309), .A1 (hfn_ipo_n23), .A2 (B[26]));
AND2_X1 i_0_1_210 (.ZN (n_0_308), .A1 (hfn_ipo_n23), .A2 (B[25]));
AND2_X1 i_0_1_209 (.ZN (n_0_307), .A1 (hfn_ipo_n23), .A2 (B[24]));
AND2_X1 i_0_1_208 (.ZN (n_0_306), .A1 (hfn_ipo_n23), .A2 (B[23]));
AND2_X1 i_0_1_207 (.ZN (n_0_305), .A1 (hfn_ipo_n23), .A2 (B[22]));
AND2_X1 i_0_1_206 (.ZN (n_0_304), .A1 (hfn_ipo_n23), .A2 (B[21]));
AND2_X1 i_0_1_205 (.ZN (n_0_303), .A1 (hfn_ipo_n23), .A2 (B[20]));
AND2_X1 i_0_1_204 (.ZN (n_0_302), .A1 (hfn_ipo_n23), .A2 (B[19]));
AND2_X1 i_0_1_203 (.ZN (n_0_301), .A1 (hfn_ipo_n23), .A2 (B[18]));
AND2_X1 i_0_1_202 (.ZN (n_0_300), .A1 (hfn_ipo_n23), .A2 (B[17]));
AND2_X1 i_0_1_201 (.ZN (n_0_299), .A1 (hfn_ipo_n23), .A2 (B[16]));
AND2_X1 i_0_1_200 (.ZN (n_0_298), .A1 (hfn_ipo_n22), .A2 (B[15]));
AND2_X1 i_0_1_199 (.ZN (n_0_297), .A1 (hfn_ipo_n22), .A2 (B[14]));
AND2_X1 i_0_1_198 (.ZN (n_0_296), .A1 (hfn_ipo_n22), .A2 (B[13]));
AND2_X1 i_0_1_197 (.ZN (n_0_295), .A1 (hfn_ipo_n22), .A2 (B[12]));
AND2_X1 i_0_1_196 (.ZN (n_0_294), .A1 (hfn_ipo_n22), .A2 (B[11]));
AND2_X1 i_0_1_195 (.ZN (n_0_293), .A1 (hfn_ipo_n22), .A2 (B[10]));
AND2_X1 i_0_1_194 (.ZN (n_0_292), .A1 (hfn_ipo_n22), .A2 (B[9]));
AND2_X1 i_0_1_193 (.ZN (n_0_291), .A1 (hfn_ipo_n22), .A2 (B[8]));
AND2_X1 i_0_1_192 (.ZN (n_0_290), .A1 (hfn_ipo_n23), .A2 (B[7]));
AND2_X1 i_0_1_191 (.ZN (n_0_289), .A1 (hfn_ipo_n23), .A2 (B[6]));
AND2_X1 i_0_1_190 (.ZN (n_0_288), .A1 (hfn_ipo_n22), .A2 (B[5]));
AND2_X1 i_0_1_189 (.ZN (n_0_287), .A1 (hfn_ipo_n22), .A2 (B[4]));
AND2_X1 i_0_1_188 (.ZN (n_0_286), .A1 (hfn_ipo_n22), .A2 (B[3]));
AND2_X1 i_0_1_187 (.ZN (n_0_285), .A1 (hfn_ipo_n22), .A2 (B[2]));
AND2_X1 i_0_1_186 (.ZN (n_0_284), .A1 (hfn_ipo_n22), .A2 (B[1]));
AND2_X1 i_0_1_185 (.ZN (n_0_283), .A1 (hfn_ipo_n22), .A2 (B[0]));
NOR2_X1 i_0_1_3 (.ZN (n_0_281), .A1 (CLOCK_opt_ipo_n1683), .A2 (reset));
AND2_X1 i_0_1_181 (.ZN (n_0_280), .A1 (hfn_ipo_n23), .A2 (A[30]));
AND2_X1 i_0_1_180 (.ZN (n_0_279), .A1 (hfn_ipo_n22), .A2 (A[29]));
AND2_X1 i_0_1_179 (.ZN (n_0_278), .A1 (hfn_ipo_n22), .A2 (A[28]));
AND2_X1 i_0_1_178 (.ZN (n_0_277), .A1 (hfn_ipo_n23), .A2 (A[27]));
AND2_X1 i_0_1_177 (.ZN (n_0_276), .A1 (hfn_ipo_n23), .A2 (A[26]));
AND2_X1 i_0_1_176 (.ZN (n_0_275), .A1 (hfn_ipo_n23), .A2 (A[25]));
AND2_X1 i_0_1_175 (.ZN (n_0_274), .A1 (hfn_ipo_n22), .A2 (A[24]));
AND2_X1 i_0_1_174 (.ZN (n_0_273), .A1 (hfn_ipo_n22), .A2 (A[23]));
AND2_X1 i_0_1_173 (.ZN (n_0_272), .A1 (hfn_ipo_n22), .A2 (A[22]));
AND2_X1 i_0_1_172 (.ZN (n_0_271), .A1 (hfn_ipo_n22), .A2 (A[21]));
AND2_X1 i_0_1_171 (.ZN (n_0_270), .A1 (hfn_ipo_n22), .A2 (A[20]));
AND2_X1 i_0_1_170 (.ZN (n_0_269), .A1 (hfn_ipo_n22), .A2 (A[19]));
AND2_X1 i_0_1_169 (.ZN (n_0_268), .A1 (hfn_ipo_n22), .A2 (A[18]));
AND2_X1 i_0_1_168 (.ZN (n_0_267), .A1 (hfn_ipo_n22), .A2 (A[17]));
AND2_X1 i_0_1_167 (.ZN (n_0_266), .A1 (hfn_ipo_n22), .A2 (A[16]));
AND2_X1 i_0_1_166 (.ZN (n_0_265), .A1 (hfn_ipo_n22), .A2 (A[15]));
AND2_X1 i_0_1_165 (.ZN (n_0_264), .A1 (hfn_ipo_n22), .A2 (A[14]));
AND2_X1 i_0_1_164 (.ZN (n_0_263), .A1 (hfn_ipo_n22), .A2 (A[13]));
AND2_X1 i_0_1_163 (.ZN (n_0_262), .A1 (hfn_ipo_n22), .A2 (A[12]));
AND2_X1 i_0_1_162 (.ZN (n_0_261), .A1 (hfn_ipo_n22), .A2 (A[11]));
AND2_X1 i_0_1_161 (.ZN (n_0_260), .A1 (hfn_ipo_n22), .A2 (A[10]));
AND2_X1 i_0_1_160 (.ZN (n_0_259), .A1 (hfn_ipo_n22), .A2 (A[9]));
AND2_X4 i_0_1_159 (.ZN (n_0_258), .A1 (hfn_ipo_n22), .A2 (A[8]));
AND2_X1 i_0_1_158 (.ZN (n_0_257), .A1 (hfn_ipo_n23), .A2 (A[7]));
AND2_X1 i_0_1_157 (.ZN (n_0_255), .A1 (hfn_ipo_n23), .A2 (A[6]));
AND2_X1 i_0_1_156 (.ZN (n_0_254), .A1 (hfn_ipo_n23), .A2 (A[5]));
AND2_X1 i_0_1_155 (.ZN (n_0_253), .A1 (hfn_ipo_n23), .A2 (A[4]));
AND2_X1 i_0_1_154 (.ZN (n_0_252), .A1 (hfn_ipo_n23), .A2 (A[3]));
AND2_X1 i_0_1_153 (.ZN (n_0_251), .A1 (hfn_ipo_n23), .A2 (A[2]));
AND2_X1 i_0_1_152 (.ZN (n_0_250), .A1 (hfn_ipo_n23), .A2 (A[1]));
AND2_X4 i_0_1_151 (.ZN (n_0_249), .A1 (hfn_ipo_n23), .A2 (A[0]));
AND2_X1 i_0_1_0 (.ZN (n_0_184), .A1 (hfn_ipo_n23), .A2 (n_0_316));
datapath__0_131 i_0_13 (.p_0 ({n_0_183, n_0_182, n_0_181, n_0_180, n_0_179, n_0_178, 
    n_0_177, n_0_176, n_0_175, n_0_174, n_0_173, n_0_172, n_0_171, n_0_170, n_0_169, 
    n_0_168, n_0_167, n_0_166, n_0_165, n_0_164, n_0_163, n_0_162, n_0_161, n_0_160, 
    n_0_159, n_0_158, n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, uc_2161}), .B_in ({
    drc_ipo_n27, n_0_63, n_0_64, n_0_65, n_0_66, n_0_67, n_0_68, n_0_69, n_0_70, 
    n_0_71, n_0_72, n_0_73, n_0_74, n_0_75, n_0_76, n_0_77, n_0_78, n_0_79, n_0_80, 
    n_0_81, n_0_82, n_0_83, n_0_84, n_0_85, opt_ipo_n1541, n_0_87, n_0_88, n_0_89, 
    n_0_90, n_0_91, n_0_92, slo__n345}), .opt_ipoPP_0 (n_0_72), .opt_ipoPP_2 (opt_ipo_n1540));
datapath__0_129 i_0_11 (.p_0 ({uc_2159, n_0_152, n_0_151, n_0_150, n_0_149, n_0_148, 
    n_0_147, n_0_146, n_0_145, n_0_144, n_0_143, n_0_142, n_0_141, n_0_140, n_0_139, 
    n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, 
    n_0_129, n_0_128, n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, uc_2160}), .A_in ({
    uc_2158, n_0_93, n_0_94, n_0_95, n_0_96, n_0_97, n_0_98, n_0_99, n_0_100, n_0_101, 
    n_0_102, n_0_103, n_0_104, n_0_105, n_0_106, n_0_107, n_0_108, n_0_109, n_0_110, 
    n_0_111, n_0_112, opt_ipo_n1364, n_0_114, n_0_115, n_0_116, n_0_117, n_0_118, 
    n_0_119, n_0_120, n_0_121, n_0_122, n_0_256}), .opt_ipoPP_2 (opt_ipo_n1363));
DLH_X2 \A_in_reg[0]  (.Q (n_0_256), .D (n_0_249), .G (CTS_n1730));
DLH_X2 \A_in_reg[1]  (.Q (n_0_122), .D (n_0_250), .G (CTS_n1730));
DLH_X2 \A_in_reg[2]  (.Q (n_0_121), .D (n_0_251), .G (CTS_n1730));
DLH_X2 \A_in_reg[3]  (.Q (n_0_120), .D (n_0_252), .G (CTS_n1730));
DLH_X2 \A_in_reg[4]  (.Q (n_0_119), .D (n_0_253), .G (CTS_n1730));
DLH_X1 \A_in_reg[5]  (.Q (n_0_118), .D (n_0_254), .G (CTS_n1730));
DLH_X2 \A_in_reg[6]  (.Q (n_0_117), .D (n_0_255), .G (CTS_n1730));
DLH_X2 \A_in_reg[7]  (.Q (n_0_116), .D (n_0_257), .G (CTS_n1730));
DLH_X1 \A_in_reg[8]  (.Q (n_0_115), .D (n_0_258), .G (CTS_n1730));
DLH_X2 \A_in_reg[9]  (.Q (n_0_114), .D (n_0_259), .G (CTS_n1730));
DLH_X1 \A_in_reg[10]  (.Q (n_0_113), .D (n_0_260), .G (CTS_n1730));
DLH_X1 \A_in_reg[11]  (.Q (n_0_112), .D (n_0_261), .G (CTS_n1730));
DLH_X1 \A_in_reg[12]  (.Q (n_0_111), .D (n_0_262), .G (CTS_n1730));
DLH_X1 \A_in_reg[13]  (.Q (n_0_110), .D (n_0_263), .G (CTS_n1730));
DLH_X1 \A_in_reg[14]  (.Q (n_0_109), .D (n_0_264), .G (CTS_n1730));
DLH_X2 \A_in_reg[15]  (.Q (n_0_108), .D (n_0_265), .G (CTS_n1730));
DLH_X2 \A_in_reg[16]  (.Q (n_0_107), .D (n_0_266), .G (CTS_n1730));
DLH_X1 \A_in_reg[17]  (.Q (n_0_106), .D (n_0_267), .G (CTS_n1730));
DLH_X2 \A_in_reg[18]  (.Q (n_0_105), .D (n_0_268), .G (CTS_n1730));
DLH_X1 \A_in_reg[19]  (.Q (n_0_104), .D (n_0_269), .G (CTS_n1730));
DLH_X1 \A_in_reg[20]  (.Q (n_0_103), .D (n_0_270), .G (CTS_n1730));
DLH_X2 \A_in_reg[21]  (.Q (n_0_102), .D (n_0_271), .G (CTS_n1730));
DLH_X1 \A_in_reg[22]  (.Q (n_0_101), .D (n_0_272), .G (CTS_n1730));
DLH_X1 \A_in_reg[23]  (.Q (n_0_100), .D (n_0_273), .G (CTS_n1730));
DLH_X2 \A_in_reg[24]  (.Q (n_0_99), .D (n_0_274), .G (CTS_n1730));
DLH_X1 \A_in_reg[25]  (.Q (n_0_98), .D (n_0_275), .G (CTS_n1730));
DLH_X1 \A_in_reg[26]  (.Q (n_0_97), .D (n_0_276), .G (CTS_n1730));
DLH_X1 \A_in_reg[27]  (.Q (n_0_96), .D (n_0_277), .G (CTS_n1730));
DLH_X1 \A_in_reg[28]  (.Q (n_0_95), .D (n_0_278), .G (CTS_n1730));
DLH_X1 \A_in_reg[29]  (.Q (n_0_94), .D (n_0_279), .G (CTS_n1730));
DLH_X1 \A_in_reg[30]  (.Q (n_0_93), .D (n_0_280), .G (CTS_n1730));
DLH_X1 \A_in_reg[31]  (.Q (A_in), .D (n_0_281), .G (CTS_n1730));
DLH_X1 \B_in_reg[0]  (.Q (slo__n345), .D (n_0_283), .G (CTS_n1730));
DLH_X2 \B_in_reg[1]  (.Q (n_0_92), .D (n_0_284), .G (CTS_n1730));
DLH_X2 \B_in_reg[2]  (.Q (n_0_91), .D (n_0_285), .G (CTS_n1730));
DLH_X2 \B_in_reg[3]  (.Q (n_0_90), .D (n_0_286), .G (CTS_n1730));
DLH_X2 \B_in_reg[4]  (.Q (n_0_89), .D (n_0_287), .G (CTS_n1730));
DLH_X1 \B_in_reg[5]  (.Q (n_0_88), .D (n_0_288), .G (CTS_n1730));
DLH_X1 \B_in_reg[6]  (.Q (n_0_87), .D (n_0_289), .G (CTS_n1730));
DLH_X1 \B_in_reg[7]  (.Q (n_0_86), .D (n_0_290), .G (CTS_n1730));
DLH_X1 \B_in_reg[8]  (.Q (n_0_85), .D (n_0_291), .G (CTS_n1730));
DLH_X1 \B_in_reg[9]  (.Q (n_0_84), .D (n_0_292), .G (CTS_n1730));
DLH_X1 \B_in_reg[10]  (.Q (n_0_83), .D (n_0_293), .G (CTS_n1730));
DLH_X1 \B_in_reg[11]  (.Q (n_0_82), .D (n_0_294), .G (CTS_n1730));
DLH_X2 \B_in_reg[12]  (.Q (n_0_81), .D (n_0_295), .G (CTS_n1730));
DLH_X2 \B_in_reg[13]  (.Q (n_0_80), .D (n_0_296), .G (CTS_n1730));
DLH_X1 \B_in_reg[14]  (.Q (n_0_79), .D (n_0_297), .G (CTS_n1730));
DLH_X1 \B_in_reg[15]  (.Q (n_0_78), .D (n_0_298), .G (CTS_n1730));
DLH_X1 \B_in_reg[16]  (.Q (n_0_77), .D (n_0_299), .G (CTS_n1730));
DLH_X1 \B_in_reg[17]  (.Q (n_0_76), .D (n_0_300), .G (CTS_n1730));
DLH_X1 \B_in_reg[18]  (.Q (n_0_75), .D (n_0_301), .G (CTS_n1730));
DLH_X1 \B_in_reg[19]  (.Q (n_0_74), .D (n_0_302), .G (CTS_n1730));
DLH_X1 \B_in_reg[20]  (.Q (n_0_73), .D (n_0_303), .G (CTS_n1730));
DLH_X2 \B_in_reg[21]  (.Q (n_0_72), .D (n_0_304), .G (CTS_n1730));
DLH_X1 \B_in_reg[22]  (.Q (n_0_71), .D (n_0_305), .G (CTS_n1730));
DLH_X1 \B_in_reg[23]  (.Q (n_0_70), .D (n_0_306), .G (CTS_n1730));
DLH_X1 \B_in_reg[24]  (.Q (n_0_69), .D (n_0_307), .G (CTS_n1730));
DLH_X1 \B_in_reg[25]  (.Q (n_0_68), .D (n_0_308), .G (CTS_n1730));
DLH_X1 \B_in_reg[26]  (.Q (n_0_67), .D (n_0_309), .G (CTS_n1730));
DLH_X1 \B_in_reg[27]  (.Q (n_0_66), .D (n_0_310), .G (CTS_n1730));
DLH_X1 \B_in_reg[28]  (.Q (n_0_65), .D (n_0_311), .G (CTS_n1730));
DLH_X1 \B_in_reg[29]  (.Q (n_0_64), .D (n_0_312), .G (CTS_n1730));
DLH_X1 \B_in_reg[30]  (.Q (n_0_63), .D (n_0_313), .G (CTS_n1730));
DLH_X1 \B_in_reg[31]  (.Q (B_in), .D (n_0_314), .G (CTS_n1730));
DLH_X1 \Res_reg[0]  (.Q (Res[0]), .D (n_0_184), .G (n_0_315));
DLH_X1 \Res_reg[1]  (.Q (Res[1]), .D (n_0_185), .G (n_0_315));
DLH_X1 \Res_reg[2]  (.Q (Res[2]), .D (n_0_186), .G (n_0_315));
DLH_X1 \Res_reg[3]  (.Q (Res[3]), .D (n_0_187), .G (n_0_315));
DLH_X1 \Res_reg[4]  (.Q (Res[4]), .D (n_0_188), .G (n_0_315));
DLH_X1 \Res_reg[5]  (.Q (Res[5]), .D (n_0_189), .G (n_0_315));
DLH_X1 \Res_reg[6]  (.Q (Res[6]), .D (n_0_190), .G (n_0_315));
DLH_X1 \Res_reg[7]  (.Q (Res[7]), .D (n_0_191), .G (n_0_315));
DLH_X1 \Res_reg[8]  (.Q (Res[8]), .D (n_0_192), .G (n_0_315));
DLH_X1 \Res_reg[9]  (.Q (Res[9]), .D (n_0_193), .G (n_0_315));
DLH_X1 \Res_reg[10]  (.Q (Res[10]), .D (n_0_194), .G (n_0_315));
DLH_X1 \Res_reg[11]  (.Q (Res[11]), .D (n_0_195), .G (n_0_315));
DLH_X1 \Res_reg[12]  (.Q (Res[12]), .D (n_0_196), .G (n_0_315));
DLH_X1 \Res_reg[13]  (.Q (Res[13]), .D (n_0_197), .G (n_0_315));
DLH_X1 \Res_reg[14]  (.Q (Res[14]), .D (n_0_198), .G (n_0_315));
DLH_X1 \Res_reg[15]  (.Q (Res[15]), .D (n_0_199), .G (n_0_315));
DLH_X1 \Res_reg[16]  (.Q (Res[16]), .D (n_0_200), .G (n_0_315));
DLH_X1 \Res_reg[17]  (.Q (Res[17]), .D (n_0_201), .G (n_0_315));
DLH_X1 \Res_reg[18]  (.Q (Res[18]), .D (n_0_202), .G (n_0_315));
DLH_X1 \Res_reg[19]  (.Q (Res[19]), .D (n_0_203), .G (n_0_315));
DLH_X1 \Res_reg[20]  (.Q (Res[20]), .D (n_0_204), .G (n_0_315));
DLH_X1 \Res_reg[21]  (.Q (Res[21]), .D (n_0_205), .G (n_0_315));
DLH_X1 \Res_reg[22]  (.Q (Res[22]), .D (n_0_206), .G (n_0_315));
DLH_X1 \Res_reg[23]  (.Q (Res[23]), .D (n_0_207), .G (n_0_315));
DLH_X1 \Res_reg[24]  (.Q (Res[24]), .D (n_0_208), .G (n_0_315));
DLH_X1 \Res_reg[25]  (.Q (Res[25]), .D (n_0_209), .G (n_0_315));
DLH_X1 \Res_reg[26]  (.Q (Res[26]), .D (n_0_210), .G (n_0_315));
DLH_X1 \Res_reg[27]  (.Q (Res[27]), .D (n_0_211), .G (n_0_315));
DLH_X1 \Res_reg[28]  (.Q (Res[28]), .D (n_0_212), .G (n_0_315));
DLH_X1 \Res_reg[29]  (.Q (Res[29]), .D (n_0_213), .G (n_0_315));
DLH_X1 \Res_reg[30]  (.Q (Res[30]), .D (n_0_214), .G (n_0_315));
DLH_X1 \Res_reg[31]  (.Q (Res[31]), .D (n_0_215), .G (n_0_315));
DLH_X1 \Res_reg[32]  (.Q (Res[32]), .D (n_0_216), .G (n_0_315));
DLH_X1 \Res_reg[33]  (.Q (Res[33]), .D (n_0_217), .G (n_0_315));
DLH_X1 \Res_reg[34]  (.Q (Res[34]), .D (n_0_218), .G (n_0_315));
DLH_X1 \Res_reg[35]  (.Q (Res[35]), .D (n_0_219), .G (n_0_315));
DLH_X1 \Res_reg[36]  (.Q (Res[36]), .D (n_0_220), .G (n_0_315));
DLH_X1 \Res_reg[37]  (.Q (Res[37]), .D (n_0_221), .G (n_0_315));
DLH_X1 \Res_reg[38]  (.Q (Res[38]), .D (n_0_222), .G (n_0_315));
DLH_X1 \Res_reg[39]  (.Q (Res[39]), .D (n_0_223), .G (n_0_315));
DLH_X1 \Res_reg[40]  (.Q (Res[40]), .D (n_0_224), .G (n_0_315));
DLH_X1 \Res_reg[41]  (.Q (Res[41]), .D (n_0_226), .G (n_0_315));
DLH_X1 \Res_reg[42]  (.Q (Res[42]), .D (n_0_227), .G (n_0_315));
DLH_X1 \Res_reg[43]  (.Q (Res[43]), .D (n_0_228), .G (n_0_315));
DLH_X1 \Res_reg[44]  (.Q (Res[44]), .D (n_0_229), .G (n_0_315));
DLH_X1 \Res_reg[45]  (.Q (Res[45]), .D (n_0_230), .G (n_0_315));
DLH_X1 \Res_reg[46]  (.Q (Res[46]), .D (n_0_231), .G (n_0_315));
DLH_X1 \Res_reg[47]  (.Q (Res[47]), .D (n_0_232), .G (n_0_315));
DLH_X1 \Res_reg[48]  (.Q (Res[48]), .D (n_0_233), .G (n_0_315));
DLH_X1 \Res_reg[49]  (.Q (Res[49]), .D (n_0_234), .G (n_0_315));
DLH_X1 \Res_reg[50]  (.Q (Res[50]), .D (n_0_235), .G (n_0_315));
DLH_X1 \Res_reg[51]  (.Q (Res[51]), .D (n_0_236), .G (n_0_315));
DLH_X1 \Res_reg[52]  (.Q (Res[52]), .D (n_0_237), .G (n_0_315));
DLH_X1 \Res_reg[53]  (.Q (Res[53]), .D (n_0_238), .G (n_0_315));
DLH_X1 \Res_reg[54]  (.Q (Res[54]), .D (n_0_239), .G (n_0_315));
DLH_X1 \Res_reg[55]  (.Q (Res[55]), .D (opt_ipo_n1547), .G (n_0_315));
DLH_X1 \Res_reg[56]  (.Q (Res[56]), .D (n_0_241), .G (n_0_315));
DLH_X1 \Res_reg[57]  (.Q (Res[57]), .D (n_0_242), .G (n_0_315));
DLH_X1 \Res_reg[58]  (.Q (Res[58]), .D (n_0_243), .G (n_0_315));
DLH_X2 \Res_reg[59]  (.Q (Res[59]), .D (n_0_244), .G (n_0_315));
DLH_X1 \Res_reg[60]  (.Q (Res[60]), .D (opt_ipo_n1569), .G (n_0_315));
DLH_X1 \Res_reg[61]  (.Q (Res[61]), .D (n_0_246), .G (n_0_315));
DLH_X1 \Res_reg[62]  (.Q (Res[62]), .D (n_0_247), .G (n_0_315));
DLH_X2 \Res_reg[63]  (.Q (sgo__n28), .D (n_0_248), .G (n_0_315));
datapath__0_119 i_0_0 (.p_0 ({n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, 
    n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, 
    n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, 
    n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, 
    n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
    n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, 
    n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, uc_2157}), .Res_imm ({\Res_imm[63] , opt_ipo_n1365, 
    CLOCK_opt_ipo_n1670, \Res_imm[60] , CLOCK_slo___n3239, \Res_imm[58] , \Res_imm[57] , 
    \Res_imm[56] , \Res_imm[55] , \Res_imm[54] , \Res_imm[53] , \Res_imm[52] , \Res_imm[51] , 
    \Res_imm[50] , \Res_imm[49] , \Res_imm[48] , \Res_imm[47] , \Res_imm[46] , \Res_imm[45] , 
    \Res_imm[44] , \Res_imm[43] , \Res_imm[42] , \Res_imm[41] , \Res_imm[40] , \Res_imm[39] , 
    \Res_imm[38] , \Res_imm[37] , \Res_imm[36] , \Res_imm[35] , \Res_imm[34] , \Res_imm[33] , 
    \Res_imm[32] , \Res_imm[31] , \Res_imm[30] , \Res_imm[29] , CLOCK_slo___n2653, 
    \Res_imm[27] , \Res_imm[26] , \Res_imm[25] , \Res_imm[24] , \Res_imm[23] , \Res_imm[22] , 
    \Res_imm[21] , \Res_imm[20] , \Res_imm[19] , \Res_imm[18] , \Res_imm[17] , \Res_imm[16] , 
    \Res_imm[15] , \Res_imm[14] , \Res_imm[13] , \Res_imm[12] , \Res_imm[11] , \Res_imm[10] , 
    \Res_imm[9] , \secondStage_Res[8] , \secondStage_Res[7] , \secondStage_Res[6] , 
    \secondStage_Res[5] , \secondStage_Res[4] , \secondStage_Res[3] , \secondStage_Res[2] , 
    \secondStage_Res[1] , n_0_316}), .opt_ipoPP_0 (opt_ipo_n1344), .opt_ipoPP_3 (opt_ipo_n1361));
addResWithCarry thirdStage (.Res_out ({\Res_imm[63] , \Res_imm[62] , \Res_imm[61] , 
    \Res_imm[60] , CLOCK_slo___n3239, \Res_imm[58] , \Res_imm[57] , \Res_imm[56] , 
    \Res_imm[55] , \Res_imm[54] , \Res_imm[53] , \Res_imm[52] , \Res_imm[51] , \Res_imm[50] , 
    \Res_imm[49] , \Res_imm[48] , \Res_imm[47] , \Res_imm[46] , \Res_imm[45] , \Res_imm[44] , 
    \Res_imm[43] , \Res_imm[42] , \Res_imm[41] , \Res_imm[40] , \Res_imm[39] , \Res_imm[38] , 
    \Res_imm[37] , \Res_imm[36] , \Res_imm[35] , \Res_imm[34] , \Res_imm[33] , \Res_imm[32] , 
    \Res_imm[31] , \Res_imm[30] , \Res_imm[29] , CLOCK_slo___n2653, \Res_imm[27] , 
    \Res_imm[26] , \Res_imm[25] , \Res_imm[24] , \Res_imm[23] , \Res_imm[22] , \Res_imm[21] , 
    \Res_imm[20] , \Res_imm[19] , \Res_imm[18] , \Res_imm[17] , \Res_imm[16] , \Res_imm[15] , 
    \Res_imm[14] , \Res_imm[13] , \Res_imm[12] , \Res_imm[11] , \Res_imm[10] , \Res_imm[9] , 
    uc_2127, uc_2128, uc_2129, uc_2130, uc_2131, uc_2132, uc_2133, uc_2134, uc_2135})
    , .Res_in ({uc_2136, uc_2137, \secondStage_Res[61] , \secondStage_Res[60] , \secondStage_Res[59] , 
    \secondStage_Res[58] , \secondStage_Res[57] , \secondStage_Res[56] , \secondStage_Res[55] , 
    \secondStage_Res[54] , \secondStage_Res[53] , \secondStage_Res[52] , \secondStage_Res[51] , 
    \secondStage_Res[50] , \secondStage_Res[49] , \secondStage_Res[48] , \secondStage_Res[47] , 
    \secondStage_Res[46] , \secondStage_Res[45] , \secondStage_Res[44] , \secondStage_Res[43] , 
    \secondStage_Res[42] , \secondStage_Res[41] , \secondStage_Res[40] , \secondStage_Res[39] , 
    \secondStage_Res[38] , \secondStage_Res[37] , \secondStage_Res[36] , \secondStage_Res[35] , 
    \secondStage_Res[34] , \secondStage_Res[33] , \secondStage_Res[32] , \secondStage_Res[31] , 
    \secondStage_Res[30] , \secondStage_Res[29] , \secondStage_Res[28] , \secondStage_Res[27] , 
    \secondStage_Res[26] , \secondStage_Res[25] , \secondStage_Res[24] , \secondStage_Res[23] , 
    \secondStage_Res[22] , \secondStage_Res[21] , \secondStage_Res[20] , \secondStage_Res[19] , 
    \secondStage_Res[18] , \secondStage_Res[17] , \secondStage_Res[16] , \secondStage_Res[15] , 
    \secondStage_Res[14] , \secondStage_Res[13] , \secondStage_Res[12] , \secondStage_Res[11] , 
    \secondStage_Res[10] , \secondStage_Res[9] , uc_2138, uc_2139, uc_2140, uc_2141, 
    uc_2142, uc_2143, uc_2144, uc_2145, uc_2146}), .carry_in ({uc_2147, \secondStage_carry[62] , 
    \secondStage_carry[61] , \secondStage_carry[60] , \secondStage_carry[59] , \secondStage_carry[58] , 
    \secondStage_carry[57] , \secondStage_carry[56] , \secondStage_carry[55] , \secondStage_carry[54] , 
    \secondStage_carry[53] , \secondStage_carry[52] , \secondStage_carry[51] , \secondStage_carry[50] , 
    \secondStage_carry[49] , \secondStage_carry[48] , \secondStage_carry[47] , \secondStage_carry[46] , 
    \secondStage_carry[45] , \secondStage_carry[44] , \secondStage_carry[43] , \secondStage_carry[42] , 
    \secondStage_carry[41] , \secondStage_carry[40] , \secondStage_carry[39] , \secondStage_carry[38] , 
    \secondStage_carry[37] , \secondStage_carry[36] , \secondStage_carry[35] , \secondStage_carry[34] , 
    \secondStage_carry[33] , \secondStage_carry[32] , \secondStage_carry[31] , \secondStage_carry[30] , 
    \secondStage_carry[29] , \secondStage_carry[28] , \secondStage_carry[27] , \secondStage_carry[26] , 
    \secondStage_carry[25] , \secondStage_carry[24] , \secondStage_carry[23] , \secondStage_carry[22] , 
    \secondStage_carry[21] , \secondStage_carry[20] , \secondStage_carry[19] , \secondStage_carry[18] , 
    \secondStage_carry[17] , \secondStage_carry[16] , \secondStage_carry[15] , \secondStage_carry[14] , 
    \secondStage_carry[13] , \secondStage_carry[12] , \secondStage_carry[11] , \secondStage_carry[10] , 
    \secondStage_carry[9] , uc_2148, uc_2149, uc_2150, uc_2151, uc_2152, uc_2153, 
    uc_2154, uc_2155, uc_2156}));
multiplyAllBits firstStage (.normalizedWires ({uc_1070, uc_1071, \normalizedWires[2045] , 
    \normalizedWires[2044] , \normalizedWires[2043] , \normalizedWires[2042] , \normalizedWires[2041] , 
    \normalizedWires[2040] , \normalizedWires[2039] , \normalizedWires[2038] , \normalizedWires[2037] , 
    \normalizedWires[2036] , \normalizedWires[2035] , \normalizedWires[2034] , \normalizedWires[2033] , 
    \normalizedWires[2032] , \normalizedWires[2031] , \normalizedWires[2030] , \normalizedWires[2029] , 
    \normalizedWires[2028] , \normalizedWires[2027] , \normalizedWires[2026] , \normalizedWires[2025] , 
    \normalizedWires[2024] , \normalizedWires[2023] , \normalizedWires[2022] , \normalizedWires[2021] , 
    \normalizedWires[2020] , \normalizedWires[2019] , \normalizedWires[2018] , \normalizedWires[2017] , 
    \normalizedWires[2016] , \normalizedWires[2015] , uc_1072, uc_1073, uc_1074, 
    uc_1075, uc_1076, uc_1077, uc_1078, uc_1079, uc_1080, uc_1081, uc_1082, uc_1083, 
    uc_1084, uc_1085, uc_1086, uc_1087, uc_1088, uc_1089, uc_1090, uc_1091, uc_1092, 
    uc_1093, uc_1094, uc_1095, uc_1096, uc_1097, uc_1098, uc_1099, uc_1100, uc_1101, 
    uc_1102, uc_1103, uc_1104, uc_1105, \normalizedWires[1980] , \normalizedWires[1979] , 
    \normalizedWires[1978] , \normalizedWires[1977] , \normalizedWires[1976] , \normalizedWires[1975] , 
    \normalizedWires[1974] , \normalizedWires[1973] , \normalizedWires[1972] , \normalizedWires[1971] , 
    \normalizedWires[1970] , \normalizedWires[1969] , \normalizedWires[1968] , \normalizedWires[1967] , 
    \normalizedWires[1966] , \normalizedWires[1965] , \normalizedWires[1964] , \normalizedWires[1963] , 
    \normalizedWires[1962] , \normalizedWires[1961] , \normalizedWires[1960] , \normalizedWires[1959] , 
    \normalizedWires[1958] , \normalizedWires[1957] , \normalizedWires[1956] , \normalizedWires[1955] , 
    \normalizedWires[1954] , \normalizedWires[1953] , \normalizedWires[1952] , \normalizedWires[1951] , 
    \normalizedWires[1950] , uc_1106, uc_1107, uc_1108, uc_1109, uc_1110, uc_1111, 
    uc_1112, uc_1113, uc_1114, uc_1115, uc_1116, uc_1117, uc_1118, uc_1119, uc_1120, 
    uc_1121, uc_1122, uc_1123, uc_1124, uc_1125, uc_1126, uc_1127, uc_1128, uc_1129, 
    uc_1130, uc_1131, uc_1132, uc_1133, uc_1134, uc_1135, uc_1136, uc_1137, uc_1138, 
    uc_1139, \normalizedWires[1915] , \normalizedWires[1914] , \normalizedWires[1913] , 
    \normalizedWires[1912] , \normalizedWires[1911] , \normalizedWires[1910] , \normalizedWires[1909] , 
    \normalizedWires[1908] , \normalizedWires[1907] , \normalizedWires[1906] , \normalizedWires[1905] , 
    \normalizedWires[1904] , \normalizedWires[1903] , \normalizedWires[1902] , \normalizedWires[1901] , 
    \normalizedWires[1900] , \normalizedWires[1899] , \normalizedWires[1898] , \normalizedWires[1897] , 
    \normalizedWires[1896] , \normalizedWires[1895] , \normalizedWires[1894] , \normalizedWires[1893] , 
    \normalizedWires[1892] , \normalizedWires[1891] , \normalizedWires[1890] , \normalizedWires[1889] , 
    \normalizedWires[1888] , \normalizedWires[1887] , \normalizedWires[1886] , \normalizedWires[1885] , 
    uc_1140, uc_1141, uc_1142, uc_1143, uc_1144, uc_1145, uc_1146, uc_1147, uc_1148, 
    uc_1149, uc_1150, uc_1151, uc_1152, uc_1153, uc_1154, uc_1155, uc_1156, uc_1157, 
    uc_1158, uc_1159, uc_1160, uc_1161, uc_1162, uc_1163, uc_1164, uc_1165, uc_1166, 
    uc_1167, uc_1168, uc_1169, uc_1170, uc_1171, uc_1172, uc_1173, \normalizedWires[1850] , 
    \normalizedWires[1849] , \normalizedWires[1848] , \normalizedWires[1847] , \normalizedWires[1846] , 
    \normalizedWires[1845] , \normalizedWires[1844] , \normalizedWires[1843] , \normalizedWires[1842] , 
    \normalizedWires[1841] , \normalizedWires[1840] , \normalizedWires[1839] , \normalizedWires[1838] , 
    \normalizedWires[1837] , \normalizedWires[1836] , \normalizedWires[1835] , \normalizedWires[1834] , 
    \normalizedWires[1833] , \normalizedWires[1832] , \normalizedWires[1831] , \normalizedWires[1830] , 
    \normalizedWires[1829] , \normalizedWires[1828] , \normalizedWires[1827] , \normalizedWires[1826] , 
    \normalizedWires[1825] , \normalizedWires[1824] , \normalizedWires[1823] , \normalizedWires[1822] , 
    \normalizedWires[1821] , \normalizedWires[1820] , uc_1174, uc_1175, uc_1176, 
    uc_1177, uc_1178, uc_1179, uc_1180, uc_1181, uc_1182, uc_1183, uc_1184, uc_1185, 
    uc_1186, uc_1187, uc_1188, uc_1189, uc_1190, uc_1191, uc_1192, uc_1193, uc_1194, 
    uc_1195, uc_1196, uc_1197, uc_1198, uc_1199, uc_1200, uc_1201, uc_1202, uc_1203, 
    uc_1204, uc_1205, uc_1206, uc_1207, \normalizedWires[1785] , \normalizedWires[1784] , 
    \normalizedWires[1783] , \normalizedWires[1782] , \normalizedWires[1781] , \normalizedWires[1780] , 
    \normalizedWires[1779] , \normalizedWires[1778] , \normalizedWires[1777] , \normalizedWires[1776] , 
    \normalizedWires[1775] , \normalizedWires[1774] , \normalizedWires[1773] , \normalizedWires[1772] , 
    \normalizedWires[1771] , \normalizedWires[1770] , \normalizedWires[1769] , \normalizedWires[1768] , 
    \normalizedWires[1767] , \normalizedWires[1766] , \normalizedWires[1765] , \normalizedWires[1764] , 
    \normalizedWires[1763] , \normalizedWires[1762] , \normalizedWires[1761] , \normalizedWires[1760] , 
    \normalizedWires[1759] , \normalizedWires[1758] , \normalizedWires[1757] , \normalizedWires[1756] , 
    \normalizedWires[1755] , uc_1208, uc_1209, uc_1210, uc_1211, uc_1212, uc_1213, 
    uc_1214, uc_1215, uc_1216, uc_1217, uc_1218, uc_1219, uc_1220, uc_1221, uc_1222, 
    uc_1223, uc_1224, uc_1225, uc_1226, uc_1227, uc_1228, uc_1229, uc_1230, uc_1231, 
    uc_1232, uc_1233, uc_1234, uc_1235, uc_1236, uc_1237, uc_1238, uc_1239, uc_1240, 
    uc_1241, \normalizedWires[1720] , \normalizedWires[1719] , \normalizedWires[1718] , 
    \normalizedWires[1717] , \normalizedWires[1716] , \normalizedWires[1715] , \normalizedWires[1714] , 
    \normalizedWires[1713] , \normalizedWires[1712] , \normalizedWires[1711] , \normalizedWires[1710] , 
    \normalizedWires[1709] , \normalizedWires[1708] , \normalizedWires[1707] , \normalizedWires[1706] , 
    \normalizedWires[1705] , \normalizedWires[1704] , \normalizedWires[1703] , \normalizedWires[1702] , 
    \normalizedWires[1701] , \normalizedWires[1700] , \normalizedWires[1699] , \normalizedWires[1698] , 
    \normalizedWires[1697] , \normalizedWires[1696] , \normalizedWires[1695] , \normalizedWires[1694] , 
    \normalizedWires[1693] , \normalizedWires[1692] , \normalizedWires[1691] , \normalizedWires[1690] , 
    uc_1242, uc_1243, uc_1244, uc_1245, uc_1246, uc_1247, uc_1248, uc_1249, uc_1250, 
    uc_1251, uc_1252, uc_1253, uc_1254, uc_1255, uc_1256, uc_1257, uc_1258, uc_1259, 
    uc_1260, uc_1261, uc_1262, uc_1263, uc_1264, uc_1265, uc_1266, uc_1267, uc_1268, 
    uc_1269, uc_1270, uc_1271, uc_1272, uc_1273, uc_1274, uc_1275, \normalizedWires[1655] , 
    \normalizedWires[1654] , \normalizedWires[1653] , \normalizedWires[1652] , \normalizedWires[1651] , 
    \normalizedWires[1650] , \normalizedWires[1649] , \normalizedWires[1648] , \normalizedWires[1647] , 
    \normalizedWires[1646] , \normalizedWires[1645] , \normalizedWires[1644] , \normalizedWires[1643] , 
    \normalizedWires[1642] , \normalizedWires[1641] , \normalizedWires[1640] , \normalizedWires[1639] , 
    \normalizedWires[1638] , \normalizedWires[1637] , \normalizedWires[1636] , \normalizedWires[1635] , 
    \normalizedWires[1634] , \normalizedWires[1633] , \normalizedWires[1632] , \normalizedWires[1631] , 
    \normalizedWires[1630] , \normalizedWires[1629] , \normalizedWires[1628] , \normalizedWires[1627] , 
    \normalizedWires[1626] , \normalizedWires[1625] , uc_1276, uc_1277, uc_1278, 
    uc_1279, uc_1280, uc_1281, uc_1282, uc_1283, uc_1284, uc_1285, uc_1286, uc_1287, 
    uc_1288, uc_1289, uc_1290, uc_1291, uc_1292, uc_1293, uc_1294, uc_1295, uc_1296, 
    uc_1297, uc_1298, uc_1299, uc_1300, uc_1301, uc_1302, uc_1303, uc_1304, uc_1305, 
    uc_1306, uc_1307, uc_1308, uc_1309, \normalizedWires[1590] , \normalizedWires[1589] , 
    \normalizedWires[1588] , \normalizedWires[1587] , \normalizedWires[1586] , \normalizedWires[1585] , 
    \normalizedWires[1584] , \normalizedWires[1583] , \normalizedWires[1582] , \normalizedWires[1581] , 
    \normalizedWires[1580] , \normalizedWires[1579] , \normalizedWires[1578] , \normalizedWires[1577] , 
    \normalizedWires[1576] , \normalizedWires[1575] , \normalizedWires[1574] , \normalizedWires[1573] , 
    \normalizedWires[1572] , \normalizedWires[1571] , \normalizedWires[1570] , \normalizedWires[1569] , 
    \normalizedWires[1568] , \normalizedWires[1567] , \normalizedWires[1566] , \normalizedWires[1565] , 
    \normalizedWires[1564] , \normalizedWires[1563] , \normalizedWires[1562] , \normalizedWires[1561] , 
    \normalizedWires[1560] , uc_1310, uc_1311, uc_1312, uc_1313, uc_1314, uc_1315, 
    uc_1316, uc_1317, uc_1318, uc_1319, uc_1320, uc_1321, uc_1322, uc_1323, uc_1324, 
    uc_1325, uc_1326, uc_1327, uc_1328, uc_1329, uc_1330, uc_1331, uc_1332, uc_1333, 
    uc_1334, uc_1335, uc_1336, uc_1337, uc_1338, uc_1339, uc_1340, uc_1341, uc_1342, 
    uc_1343, \normalizedWires[1525] , \normalizedWires[1524] , \normalizedWires[1523] , 
    \normalizedWires[1522] , \normalizedWires[1521] , \normalizedWires[1520] , \normalizedWires[1519] , 
    \normalizedWires[1518] , \normalizedWires[1517] , \normalizedWires[1516] , \normalizedWires[1515] , 
    \normalizedWires[1514] , \normalizedWires[1513] , \normalizedWires[1512] , \normalizedWires[1511] , 
    \normalizedWires[1510] , \normalizedWires[1509] , \normalizedWires[1508] , \normalizedWires[1507] , 
    \normalizedWires[1506] , \normalizedWires[1505] , \normalizedWires[1504] , \normalizedWires[1503] , 
    \normalizedWires[1502] , \normalizedWires[1501] , \normalizedWires[1500] , \normalizedWires[1499] , 
    \normalizedWires[1498] , \normalizedWires[1497] , \normalizedWires[1496] , \normalizedWires[1495] , 
    uc_1344, uc_1345, uc_1346, uc_1347, uc_1348, uc_1349, uc_1350, uc_1351, uc_1352, 
    uc_1353, uc_1354, uc_1355, uc_1356, uc_1357, uc_1358, uc_1359, uc_1360, uc_1361, 
    uc_1362, uc_1363, uc_1364, uc_1365, uc_1366, uc_1367, uc_1368, uc_1369, uc_1370, 
    uc_1371, uc_1372, uc_1373, uc_1374, uc_1375, uc_1376, uc_1377, \normalizedWires[1460] , 
    \normalizedWires[1459] , \normalizedWires[1458] , \normalizedWires[1457] , \normalizedWires[1456] , 
    \normalizedWires[1455] , \normalizedWires[1454] , \normalizedWires[1453] , \normalizedWires[1452] , 
    \normalizedWires[1451] , \normalizedWires[1450] , \normalizedWires[1449] , \normalizedWires[1448] , 
    \normalizedWires[1447] , \normalizedWires[1446] , \normalizedWires[1445] , \normalizedWires[1444] , 
    \normalizedWires[1443] , \normalizedWires[1442] , \normalizedWires[1441] , \normalizedWires[1440] , 
    \normalizedWires[1439] , \normalizedWires[1438] , \normalizedWires[1437] , \normalizedWires[1436] , 
    \normalizedWires[1435] , \normalizedWires[1434] , \normalizedWires[1433] , \normalizedWires[1432] , 
    \normalizedWires[1431] , \normalizedWires[1430] , uc_1378, uc_1379, uc_1380, 
    uc_1381, uc_1382, uc_1383, uc_1384, uc_1385, uc_1386, uc_1387, uc_1388, uc_1389, 
    uc_1390, uc_1391, uc_1392, uc_1393, uc_1394, uc_1395, uc_1396, uc_1397, uc_1398, 
    uc_1399, uc_1400, uc_1401, uc_1402, uc_1403, uc_1404, uc_1405, uc_1406, uc_1407, 
    uc_1408, uc_1409, uc_1410, uc_1411, \normalizedWires[1395] , \normalizedWires[1394] , 
    \normalizedWires[1393] , \normalizedWires[1392] , \normalizedWires[1391] , \normalizedWires[1390] , 
    \normalizedWires[1389] , \normalizedWires[1388] , \normalizedWires[1387] , \normalizedWires[1386] , 
    \normalizedWires[1385] , \normalizedWires[1384] , \normalizedWires[1383] , \normalizedWires[1382] , 
    \normalizedWires[1381] , \normalizedWires[1380] , \normalizedWires[1379] , \normalizedWires[1378] , 
    \normalizedWires[1377] , \normalizedWires[1376] , \normalizedWires[1375] , \normalizedWires[1374] , 
    \normalizedWires[1373] , \normalizedWires[1372] , \normalizedWires[1371] , \normalizedWires[1370] , 
    \normalizedWires[1369] , \normalizedWires[1368] , \normalizedWires[1367] , \normalizedWires[1366] , 
    \normalizedWires[1365] , uc_1412, uc_1413, uc_1414, uc_1415, uc_1416, uc_1417, 
    uc_1418, uc_1419, uc_1420, uc_1421, uc_1422, uc_1423, uc_1424, uc_1425, uc_1426, 
    uc_1427, uc_1428, uc_1429, uc_1430, uc_1431, uc_1432, uc_1433, uc_1434, uc_1435, 
    uc_1436, uc_1437, uc_1438, uc_1439, uc_1440, uc_1441, uc_1442, uc_1443, uc_1444, 
    uc_1445, \normalizedWires[1330] , \normalizedWires[1329] , \normalizedWires[1328] , 
    \normalizedWires[1327] , \normalizedWires[1326] , \normalizedWires[1325] , \normalizedWires[1324] , 
    \normalizedWires[1323] , \normalizedWires[1322] , \normalizedWires[1321] , \normalizedWires[1320] , 
    \normalizedWires[1319] , \normalizedWires[1318] , \normalizedWires[1317] , \normalizedWires[1316] , 
    \normalizedWires[1315] , \normalizedWires[1314] , \normalizedWires[1313] , \normalizedWires[1312] , 
    \normalizedWires[1311] , \normalizedWires[1310] , \normalizedWires[1309] , \normalizedWires[1308] , 
    \normalizedWires[1307] , \normalizedWires[1306] , \normalizedWires[1305] , \normalizedWires[1304] , 
    \normalizedWires[1303] , \normalizedWires[1302] , \normalizedWires[1301] , \normalizedWires[1300] , 
    uc_1446, uc_1447, uc_1448, uc_1449, uc_1450, uc_1451, uc_1452, uc_1453, uc_1454, 
    uc_1455, uc_1456, uc_1457, uc_1458, uc_1459, uc_1460, uc_1461, uc_1462, uc_1463, 
    uc_1464, uc_1465, uc_1466, uc_1467, uc_1468, uc_1469, uc_1470, uc_1471, uc_1472, 
    uc_1473, uc_1474, uc_1475, uc_1476, uc_1477, uc_1478, uc_1479, \normalizedWires[1265] , 
    \normalizedWires[1264] , \normalizedWires[1263] , \normalizedWires[1262] , \normalizedWires[1261] , 
    \normalizedWires[1260] , \normalizedWires[1259] , \normalizedWires[1258] , \normalizedWires[1257] , 
    \normalizedWires[1256] , \normalizedWires[1255] , \normalizedWires[1254] , \normalizedWires[1253] , 
    \normalizedWires[1252] , \normalizedWires[1251] , \normalizedWires[1250] , \normalizedWires[1249] , 
    \normalizedWires[1248] , \normalizedWires[1247] , \normalizedWires[1246] , \normalizedWires[1245] , 
    \normalizedWires[1244] , \normalizedWires[1243] , \normalizedWires[1242] , \normalizedWires[1241] , 
    \normalizedWires[1240] , \normalizedWires[1239] , \normalizedWires[1238] , \normalizedWires[1237] , 
    \normalizedWires[1236] , \normalizedWires[1235] , uc_1480, uc_1481, uc_1482, 
    uc_1483, uc_1484, uc_1485, uc_1486, uc_1487, uc_1488, uc_1489, uc_1490, uc_1491, 
    uc_1492, uc_1493, uc_1494, uc_1495, uc_1496, uc_1497, uc_1498, uc_1499, uc_1500, 
    uc_1501, uc_1502, uc_1503, uc_1504, uc_1505, uc_1506, uc_1507, uc_1508, uc_1509, 
    uc_1510, uc_1511, uc_1512, uc_1513, \normalizedWires[1200] , \normalizedWires[1199] , 
    \normalizedWires[1198] , \normalizedWires[1197] , \normalizedWires[1196] , \normalizedWires[1195] , 
    \normalizedWires[1194] , \normalizedWires[1193] , \normalizedWires[1192] , \normalizedWires[1191] , 
    \normalizedWires[1190] , \normalizedWires[1189] , \normalizedWires[1188] , \normalizedWires[1187] , 
    \normalizedWires[1186] , \normalizedWires[1185] , \normalizedWires[1184] , \normalizedWires[1183] , 
    \normalizedWires[1182] , \normalizedWires[1181] , \normalizedWires[1180] , \normalizedWires[1179] , 
    \normalizedWires[1178] , \normalizedWires[1177] , \normalizedWires[1176] , \normalizedWires[1175] , 
    \normalizedWires[1174] , \normalizedWires[1173] , \normalizedWires[1172] , \normalizedWires[1171] , 
    \normalizedWires[1170] , uc_1514, uc_1515, uc_1516, uc_1517, uc_1518, uc_1519, 
    uc_1520, uc_1521, uc_1522, uc_1523, uc_1524, uc_1525, uc_1526, uc_1527, uc_1528, 
    uc_1529, uc_1530, uc_1531, uc_1532, uc_1533, uc_1534, uc_1535, uc_1536, uc_1537, 
    uc_1538, uc_1539, uc_1540, uc_1541, uc_1542, uc_1543, uc_1544, uc_1545, uc_1546, 
    uc_1547, \normalizedWires[1135] , \normalizedWires[1134] , \normalizedWires[1133] , 
    \normalizedWires[1132] , \normalizedWires[1131] , \normalizedWires[1130] , \normalizedWires[1129] , 
    \normalizedWires[1128] , \normalizedWires[1127] , \normalizedWires[1126] , \normalizedWires[1125] , 
    \normalizedWires[1124] , \normalizedWires[1123] , \normalizedWires[1122] , \normalizedWires[1121] , 
    \normalizedWires[1120] , \normalizedWires[1119] , \normalizedWires[1118] , \normalizedWires[1117] , 
    \normalizedWires[1116] , \normalizedWires[1115] , \normalizedWires[1114] , \normalizedWires[1113] , 
    \normalizedWires[1112] , \normalizedWires[1111] , \normalizedWires[1110] , \normalizedWires[1109] , 
    \normalizedWires[1108] , \normalizedWires[1107] , \normalizedWires[1106] , \normalizedWires[1105] , 
    uc_1548, uc_1549, uc_1550, uc_1551, uc_1552, uc_1553, uc_1554, uc_1555, uc_1556, 
    uc_1557, uc_1558, uc_1559, uc_1560, uc_1561, uc_1562, uc_1563, uc_1564, uc_1565, 
    uc_1566, uc_1567, uc_1568, uc_1569, uc_1570, uc_1571, uc_1572, uc_1573, uc_1574, 
    uc_1575, uc_1576, uc_1577, uc_1578, uc_1579, uc_1580, uc_1581, \normalizedWires[1070] , 
    \normalizedWires[1069] , \normalizedWires[1068] , \normalizedWires[1067] , \normalizedWires[1066] , 
    \normalizedWires[1065] , \normalizedWires[1064] , \normalizedWires[1063] , \normalizedWires[1062] , 
    \normalizedWires[1061] , \normalizedWires[1060] , \normalizedWires[1059] , \normalizedWires[1058] , 
    \normalizedWires[1057] , \normalizedWires[1056] , \normalizedWires[1055] , \normalizedWires[1054] , 
    \normalizedWires[1053] , \normalizedWires[1052] , \normalizedWires[1051] , \normalizedWires[1050] , 
    \normalizedWires[1049] , \normalizedWires[1048] , \normalizedWires[1047] , \normalizedWires[1046] , 
    \normalizedWires[1045] , \normalizedWires[1044] , \normalizedWires[1043] , \normalizedWires[1042] , 
    \normalizedWires[1041] , \normalizedWires[1040] , uc_1582, uc_1583, uc_1584, 
    uc_1585, uc_1586, uc_1587, uc_1588, uc_1589, uc_1590, uc_1591, uc_1592, uc_1593, 
    uc_1594, uc_1595, uc_1596, uc_1597, uc_1598, uc_1599, uc_1600, uc_1601, uc_1602, 
    uc_1603, uc_1604, uc_1605, uc_1606, uc_1607, uc_1608, uc_1609, uc_1610, uc_1611, 
    uc_1612, uc_1613, uc_1614, uc_1615, \normalizedWires[1005] , \normalizedWires[1004] , 
    \normalizedWires[1003] , \normalizedWires[1002] , \normalizedWires[1001] , \normalizedWires[1000] , 
    \normalizedWires[999] , \normalizedWires[998] , \normalizedWires[997] , \normalizedWires[996] , 
    \normalizedWires[995] , \normalizedWires[994] , \normalizedWires[993] , \normalizedWires[992] , 
    \normalizedWires[991] , \normalizedWires[990] , \normalizedWires[989] , \normalizedWires[988] , 
    \normalizedWires[987] , \normalizedWires[986] , \normalizedWires[985] , \normalizedWires[984] , 
    \normalizedWires[983] , \normalizedWires[982] , \normalizedWires[981] , \normalizedWires[980] , 
    \normalizedWires[979] , \normalizedWires[978] , \normalizedWires[977] , \normalizedWires[976] , 
    \normalizedWires[975] , uc_1616, uc_1617, uc_1618, uc_1619, uc_1620, uc_1621, 
    uc_1622, uc_1623, uc_1624, uc_1625, uc_1626, uc_1627, uc_1628, uc_1629, uc_1630, 
    uc_1631, uc_1632, uc_1633, uc_1634, uc_1635, uc_1636, uc_1637, uc_1638, uc_1639, 
    uc_1640, uc_1641, uc_1642, uc_1643, uc_1644, uc_1645, uc_1646, uc_1647, uc_1648, 
    uc_1649, \normalizedWires[940] , \normalizedWires[939] , \normalizedWires[938] , 
    \normalizedWires[937] , \normalizedWires[936] , \normalizedWires[935] , \normalizedWires[934] , 
    \normalizedWires[933] , \normalizedWires[932] , \normalizedWires[931] , \normalizedWires[930] , 
    \normalizedWires[929] , \normalizedWires[928] , \normalizedWires[927] , \normalizedWires[926] , 
    \normalizedWires[925] , \normalizedWires[924] , \normalizedWires[923] , \normalizedWires[922] , 
    \normalizedWires[921] , \normalizedWires[920] , \normalizedWires[919] , \normalizedWires[918] , 
    \normalizedWires[917] , \normalizedWires[916] , \normalizedWires[915] , \normalizedWires[914] , 
    \normalizedWires[913] , \normalizedWires[912] , \normalizedWires[911] , \normalizedWires[910] , 
    uc_1650, uc_1651, uc_1652, uc_1653, uc_1654, uc_1655, uc_1656, uc_1657, uc_1658, 
    uc_1659, uc_1660, uc_1661, uc_1662, uc_1663, uc_1664, uc_1665, uc_1666, uc_1667, 
    uc_1668, uc_1669, uc_1670, uc_1671, uc_1672, uc_1673, uc_1674, uc_1675, uc_1676, 
    uc_1677, uc_1678, uc_1679, uc_1680, uc_1681, uc_1682, uc_1683, \normalizedWires[875] , 
    \normalizedWires[874] , \normalizedWires[873] , \normalizedWires[872] , \normalizedWires[871] , 
    \normalizedWires[870] , \normalizedWires[869] , \normalizedWires[868] , \normalizedWires[867] , 
    \normalizedWires[866] , \normalizedWires[865] , \normalizedWires[864] , \normalizedWires[863] , 
    \normalizedWires[862] , \normalizedWires[861] , \normalizedWires[860] , \normalizedWires[859] , 
    \normalizedWires[858] , \normalizedWires[857] , \normalizedWires[856] , \normalizedWires[855] , 
    \normalizedWires[854] , \normalizedWires[853] , \normalizedWires[852] , \normalizedWires[851] , 
    \normalizedWires[850] , \normalizedWires[849] , \normalizedWires[848] , \normalizedWires[847] , 
    \normalizedWires[846] , \normalizedWires[845] , uc_1684, uc_1685, uc_1686, uc_1687, 
    uc_1688, uc_1689, uc_1690, uc_1691, uc_1692, uc_1693, uc_1694, uc_1695, uc_1696, 
    uc_1697, uc_1698, uc_1699, uc_1700, uc_1701, uc_1702, uc_1703, uc_1704, uc_1705, 
    uc_1706, uc_1707, uc_1708, uc_1709, uc_1710, uc_1711, uc_1712, uc_1713, uc_1714, 
    uc_1715, uc_1716, uc_1717, \normalizedWires[810] , \normalizedWires[809] , \normalizedWires[808] , 
    \normalizedWires[807] , \normalizedWires[806] , \normalizedWires[805] , \normalizedWires[804] , 
    \normalizedWires[803] , \normalizedWires[802] , \normalizedWires[801] , \normalizedWires[800] , 
    \normalizedWires[799] , \normalizedWires[798] , \normalizedWires[797] , \normalizedWires[796] , 
    \normalizedWires[795] , \normalizedWires[794] , \normalizedWires[793] , \normalizedWires[792] , 
    \normalizedWires[791] , \normalizedWires[790] , \normalizedWires[789] , \normalizedWires[788] , 
    \normalizedWires[787] , \normalizedWires[786] , \normalizedWires[785] , \normalizedWires[784] , 
    \normalizedWires[783] , \normalizedWires[782] , \normalizedWires[781] , \normalizedWires[780] , 
    uc_1718, uc_1719, uc_1720, uc_1721, uc_1722, uc_1723, uc_1724, uc_1725, uc_1726, 
    uc_1727, uc_1728, uc_1729, uc_1730, uc_1731, uc_1732, uc_1733, uc_1734, uc_1735, 
    uc_1736, uc_1737, uc_1738, uc_1739, uc_1740, uc_1741, uc_1742, uc_1743, uc_1744, 
    uc_1745, uc_1746, uc_1747, uc_1748, uc_1749, uc_1750, uc_1751, \normalizedWires[745] , 
    \normalizedWires[744] , \normalizedWires[743] , \normalizedWires[742] , \normalizedWires[741] , 
    \normalizedWires[740] , \normalizedWires[739] , \normalizedWires[738] , \normalizedWires[737] , 
    \normalizedWires[736] , \normalizedWires[735] , \normalizedWires[734] , \normalizedWires[733] , 
    \normalizedWires[732] , \normalizedWires[731] , \normalizedWires[730] , \normalizedWires[729] , 
    \normalizedWires[728] , \normalizedWires[727] , \normalizedWires[726] , \normalizedWires[725] , 
    \normalizedWires[724] , \normalizedWires[723] , \normalizedWires[722] , \normalizedWires[721] , 
    \normalizedWires[720] , \normalizedWires[719] , \normalizedWires[718] , \normalizedWires[717] , 
    \normalizedWires[716] , \normalizedWires[715] , uc_1752, uc_1753, uc_1754, uc_1755, 
    uc_1756, uc_1757, uc_1758, uc_1759, uc_1760, uc_1761, uc_1762, uc_1763, uc_1764, 
    uc_1765, uc_1766, uc_1767, uc_1768, uc_1769, uc_1770, uc_1771, uc_1772, uc_1773, 
    uc_1774, uc_1775, uc_1776, uc_1777, uc_1778, uc_1779, uc_1780, uc_1781, uc_1782, 
    uc_1783, uc_1784, uc_1785, \normalizedWires[680] , \normalizedWires[679] , \normalizedWires[678] , 
    \normalizedWires[677] , \normalizedWires[676] , \normalizedWires[675] , \normalizedWires[674] , 
    \normalizedWires[673] , \normalizedWires[672] , \normalizedWires[671] , \normalizedWires[670] , 
    \normalizedWires[669] , \normalizedWires[668] , \normalizedWires[667] , \normalizedWires[666] , 
    \normalizedWires[665] , \normalizedWires[664] , \normalizedWires[663] , \normalizedWires[662] , 
    \normalizedWires[661] , \normalizedWires[660] , \normalizedWires[659] , \normalizedWires[658] , 
    \normalizedWires[657] , \normalizedWires[656] , \normalizedWires[655] , \normalizedWires[654] , 
    \normalizedWires[653] , \normalizedWires[652] , \normalizedWires[651] , \normalizedWires[650] , 
    uc_1786, uc_1787, uc_1788, uc_1789, uc_1790, uc_1791, uc_1792, uc_1793, uc_1794, 
    uc_1795, uc_1796, uc_1797, uc_1798, uc_1799, uc_1800, uc_1801, uc_1802, uc_1803, 
    uc_1804, uc_1805, uc_1806, uc_1807, uc_1808, uc_1809, uc_1810, uc_1811, uc_1812, 
    uc_1813, uc_1814, uc_1815, uc_1816, uc_1817, uc_1818, uc_1819, \normalizedWires[615] , 
    \normalizedWires[614] , \normalizedWires[613] , \normalizedWires[612] , \normalizedWires[611] , 
    \normalizedWires[610] , \normalizedWires[609] , \normalizedWires[608] , \normalizedWires[607] , 
    \normalizedWires[606] , \normalizedWires[605] , \normalizedWires[604] , \normalizedWires[603] , 
    \normalizedWires[602] , \normalizedWires[601] , \normalizedWires[600] , \normalizedWires[599] , 
    \normalizedWires[598] , \normalizedWires[597] , \normalizedWires[596] , \normalizedWires[595] , 
    \normalizedWires[594] , \normalizedWires[593] , \normalizedWires[592] , \normalizedWires[591] , 
    \normalizedWires[590] , \normalizedWires[589] , \normalizedWires[588] , \normalizedWires[587] , 
    \normalizedWires[586] , \normalizedWires[585] , uc_1820, uc_1821, uc_1822, uc_1823, 
    uc_1824, uc_1825, uc_1826, uc_1827, uc_1828, uc_1829, uc_1830, uc_1831, uc_1832, 
    uc_1833, uc_1834, uc_1835, uc_1836, uc_1837, uc_1838, uc_1839, uc_1840, uc_1841, 
    uc_1842, uc_1843, uc_1844, uc_1845, uc_1846, uc_1847, uc_1848, uc_1849, uc_1850, 
    uc_1851, uc_1852, uc_1853, \normalizedWires[550] , \normalizedWires[549] , \normalizedWires[548] , 
    \normalizedWires[547] , \normalizedWires[546] , \normalizedWires[545] , \normalizedWires[544] , 
    \normalizedWires[543] , \normalizedWires[542] , \normalizedWires[541] , \normalizedWires[540] , 
    \normalizedWires[539] , \normalizedWires[538] , \normalizedWires[537] , \normalizedWires[536] , 
    \normalizedWires[535] , \normalizedWires[534] , \normalizedWires[533] , \normalizedWires[532] , 
    \normalizedWires[531] , \normalizedWires[530] , \normalizedWires[529] , \normalizedWires[528] , 
    \normalizedWires[527] , \normalizedWires[526] , \normalizedWires[525] , \normalizedWires[524] , 
    \normalizedWires[523] , \normalizedWires[522] , \normalizedWires[521] , \normalizedWires[520] , 
    uc_1854, uc_1855, uc_1856, uc_1857, uc_1858, uc_1859, uc_1860, uc_1861, uc_1862, 
    uc_1863, uc_1864, uc_1865, uc_1866, uc_1867, uc_1868, uc_1869, uc_1870, uc_1871, 
    uc_1872, uc_1873, uc_1874, uc_1875, uc_1876, uc_1877, uc_1878, uc_1879, uc_1880, 
    uc_1881, uc_1882, uc_1883, uc_1884, uc_1885, uc_1886, uc_1887, \normalizedWires[485] , 
    \normalizedWires[484] , \normalizedWires[483] , \normalizedWires[482] , \normalizedWires[481] , 
    \normalizedWires[480] , \normalizedWires[479] , \normalizedWires[478] , \normalizedWires[477] , 
    \normalizedWires[476] , \normalizedWires[475] , \normalizedWires[474] , \normalizedWires[473] , 
    \normalizedWires[472] , \normalizedWires[471] , \normalizedWires[470] , \normalizedWires[469] , 
    \normalizedWires[468] , \normalizedWires[467] , \normalizedWires[466] , \normalizedWires[465] , 
    \normalizedWires[464] , \normalizedWires[463] , \normalizedWires[462] , \normalizedWires[461] , 
    \normalizedWires[460] , \normalizedWires[459] , \normalizedWires[458] , \normalizedWires[457] , 
    \normalizedWires[456] , \normalizedWires[455] , uc_1888, uc_1889, uc_1890, uc_1891, 
    uc_1892, uc_1893, uc_1894, uc_1895, uc_1896, uc_1897, uc_1898, uc_1899, uc_1900, 
    uc_1901, uc_1902, uc_1903, uc_1904, uc_1905, uc_1906, uc_1907, uc_1908, uc_1909, 
    uc_1910, uc_1911, uc_1912, uc_1913, uc_1914, uc_1915, uc_1916, uc_1917, uc_1918, 
    uc_1919, uc_1920, uc_1921, \normalizedWires[420] , \normalizedWires[419] , \normalizedWires[418] , 
    \normalizedWires[417] , \normalizedWires[416] , \normalizedWires[415] , \normalizedWires[414] , 
    \normalizedWires[413] , \normalizedWires[412] , \normalizedWires[411] , \normalizedWires[410] , 
    \normalizedWires[409] , \normalizedWires[408] , \normalizedWires[407] , \normalizedWires[406] , 
    \normalizedWires[405] , \normalizedWires[404] , \normalizedWires[403] , \normalizedWires[402] , 
    \normalizedWires[401] , \normalizedWires[400] , \normalizedWires[399] , \normalizedWires[398] , 
    \normalizedWires[397] , \normalizedWires[396] , \normalizedWires[395] , \normalizedWires[394] , 
    \normalizedWires[393] , \normalizedWires[392] , \normalizedWires[391] , \normalizedWires[390] , 
    uc_1922, uc_1923, uc_1924, uc_1925, uc_1926, uc_1927, uc_1928, uc_1929, uc_1930, 
    uc_1931, uc_1932, uc_1933, uc_1934, uc_1935, uc_1936, uc_1937, uc_1938, uc_1939, 
    uc_1940, uc_1941, uc_1942, uc_1943, uc_1944, uc_1945, uc_1946, uc_1947, uc_1948, 
    uc_1949, uc_1950, uc_1951, uc_1952, uc_1953, uc_1954, uc_1955, \normalizedWires[355] , 
    \normalizedWires[354] , \normalizedWires[353] , \normalizedWires[352] , \normalizedWires[351] , 
    \normalizedWires[350] , \normalizedWires[349] , \normalizedWires[348] , \normalizedWires[347] , 
    \normalizedWires[346] , \normalizedWires[345] , \normalizedWires[344] , \normalizedWires[343] , 
    \normalizedWires[342] , \normalizedWires[341] , \normalizedWires[340] , \normalizedWires[339] , 
    \normalizedWires[338] , \normalizedWires[337] , \normalizedWires[336] , \normalizedWires[335] , 
    \normalizedWires[334] , \normalizedWires[333] , \normalizedWires[332] , \normalizedWires[331] , 
    \normalizedWires[330] , \normalizedWires[329] , \normalizedWires[328] , \normalizedWires[327] , 
    \normalizedWires[326] , \normalizedWires[325] , uc_1956, uc_1957, uc_1958, uc_1959, 
    uc_1960, uc_1961, uc_1962, uc_1963, uc_1964, uc_1965, uc_1966, uc_1967, uc_1968, 
    uc_1969, uc_1970, uc_1971, uc_1972, uc_1973, uc_1974, uc_1975, uc_1976, uc_1977, 
    uc_1978, uc_1979, uc_1980, uc_1981, uc_1982, uc_1983, uc_1984, uc_1985, uc_1986, 
    uc_1987, uc_1988, uc_1989, \normalizedWires[290] , \normalizedWires[289] , \normalizedWires[288] , 
    \normalizedWires[287] , \normalizedWires[286] , \normalizedWires[285] , \normalizedWires[284] , 
    \normalizedWires[283] , \normalizedWires[282] , \normalizedWires[281] , \normalizedWires[280] , 
    \normalizedWires[279] , \normalizedWires[278] , \normalizedWires[277] , \normalizedWires[276] , 
    \normalizedWires[275] , \normalizedWires[274] , \normalizedWires[273] , \normalizedWires[272] , 
    \normalizedWires[271] , \normalizedWires[270] , \normalizedWires[269] , \normalizedWires[268] , 
    \normalizedWires[267] , \normalizedWires[266] , \normalizedWires[265] , \normalizedWires[264] , 
    \normalizedWires[263] , \normalizedWires[262] , \normalizedWires[261] , \normalizedWires[260] , 
    uc_1990, uc_1991, uc_1992, uc_1993, uc_1994, uc_1995, uc_1996, uc_1997, uc_1998, 
    uc_1999, uc_2000, uc_2001, uc_2002, uc_2003, uc_2004, uc_2005, uc_2006, uc_2007, 
    uc_2008, uc_2009, uc_2010, uc_2011, uc_2012, uc_2013, uc_2014, uc_2015, uc_2016, 
    uc_2017, uc_2018, uc_2019, uc_2020, uc_2021, uc_2022, uc_2023, \normalizedWires[225] , 
    \normalizedWires[224] , \normalizedWires[223] , \normalizedWires[222] , \normalizedWires[221] , 
    \normalizedWires[220] , \normalizedWires[219] , \normalizedWires[218] , \normalizedWires[217] , 
    \normalizedWires[216] , \normalizedWires[215] , \normalizedWires[214] , \normalizedWires[213] , 
    \normalizedWires[212] , \normalizedWires[211] , \normalizedWires[210] , \normalizedWires[209] , 
    \normalizedWires[208] , \normalizedWires[207] , \normalizedWires[206] , \normalizedWires[205] , 
    \normalizedWires[204] , \normalizedWires[203] , \normalizedWires[202] , \normalizedWires[201] , 
    \normalizedWires[200] , \normalizedWires[199] , \normalizedWires[198] , \normalizedWires[197] , 
    \normalizedWires[196] , \normalizedWires[195] , uc_2024, uc_2025, uc_2026, uc_2027, 
    uc_2028, uc_2029, uc_2030, uc_2031, uc_2032, uc_2033, uc_2034, uc_2035, uc_2036, 
    uc_2037, uc_2038, uc_2039, uc_2040, uc_2041, uc_2042, uc_2043, uc_2044, uc_2045, 
    uc_2046, uc_2047, uc_2048, uc_2049, uc_2050, uc_2051, uc_2052, uc_2053, uc_2054, 
    uc_2055, uc_2056, uc_2057, \normalizedWires[160] , \normalizedWires[159] , \normalizedWires[158] , 
    \normalizedWires[157] , \normalizedWires[156] , \normalizedWires[155] , \normalizedWires[154] , 
    \normalizedWires[153] , \normalizedWires[152] , \normalizedWires[151] , \normalizedWires[150] , 
    \normalizedWires[149] , \normalizedWires[148] , \normalizedWires[147] , \normalizedWires[146] , 
    \normalizedWires[145] , \normalizedWires[144] , \normalizedWires[143] , \normalizedWires[142] , 
    \normalizedWires[141] , \normalizedWires[140] , \normalizedWires[139] , \normalizedWires[138] , 
    \normalizedWires[137] , \normalizedWires[136] , \normalizedWires[135] , \normalizedWires[134] , 
    \normalizedWires[133] , \normalizedWires[132] , \normalizedWires[131] , \normalizedWires[130] , 
    uc_2058, uc_2059, uc_2060, uc_2061, uc_2062, uc_2063, uc_2064, uc_2065, uc_2066, 
    uc_2067, uc_2068, uc_2069, uc_2070, uc_2071, uc_2072, uc_2073, uc_2074, uc_2075, 
    uc_2076, uc_2077, uc_2078, uc_2079, uc_2080, uc_2081, uc_2082, uc_2083, uc_2084, 
    uc_2085, uc_2086, uc_2087, uc_2088, uc_2089, uc_2090, uc_2091, \normalizedWires[95] , 
    \normalizedWires[94] , \normalizedWires[93] , \normalizedWires[92] , \normalizedWires[91] , 
    \normalizedWires[90] , \normalizedWires[89] , \normalizedWires[88] , \normalizedWires[87] , 
    \normalizedWires[86] , \normalizedWires[85] , \normalizedWires[84] , \normalizedWires[83] , 
    \normalizedWires[82] , \normalizedWires[81] , \normalizedWires[80] , \normalizedWires[79] , 
    \normalizedWires[78] , \normalizedWires[77] , \normalizedWires[76] , \normalizedWires[75] , 
    \normalizedWires[74] , \normalizedWires[73] , \normalizedWires[72] , \normalizedWires[71] , 
    \normalizedWires[70] , \normalizedWires[69] , \normalizedWires[68] , \normalizedWires[67] , 
    \normalizedWires[66] , \normalizedWires[65] , uc_2092, uc_2093, uc_2094, uc_2095, 
    uc_2096, uc_2097, uc_2098, uc_2099, uc_2100, uc_2101, uc_2102, uc_2103, uc_2104, 
    uc_2105, uc_2106, uc_2107, uc_2108, uc_2109, uc_2110, uc_2111, uc_2112, uc_2113, 
    uc_2114, uc_2115, uc_2116, uc_2117, uc_2118, uc_2119, uc_2120, uc_2121, uc_2122, 
    uc_2123, uc_2124, uc_2125, \normalizedWires[30] , \normalizedWires[29] , \normalizedWires[28] , 
    \normalizedWires[27] , \normalizedWires[26] , \normalizedWires[25] , \normalizedWires[24] , 
    \normalizedWires[23] , \normalizedWires[22] , \normalizedWires[21] , \normalizedWires[20] , 
    \normalizedWires[19] , \normalizedWires[18] , \normalizedWires[17] , \normalizedWires[16] , 
    \normalizedWires[15] , \normalizedWires[14] , \normalizedWires[13] , \normalizedWires[12] , 
    \normalizedWires[11] , \normalizedWires[10] , \normalizedWires[9] , \normalizedWires[8] , 
    \normalizedWires[7] , \normalizedWires[6] , \normalizedWires[5] , \normalizedWires[4] , 
    \normalizedWires[3] , \normalizedWires[2] , \normalizedWires[1] , n_0_316}), .A ({
    uc_2126, \A_imm[30] , \A_imm[29] , \A_imm[28] , \A_imm[27] , CLOCK_slo__mro_n3162, 
    slo__sro_n405, CLOCK_slo__sro_n3065, CLOCK_slo__sro_n3369, \A_imm[22] , slo__sro_n667, 
    slo__sro_n363, slo__sro_n381, slo__sro_n538, CLOCK_slo__mro_n2292, slo__sro_n1079, 
    slo__sro_n1026, CLOCK_slo__mro_n2310, slo__sro_n1120, \A_imm[12] , \A_imm[11] , 
    slo__sro_n558, \A_imm[9] , \A_imm[8] , \A_imm[7] , \A_imm[6] , \A_imm[5] , \A_imm[4] , 
    \A_imm[3] , \A_imm[2] , \A_imm[1] , n_0_256}), .B ({\B_imm[31] , \B_imm[30] , 
    \B_imm[29] , \B_imm[28] , \B_imm[27] , \B_imm[26] , slo__sro_n700, CLOCK_slo__sro_n2793, 
    \B_imm[23] , slo__sro_n513, slo__sro_n1150, \B_imm[20] , \B_imm[19] , \B_imm[18] , 
    \B_imm[17] , CLOCK_slo__sro_n2682, CLOCK_slo__sro_n2298, \B_imm[14] , \B_imm[13] , 
    \B_imm[12] , \B_imm[11] , slo__sro_n420, slo__sro_n1186, \B_imm[8] , CLOCK_slo__sro_n2212, 
    CLOCK_slo__sro_n2841, \B_imm[5] , \B_imm[4] , \B_imm[3] , \B_imm[2] , \B_imm[1] , 
    slo__n619}), .B_7_PP_0 (CLOCK_slo__sro_n2212), .B_24_PP_0 (CLOCK_slo__sro_n2793)
    , .B_4_PP_0 (\B_imm[4] ));
addIntermedaiteWires secondStage (.Res ({uc_0, uc_1, \secondStage_Res[61] , \secondStage_Res[60] , 
    \secondStage_Res[59] , \secondStage_Res[58] , \secondStage_Res[57] , \secondStage_Res[56] , 
    \secondStage_Res[55] , \secondStage_Res[54] , \secondStage_Res[53] , \secondStage_Res[52] , 
    \secondStage_Res[51] , \secondStage_Res[50] , \secondStage_Res[49] , \secondStage_Res[48] , 
    \secondStage_Res[47] , \secondStage_Res[46] , \secondStage_Res[45] , \secondStage_Res[44] , 
    \secondStage_Res[43] , \secondStage_Res[42] , \secondStage_Res[41] , \secondStage_Res[40] , 
    \secondStage_Res[39] , \secondStage_Res[38] , \secondStage_Res[37] , \secondStage_Res[36] , 
    \secondStage_Res[35] , \secondStage_Res[34] , \secondStage_Res[33] , \secondStage_Res[32] , 
    \secondStage_Res[31] , \secondStage_Res[30] , \secondStage_Res[29] , \secondStage_Res[28] , 
    \secondStage_Res[27] , \secondStage_Res[26] , \secondStage_Res[25] , \secondStage_Res[24] , 
    \secondStage_Res[23] , \secondStage_Res[22] , \secondStage_Res[21] , \secondStage_Res[20] , 
    \secondStage_Res[19] , \secondStage_Res[18] , \secondStage_Res[17] , \secondStage_Res[16] , 
    \secondStage_Res[15] , \secondStage_Res[14] , \secondStage_Res[13] , \secondStage_Res[12] , 
    \secondStage_Res[11] , \secondStage_Res[10] , \secondStage_Res[9] , \secondStage_Res[8] , 
    \secondStage_Res[7] , \secondStage_Res[6] , \secondStage_Res[5] , \secondStage_Res[4] , 
    \secondStage_Res[3] , \secondStage_Res[2] , \secondStage_Res[1] , uc_2}), .carry ({
    uc_3, \secondStage_carry[62] , \secondStage_carry[61] , \secondStage_carry[60] , 
    \secondStage_carry[59] , \secondStage_carry[58] , \secondStage_carry[57] , \secondStage_carry[56] , 
    \secondStage_carry[55] , \secondStage_carry[54] , \secondStage_carry[53] , \secondStage_carry[52] , 
    \secondStage_carry[51] , \secondStage_carry[50] , \secondStage_carry[49] , \secondStage_carry[48] , 
    \secondStage_carry[47] , \secondStage_carry[46] , \secondStage_carry[45] , \secondStage_carry[44] , 
    \secondStage_carry[43] , \secondStage_carry[42] , \secondStage_carry[41] , \secondStage_carry[40] , 
    \secondStage_carry[39] , \secondStage_carry[38] , \secondStage_carry[37] , \secondStage_carry[36] , 
    \secondStage_carry[35] , \secondStage_carry[34] , \secondStage_carry[33] , \secondStage_carry[32] , 
    \secondStage_carry[31] , \secondStage_carry[30] , \secondStage_carry[29] , \secondStage_carry[28] , 
    \secondStage_carry[27] , \secondStage_carry[26] , \secondStage_carry[25] , \secondStage_carry[24] , 
    \secondStage_carry[23] , \secondStage_carry[22] , \secondStage_carry[21] , \secondStage_carry[20] , 
    \secondStage_carry[19] , \secondStage_carry[18] , \secondStage_carry[17] , \secondStage_carry[16] , 
    \secondStage_carry[15] , \secondStage_carry[14] , \secondStage_carry[13] , \secondStage_carry[12] , 
    \secondStage_carry[11] , \secondStage_carry[10] , \secondStage_carry[9] , uc_4, 
    uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12}), .normalizedWires ({uc_13, 
    uc_14, \normalizedWires[2045] , \normalizedWires[2044] , \normalizedWires[2043] , 
    \normalizedWires[2042] , \normalizedWires[2041] , \normalizedWires[2040] , \normalizedWires[2039] , 
    \normalizedWires[2038] , \normalizedWires[2037] , \normalizedWires[2036] , \normalizedWires[2035] , 
    \normalizedWires[2034] , \normalizedWires[2033] , \normalizedWires[2032] , \normalizedWires[2031] , 
    \normalizedWires[2030] , \normalizedWires[2029] , \normalizedWires[2028] , \normalizedWires[2027] , 
    \normalizedWires[2026] , \normalizedWires[2025] , \normalizedWires[2024] , \normalizedWires[2023] , 
    \normalizedWires[2022] , \normalizedWires[2021] , \normalizedWires[2020] , \normalizedWires[2019] , 
    \normalizedWires[2018] , \normalizedWires[2017] , \normalizedWires[2016] , \normalizedWires[2015] , 
    uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, 
    uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, 
    uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, 
    uc_48, \normalizedWires[1980] , \normalizedWires[1979] , \normalizedWires[1978] , 
    \normalizedWires[1977] , \normalizedWires[1976] , \normalizedWires[1975] , \normalizedWires[1974] , 
    \normalizedWires[1973] , \normalizedWires[1972] , \normalizedWires[1971] , \normalizedWires[1970] , 
    \normalizedWires[1969] , \normalizedWires[1968] , \normalizedWires[1967] , \normalizedWires[1966] , 
    \normalizedWires[1965] , \normalizedWires[1964] , \normalizedWires[1963] , \normalizedWires[1962] , 
    \normalizedWires[1961] , \normalizedWires[1960] , \normalizedWires[1959] , \normalizedWires[1958] , 
    \normalizedWires[1957] , \normalizedWires[1956] , \normalizedWires[1955] , \normalizedWires[1954] , 
    \normalizedWires[1953] , \normalizedWires[1952] , \normalizedWires[1951] , \normalizedWires[1950] , 
    uc_49, uc_50, uc_51, uc_52, uc_53, uc_54, uc_55, uc_56, uc_57, uc_58, uc_59, 
    uc_60, uc_61, uc_62, uc_63, uc_64, uc_65, uc_66, uc_67, uc_68, uc_69, uc_70, 
    uc_71, uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, uc_79, uc_80, uc_81, 
    uc_82, \normalizedWires[1915] , \normalizedWires[1914] , \normalizedWires[1913] , 
    \normalizedWires[1912] , \normalizedWires[1911] , \normalizedWires[1910] , \normalizedWires[1909] , 
    \normalizedWires[1908] , \normalizedWires[1907] , \normalizedWires[1906] , \normalizedWires[1905] , 
    \normalizedWires[1904] , \normalizedWires[1903] , \normalizedWires[1902] , \normalizedWires[1901] , 
    \normalizedWires[1900] , \normalizedWires[1899] , \normalizedWires[1898] , \normalizedWires[1897] , 
    \normalizedWires[1896] , \normalizedWires[1895] , \normalizedWires[1894] , \normalizedWires[1893] , 
    \normalizedWires[1892] , \normalizedWires[1891] , \normalizedWires[1890] , \normalizedWires[1889] , 
    \normalizedWires[1888] , \normalizedWires[1887] , \normalizedWires[1886] , \normalizedWires[1885] , 
    uc_83, uc_84, uc_85, uc_86, uc_87, uc_88, uc_89, uc_90, uc_91, uc_92, uc_93, 
    uc_94, uc_95, uc_96, uc_97, uc_98, uc_99, uc_100, uc_101, uc_102, uc_103, uc_104, 
    uc_105, uc_106, uc_107, uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, uc_114, 
    uc_115, uc_116, \normalizedWires[1850] , \normalizedWires[1849] , \normalizedWires[1848] , 
    \normalizedWires[1847] , \normalizedWires[1846] , \normalizedWires[1845] , \normalizedWires[1844] , 
    \normalizedWires[1843] , \normalizedWires[1842] , \normalizedWires[1841] , \normalizedWires[1840] , 
    \normalizedWires[1839] , \normalizedWires[1838] , \normalizedWires[1837] , \normalizedWires[1836] , 
    \normalizedWires[1835] , \normalizedWires[1834] , \normalizedWires[1833] , \normalizedWires[1832] , 
    \normalizedWires[1831] , \normalizedWires[1830] , \normalizedWires[1829] , \normalizedWires[1828] , 
    \normalizedWires[1827] , \normalizedWires[1826] , \normalizedWires[1825] , \normalizedWires[1824] , 
    \normalizedWires[1823] , \normalizedWires[1822] , \normalizedWires[1821] , \normalizedWires[1820] , 
    uc_117, uc_118, uc_119, uc_120, uc_121, uc_122, uc_123, uc_124, uc_125, uc_126, 
    uc_127, uc_128, uc_129, uc_130, uc_131, uc_132, uc_133, uc_134, uc_135, uc_136, 
    uc_137, uc_138, uc_139, uc_140, uc_141, uc_142, uc_143, uc_144, uc_145, uc_146, 
    uc_147, uc_148, uc_149, uc_150, \normalizedWires[1785] , \normalizedWires[1784] , 
    \normalizedWires[1783] , \normalizedWires[1782] , \normalizedWires[1781] , \normalizedWires[1780] , 
    \normalizedWires[1779] , \normalizedWires[1778] , \normalizedWires[1777] , \normalizedWires[1776] , 
    \normalizedWires[1775] , \normalizedWires[1774] , \normalizedWires[1773] , \normalizedWires[1772] , 
    \normalizedWires[1771] , \normalizedWires[1770] , \normalizedWires[1769] , \normalizedWires[1768] , 
    \normalizedWires[1767] , \normalizedWires[1766] , \normalizedWires[1765] , \normalizedWires[1764] , 
    \normalizedWires[1763] , \normalizedWires[1762] , \normalizedWires[1761] , \normalizedWires[1760] , 
    \normalizedWires[1759] , \normalizedWires[1758] , \normalizedWires[1757] , \normalizedWires[1756] , 
    \normalizedWires[1755] , uc_151, uc_152, uc_153, uc_154, uc_155, uc_156, uc_157, 
    uc_158, uc_159, uc_160, uc_161, uc_162, uc_163, uc_164, uc_165, uc_166, uc_167, 
    uc_168, uc_169, uc_170, uc_171, uc_172, uc_173, uc_174, uc_175, uc_176, uc_177, 
    uc_178, uc_179, uc_180, uc_181, uc_182, uc_183, uc_184, \normalizedWires[1720] , 
    \normalizedWires[1719] , \normalizedWires[1718] , \normalizedWires[1717] , \normalizedWires[1716] , 
    \normalizedWires[1715] , \normalizedWires[1714] , \normalizedWires[1713] , \normalizedWires[1712] , 
    \normalizedWires[1711] , \normalizedWires[1710] , \normalizedWires[1709] , \normalizedWires[1708] , 
    \normalizedWires[1707] , \normalizedWires[1706] , \normalizedWires[1705] , \normalizedWires[1704] , 
    \normalizedWires[1703] , \normalizedWires[1702] , \normalizedWires[1701] , \normalizedWires[1700] , 
    \normalizedWires[1699] , \normalizedWires[1698] , \normalizedWires[1697] , \normalizedWires[1696] , 
    \normalizedWires[1695] , \normalizedWires[1694] , \normalizedWires[1693] , \normalizedWires[1692] , 
    \normalizedWires[1691] , \normalizedWires[1690] , uc_185, uc_186, uc_187, uc_188, 
    uc_189, uc_190, uc_191, uc_192, uc_193, uc_194, uc_195, uc_196, uc_197, uc_198, 
    uc_199, uc_200, uc_201, uc_202, uc_203, uc_204, uc_205, uc_206, uc_207, uc_208, 
    uc_209, uc_210, uc_211, uc_212, uc_213, uc_214, uc_215, uc_216, uc_217, uc_218, 
    \normalizedWires[1655] , \normalizedWires[1654] , \normalizedWires[1653] , \normalizedWires[1652] , 
    \normalizedWires[1651] , \normalizedWires[1650] , \normalizedWires[1649] , \normalizedWires[1648] , 
    \normalizedWires[1647] , \normalizedWires[1646] , \normalizedWires[1645] , \normalizedWires[1644] , 
    \normalizedWires[1643] , \normalizedWires[1642] , \normalizedWires[1641] , \normalizedWires[1640] , 
    \normalizedWires[1639] , \normalizedWires[1638] , \normalizedWires[1637] , \normalizedWires[1636] , 
    \normalizedWires[1635] , \normalizedWires[1634] , \normalizedWires[1633] , \normalizedWires[1632] , 
    \normalizedWires[1631] , \normalizedWires[1630] , \normalizedWires[1629] , \normalizedWires[1628] , 
    \normalizedWires[1627] , \normalizedWires[1626] , \normalizedWires[1625] , uc_219, 
    uc_220, uc_221, uc_222, uc_223, uc_224, uc_225, uc_226, uc_227, uc_228, uc_229, 
    uc_230, uc_231, uc_232, uc_233, uc_234, uc_235, uc_236, uc_237, uc_238, uc_239, 
    uc_240, uc_241, uc_242, uc_243, uc_244, uc_245, uc_246, uc_247, uc_248, uc_249, 
    uc_250, uc_251, uc_252, \normalizedWires[1590] , \normalizedWires[1589] , \normalizedWires[1588] , 
    \normalizedWires[1587] , \normalizedWires[1586] , \normalizedWires[1585] , \normalizedWires[1584] , 
    \normalizedWires[1583] , \normalizedWires[1582] , \normalizedWires[1581] , \normalizedWires[1580] , 
    \normalizedWires[1579] , \normalizedWires[1578] , \normalizedWires[1577] , \normalizedWires[1576] , 
    \normalizedWires[1575] , \normalizedWires[1574] , \normalizedWires[1573] , \normalizedWires[1572] , 
    \normalizedWires[1571] , \normalizedWires[1570] , \normalizedWires[1569] , \normalizedWires[1568] , 
    \normalizedWires[1567] , \normalizedWires[1566] , \normalizedWires[1565] , \normalizedWires[1564] , 
    \normalizedWires[1563] , \normalizedWires[1562] , \normalizedWires[1561] , \normalizedWires[1560] , 
    uc_253, uc_254, uc_255, uc_256, uc_257, uc_258, uc_259, uc_260, uc_261, uc_262, 
    uc_263, uc_264, uc_265, uc_266, uc_267, uc_268, uc_269, uc_270, uc_271, uc_272, 
    uc_273, uc_274, uc_275, uc_276, uc_277, uc_278, uc_279, uc_280, uc_281, uc_282, 
    uc_283, uc_284, uc_285, uc_286, \normalizedWires[1525] , \normalizedWires[1524] , 
    \normalizedWires[1523] , \normalizedWires[1522] , \normalizedWires[1521] , \normalizedWires[1520] , 
    \normalizedWires[1519] , \normalizedWires[1518] , \normalizedWires[1517] , \normalizedWires[1516] , 
    \normalizedWires[1515] , \normalizedWires[1514] , \normalizedWires[1513] , \normalizedWires[1512] , 
    \normalizedWires[1511] , \normalizedWires[1510] , \normalizedWires[1509] , \normalizedWires[1508] , 
    \normalizedWires[1507] , \normalizedWires[1506] , \normalizedWires[1505] , \normalizedWires[1504] , 
    \normalizedWires[1503] , \normalizedWires[1502] , \normalizedWires[1501] , \normalizedWires[1500] , 
    \normalizedWires[1499] , \normalizedWires[1498] , \normalizedWires[1497] , \normalizedWires[1496] , 
    \normalizedWires[1495] , uc_287, uc_288, uc_289, uc_290, uc_291, uc_292, uc_293, 
    uc_294, uc_295, uc_296, uc_297, uc_298, uc_299, uc_300, uc_301, uc_302, uc_303, 
    uc_304, uc_305, uc_306, uc_307, uc_308, uc_309, uc_310, uc_311, uc_312, uc_313, 
    uc_314, uc_315, uc_316, uc_317, uc_318, uc_319, uc_320, \normalizedWires[1460] , 
    \normalizedWires[1459] , \normalizedWires[1458] , \normalizedWires[1457] , \normalizedWires[1456] , 
    \normalizedWires[1455] , \normalizedWires[1454] , \normalizedWires[1453] , \normalizedWires[1452] , 
    \normalizedWires[1451] , \normalizedWires[1450] , \normalizedWires[1449] , \normalizedWires[1448] , 
    \normalizedWires[1447] , \normalizedWires[1446] , \normalizedWires[1445] , \normalizedWires[1444] , 
    \normalizedWires[1443] , \normalizedWires[1442] , \normalizedWires[1441] , \normalizedWires[1440] , 
    \normalizedWires[1439] , \normalizedWires[1438] , \normalizedWires[1437] , \normalizedWires[1436] , 
    \normalizedWires[1435] , \normalizedWires[1434] , \normalizedWires[1433] , \normalizedWires[1432] , 
    \normalizedWires[1431] , \normalizedWires[1430] , uc_321, uc_322, uc_323, uc_324, 
    uc_325, uc_326, uc_327, uc_328, uc_329, uc_330, uc_331, uc_332, uc_333, uc_334, 
    uc_335, uc_336, uc_337, uc_338, uc_339, uc_340, uc_341, uc_342, uc_343, uc_344, 
    uc_345, uc_346, uc_347, uc_348, uc_349, uc_350, uc_351, uc_352, uc_353, uc_354, 
    \normalizedWires[1395] , \normalizedWires[1394] , \normalizedWires[1393] , \normalizedWires[1392] , 
    \normalizedWires[1391] , \normalizedWires[1390] , \normalizedWires[1389] , \normalizedWires[1388] , 
    \normalizedWires[1387] , \normalizedWires[1386] , \normalizedWires[1385] , \normalizedWires[1384] , 
    \normalizedWires[1383] , \normalizedWires[1382] , \normalizedWires[1381] , \normalizedWires[1380] , 
    \normalizedWires[1379] , \normalizedWires[1378] , \normalizedWires[1377] , \normalizedWires[1376] , 
    \normalizedWires[1375] , \normalizedWires[1374] , \normalizedWires[1373] , \normalizedWires[1372] , 
    \normalizedWires[1371] , \normalizedWires[1370] , \normalizedWires[1369] , \normalizedWires[1368] , 
    \normalizedWires[1367] , \normalizedWires[1366] , \normalizedWires[1365] , uc_355, 
    uc_356, uc_357, uc_358, uc_359, uc_360, uc_361, uc_362, uc_363, uc_364, uc_365, 
    uc_366, uc_367, uc_368, uc_369, uc_370, uc_371, uc_372, uc_373, uc_374, uc_375, 
    uc_376, uc_377, uc_378, uc_379, uc_380, uc_381, uc_382, uc_383, uc_384, uc_385, 
    uc_386, uc_387, uc_388, \normalizedWires[1330] , \normalizedWires[1329] , \normalizedWires[1328] , 
    \normalizedWires[1327] , \normalizedWires[1326] , \normalizedWires[1325] , \normalizedWires[1324] , 
    \normalizedWires[1323] , \normalizedWires[1322] , \normalizedWires[1321] , \normalizedWires[1320] , 
    \normalizedWires[1319] , \normalizedWires[1318] , \normalizedWires[1317] , \normalizedWires[1316] , 
    \normalizedWires[1315] , \normalizedWires[1314] , \normalizedWires[1313] , \normalizedWires[1312] , 
    \normalizedWires[1311] , \normalizedWires[1310] , \normalizedWires[1309] , \normalizedWires[1308] , 
    \normalizedWires[1307] , \normalizedWires[1306] , \normalizedWires[1305] , \normalizedWires[1304] , 
    \normalizedWires[1303] , \normalizedWires[1302] , \normalizedWires[1301] , \normalizedWires[1300] , 
    uc_389, uc_390, uc_391, uc_392, uc_393, uc_394, uc_395, uc_396, uc_397, uc_398, 
    uc_399, uc_400, uc_401, uc_402, uc_403, uc_404, uc_405, uc_406, uc_407, uc_408, 
    uc_409, uc_410, uc_411, uc_412, uc_413, uc_414, uc_415, uc_416, uc_417, uc_418, 
    uc_419, uc_420, uc_421, uc_422, \normalizedWires[1265] , \normalizedWires[1264] , 
    \normalizedWires[1263] , \normalizedWires[1262] , \normalizedWires[1261] , \normalizedWires[1260] , 
    \normalizedWires[1259] , \normalizedWires[1258] , \normalizedWires[1257] , \normalizedWires[1256] , 
    \normalizedWires[1255] , \normalizedWires[1254] , \normalizedWires[1253] , \normalizedWires[1252] , 
    \normalizedWires[1251] , \normalizedWires[1250] , \normalizedWires[1249] , \normalizedWires[1248] , 
    \normalizedWires[1247] , \normalizedWires[1246] , \normalizedWires[1245] , \normalizedWires[1244] , 
    \normalizedWires[1243] , \normalizedWires[1242] , \normalizedWires[1241] , \normalizedWires[1240] , 
    \normalizedWires[1239] , \normalizedWires[1238] , \normalizedWires[1237] , \normalizedWires[1236] , 
    \normalizedWires[1235] , uc_423, uc_424, uc_425, uc_426, uc_427, uc_428, uc_429, 
    uc_430, uc_431, uc_432, uc_433, uc_434, uc_435, uc_436, uc_437, uc_438, uc_439, 
    uc_440, uc_441, uc_442, uc_443, uc_444, uc_445, uc_446, uc_447, uc_448, uc_449, 
    uc_450, uc_451, uc_452, uc_453, uc_454, uc_455, uc_456, \normalizedWires[1200] , 
    \normalizedWires[1199] , \normalizedWires[1198] , \normalizedWires[1197] , \normalizedWires[1196] , 
    \normalizedWires[1195] , \normalizedWires[1194] , \normalizedWires[1193] , \normalizedWires[1192] , 
    \normalizedWires[1191] , \normalizedWires[1190] , \normalizedWires[1189] , \normalizedWires[1188] , 
    \normalizedWires[1187] , \normalizedWires[1186] , \normalizedWires[1185] , \normalizedWires[1184] , 
    \normalizedWires[1183] , \normalizedWires[1182] , \normalizedWires[1181] , \normalizedWires[1180] , 
    \normalizedWires[1179] , \normalizedWires[1178] , \normalizedWires[1177] , \normalizedWires[1176] , 
    \normalizedWires[1175] , \normalizedWires[1174] , \normalizedWires[1173] , \normalizedWires[1172] , 
    \normalizedWires[1171] , \normalizedWires[1170] , uc_457, uc_458, uc_459, uc_460, 
    uc_461, uc_462, uc_463, uc_464, uc_465, uc_466, uc_467, uc_468, uc_469, uc_470, 
    uc_471, uc_472, uc_473, uc_474, uc_475, uc_476, uc_477, uc_478, uc_479, uc_480, 
    uc_481, uc_482, uc_483, uc_484, uc_485, uc_486, uc_487, uc_488, uc_489, uc_490, 
    \normalizedWires[1135] , \normalizedWires[1134] , \normalizedWires[1133] , \normalizedWires[1132] , 
    \normalizedWires[1131] , \normalizedWires[1130] , \normalizedWires[1129] , \normalizedWires[1128] , 
    \normalizedWires[1127] , \normalizedWires[1126] , \normalizedWires[1125] , \normalizedWires[1124] , 
    \normalizedWires[1123] , \normalizedWires[1122] , \normalizedWires[1121] , \normalizedWires[1120] , 
    \normalizedWires[1119] , \normalizedWires[1118] , \normalizedWires[1117] , \normalizedWires[1116] , 
    \normalizedWires[1115] , \normalizedWires[1114] , \normalizedWires[1113] , \normalizedWires[1112] , 
    \normalizedWires[1111] , \normalizedWires[1110] , \normalizedWires[1109] , \normalizedWires[1108] , 
    \normalizedWires[1107] , \normalizedWires[1106] , \normalizedWires[1105] , uc_491, 
    uc_492, uc_493, uc_494, uc_495, uc_496, uc_497, uc_498, uc_499, uc_500, uc_501, 
    uc_502, uc_503, uc_504, uc_505, uc_506, uc_507, uc_508, uc_509, uc_510, uc_511, 
    uc_512, uc_513, uc_514, uc_515, uc_516, uc_517, uc_518, uc_519, uc_520, uc_521, 
    uc_522, uc_523, uc_524, \normalizedWires[1070] , \normalizedWires[1069] , \normalizedWires[1068] , 
    \normalizedWires[1067] , \normalizedWires[1066] , \normalizedWires[1065] , \normalizedWires[1064] , 
    \normalizedWires[1063] , \normalizedWires[1062] , \normalizedWires[1061] , \normalizedWires[1060] , 
    \normalizedWires[1059] , \normalizedWires[1058] , \normalizedWires[1057] , \normalizedWires[1056] , 
    \normalizedWires[1055] , \normalizedWires[1054] , \normalizedWires[1053] , \normalizedWires[1052] , 
    \normalizedWires[1051] , \normalizedWires[1050] , \normalizedWires[1049] , \normalizedWires[1048] , 
    \normalizedWires[1047] , \normalizedWires[1046] , \normalizedWires[1045] , \normalizedWires[1044] , 
    \normalizedWires[1043] , \normalizedWires[1042] , \normalizedWires[1041] , \normalizedWires[1040] , 
    uc_525, uc_526, uc_527, uc_528, uc_529, uc_530, uc_531, uc_532, uc_533, uc_534, 
    uc_535, uc_536, uc_537, uc_538, uc_539, uc_540, uc_541, uc_542, uc_543, uc_544, 
    uc_545, uc_546, uc_547, uc_548, uc_549, uc_550, uc_551, uc_552, uc_553, uc_554, 
    uc_555, uc_556, uc_557, uc_558, \normalizedWires[1005] , \normalizedWires[1004] , 
    \normalizedWires[1003] , \normalizedWires[1002] , \normalizedWires[1001] , \normalizedWires[1000] , 
    \normalizedWires[999] , \normalizedWires[998] , \normalizedWires[997] , \normalizedWires[996] , 
    \normalizedWires[995] , \normalizedWires[994] , \normalizedWires[993] , \normalizedWires[992] , 
    \normalizedWires[991] , \normalizedWires[990] , \normalizedWires[989] , \normalizedWires[988] , 
    \normalizedWires[987] , \normalizedWires[986] , \normalizedWires[985] , \normalizedWires[984] , 
    \normalizedWires[983] , \normalizedWires[982] , \normalizedWires[981] , \normalizedWires[980] , 
    \normalizedWires[979] , \normalizedWires[978] , \normalizedWires[977] , \normalizedWires[976] , 
    \normalizedWires[975] , uc_559, uc_560, uc_561, uc_562, uc_563, uc_564, uc_565, 
    uc_566, uc_567, uc_568, uc_569, uc_570, uc_571, uc_572, uc_573, uc_574, uc_575, 
    uc_576, uc_577, uc_578, uc_579, uc_580, uc_581, uc_582, uc_583, uc_584, uc_585, 
    uc_586, uc_587, uc_588, uc_589, uc_590, uc_591, uc_592, \normalizedWires[940] , 
    \normalizedWires[939] , \normalizedWires[938] , \normalizedWires[937] , \normalizedWires[936] , 
    \normalizedWires[935] , \normalizedWires[934] , \normalizedWires[933] , \normalizedWires[932] , 
    \normalizedWires[931] , \normalizedWires[930] , \normalizedWires[929] , \normalizedWires[928] , 
    \normalizedWires[927] , \normalizedWires[926] , \normalizedWires[925] , \normalizedWires[924] , 
    \normalizedWires[923] , \normalizedWires[922] , \normalizedWires[921] , \normalizedWires[920] , 
    \normalizedWires[919] , \normalizedWires[918] , \normalizedWires[917] , \normalizedWires[916] , 
    \normalizedWires[915] , \normalizedWires[914] , \normalizedWires[913] , \normalizedWires[912] , 
    \normalizedWires[911] , \normalizedWires[910] , uc_593, uc_594, uc_595, uc_596, 
    uc_597, uc_598, uc_599, uc_600, uc_601, uc_602, uc_603, uc_604, uc_605, uc_606, 
    uc_607, uc_608, uc_609, uc_610, uc_611, uc_612, uc_613, uc_614, uc_615, uc_616, 
    uc_617, uc_618, uc_619, uc_620, uc_621, uc_622, uc_623, uc_624, uc_625, uc_626, 
    \normalizedWires[875] , \normalizedWires[874] , \normalizedWires[873] , \normalizedWires[872] , 
    \normalizedWires[871] , \normalizedWires[870] , \normalizedWires[869] , \normalizedWires[868] , 
    \normalizedWires[867] , \normalizedWires[866] , \normalizedWires[865] , \normalizedWires[864] , 
    \normalizedWires[863] , \normalizedWires[862] , \normalizedWires[861] , \normalizedWires[860] , 
    \normalizedWires[859] , \normalizedWires[858] , \normalizedWires[857] , \normalizedWires[856] , 
    \normalizedWires[855] , \normalizedWires[854] , \normalizedWires[853] , \normalizedWires[852] , 
    \normalizedWires[851] , \normalizedWires[850] , \normalizedWires[849] , \normalizedWires[848] , 
    \normalizedWires[847] , \normalizedWires[846] , \normalizedWires[845] , uc_627, 
    uc_628, uc_629, uc_630, uc_631, uc_632, uc_633, uc_634, uc_635, uc_636, uc_637, 
    uc_638, uc_639, uc_640, uc_641, uc_642, uc_643, uc_644, uc_645, uc_646, uc_647, 
    uc_648, uc_649, uc_650, uc_651, uc_652, uc_653, uc_654, uc_655, uc_656, uc_657, 
    uc_658, uc_659, uc_660, \normalizedWires[810] , \normalizedWires[809] , \normalizedWires[808] , 
    \normalizedWires[807] , \normalizedWires[806] , \normalizedWires[805] , \normalizedWires[804] , 
    \normalizedWires[803] , \normalizedWires[802] , \normalizedWires[801] , \normalizedWires[800] , 
    \normalizedWires[799] , \normalizedWires[798] , \normalizedWires[797] , \normalizedWires[796] , 
    \normalizedWires[795] , \normalizedWires[794] , \normalizedWires[793] , \normalizedWires[792] , 
    \normalizedWires[791] , \normalizedWires[790] , \normalizedWires[789] , \normalizedWires[788] , 
    \normalizedWires[787] , \normalizedWires[786] , \normalizedWires[785] , \normalizedWires[784] , 
    \normalizedWires[783] , \normalizedWires[782] , \normalizedWires[781] , \normalizedWires[780] , 
    uc_661, uc_662, uc_663, uc_664, uc_665, uc_666, uc_667, uc_668, uc_669, uc_670, 
    uc_671, uc_672, uc_673, uc_674, uc_675, uc_676, uc_677, uc_678, uc_679, uc_680, 
    uc_681, uc_682, uc_683, uc_684, uc_685, uc_686, uc_687, uc_688, uc_689, uc_690, 
    uc_691, uc_692, uc_693, uc_694, \normalizedWires[745] , \normalizedWires[744] , 
    \normalizedWires[743] , \normalizedWires[742] , \normalizedWires[741] , \normalizedWires[740] , 
    \normalizedWires[739] , \normalizedWires[738] , \normalizedWires[737] , \normalizedWires[736] , 
    \normalizedWires[735] , \normalizedWires[734] , \normalizedWires[733] , \normalizedWires[732] , 
    \normalizedWires[731] , \normalizedWires[730] , \normalizedWires[729] , \normalizedWires[728] , 
    \normalizedWires[727] , \normalizedWires[726] , \normalizedWires[725] , \normalizedWires[724] , 
    \normalizedWires[723] , \normalizedWires[722] , \normalizedWires[721] , \normalizedWires[720] , 
    \normalizedWires[719] , \normalizedWires[718] , \normalizedWires[717] , \normalizedWires[716] , 
    \normalizedWires[715] , uc_695, uc_696, uc_697, uc_698, uc_699, uc_700, uc_701, 
    uc_702, uc_703, uc_704, uc_705, uc_706, uc_707, uc_708, uc_709, uc_710, uc_711, 
    uc_712, uc_713, uc_714, uc_715, uc_716, uc_717, uc_718, uc_719, uc_720, uc_721, 
    uc_722, uc_723, uc_724, uc_725, uc_726, uc_727, uc_728, \normalizedWires[680] , 
    \normalizedWires[679] , \normalizedWires[678] , \normalizedWires[677] , \normalizedWires[676] , 
    \normalizedWires[675] , \normalizedWires[674] , \normalizedWires[673] , \normalizedWires[672] , 
    \normalizedWires[671] , \normalizedWires[670] , \normalizedWires[669] , \normalizedWires[668] , 
    \normalizedWires[667] , \normalizedWires[666] , \normalizedWires[665] , \normalizedWires[664] , 
    \normalizedWires[663] , \normalizedWires[662] , \normalizedWires[661] , \normalizedWires[660] , 
    \normalizedWires[659] , \normalizedWires[658] , \normalizedWires[657] , \normalizedWires[656] , 
    \normalizedWires[655] , \normalizedWires[654] , \normalizedWires[653] , \normalizedWires[652] , 
    \normalizedWires[651] , \normalizedWires[650] , uc_729, uc_730, uc_731, uc_732, 
    uc_733, uc_734, uc_735, uc_736, uc_737, uc_738, uc_739, uc_740, uc_741, uc_742, 
    uc_743, uc_744, uc_745, uc_746, uc_747, uc_748, uc_749, uc_750, uc_751, uc_752, 
    uc_753, uc_754, uc_755, uc_756, uc_757, uc_758, uc_759, uc_760, uc_761, uc_762, 
    \normalizedWires[615] , \normalizedWires[614] , \normalizedWires[613] , \normalizedWires[612] , 
    \normalizedWires[611] , \normalizedWires[610] , \normalizedWires[609] , \normalizedWires[608] , 
    \normalizedWires[607] , \normalizedWires[606] , \normalizedWires[605] , \normalizedWires[604] , 
    \normalizedWires[603] , \normalizedWires[602] , \normalizedWires[601] , \normalizedWires[600] , 
    \normalizedWires[599] , \normalizedWires[598] , \normalizedWires[597] , \normalizedWires[596] , 
    \normalizedWires[595] , \normalizedWires[594] , \normalizedWires[593] , \normalizedWires[592] , 
    \normalizedWires[591] , \normalizedWires[590] , \normalizedWires[589] , \normalizedWires[588] , 
    \normalizedWires[587] , \normalizedWires[586] , \normalizedWires[585] , uc_763, 
    uc_764, uc_765, uc_766, uc_767, uc_768, uc_769, uc_770, uc_771, uc_772, uc_773, 
    uc_774, uc_775, uc_776, uc_777, uc_778, uc_779, uc_780, uc_781, uc_782, uc_783, 
    uc_784, uc_785, uc_786, uc_787, uc_788, uc_789, uc_790, uc_791, uc_792, uc_793, 
    uc_794, uc_795, uc_796, \normalizedWires[550] , \normalizedWires[549] , \normalizedWires[548] , 
    \normalizedWires[547] , \normalizedWires[546] , \normalizedWires[545] , \normalizedWires[544] , 
    \normalizedWires[543] , \normalizedWires[542] , \normalizedWires[541] , \normalizedWires[540] , 
    \normalizedWires[539] , \normalizedWires[538] , \normalizedWires[537] , \normalizedWires[536] , 
    \normalizedWires[535] , \normalizedWires[534] , \normalizedWires[533] , \normalizedWires[532] , 
    \normalizedWires[531] , \normalizedWires[530] , \normalizedWires[529] , \normalizedWires[528] , 
    \normalizedWires[527] , \normalizedWires[526] , \normalizedWires[525] , \normalizedWires[524] , 
    \normalizedWires[523] , \normalizedWires[522] , \normalizedWires[521] , \normalizedWires[520] , 
    uc_797, uc_798, uc_799, uc_800, uc_801, uc_802, uc_803, uc_804, uc_805, uc_806, 
    uc_807, uc_808, uc_809, uc_810, uc_811, uc_812, uc_813, uc_814, uc_815, uc_816, 
    uc_817, uc_818, uc_819, uc_820, uc_821, uc_822, uc_823, uc_824, uc_825, uc_826, 
    uc_827, uc_828, uc_829, uc_830, \normalizedWires[485] , \normalizedWires[484] , 
    \normalizedWires[483] , \normalizedWires[482] , \normalizedWires[481] , \normalizedWires[480] , 
    \normalizedWires[479] , \normalizedWires[478] , \normalizedWires[477] , \normalizedWires[476] , 
    \normalizedWires[475] , \normalizedWires[474] , \normalizedWires[473] , \normalizedWires[472] , 
    \normalizedWires[471] , \normalizedWires[470] , \normalizedWires[469] , \normalizedWires[468] , 
    \normalizedWires[467] , \normalizedWires[466] , \normalizedWires[465] , \normalizedWires[464] , 
    \normalizedWires[463] , \normalizedWires[462] , \normalizedWires[461] , \normalizedWires[460] , 
    \normalizedWires[459] , \normalizedWires[458] , \normalizedWires[457] , \normalizedWires[456] , 
    \normalizedWires[455] , uc_831, uc_832, uc_833, uc_834, uc_835, uc_836, uc_837, 
    uc_838, uc_839, uc_840, uc_841, uc_842, uc_843, uc_844, uc_845, uc_846, uc_847, 
    uc_848, uc_849, uc_850, uc_851, uc_852, uc_853, uc_854, uc_855, uc_856, uc_857, 
    uc_858, uc_859, uc_860, uc_861, uc_862, uc_863, uc_864, \normalizedWires[420] , 
    \normalizedWires[419] , \normalizedWires[418] , \normalizedWires[417] , \normalizedWires[416] , 
    \normalizedWires[415] , \normalizedWires[414] , \normalizedWires[413] , \normalizedWires[412] , 
    \normalizedWires[411] , \normalizedWires[410] , \normalizedWires[409] , \normalizedWires[408] , 
    \normalizedWires[407] , \normalizedWires[406] , \normalizedWires[405] , \normalizedWires[404] , 
    \normalizedWires[403] , \normalizedWires[402] , \normalizedWires[401] , \normalizedWires[400] , 
    \normalizedWires[399] , \normalizedWires[398] , \normalizedWires[397] , \normalizedWires[396] , 
    \normalizedWires[395] , \normalizedWires[394] , \normalizedWires[393] , \normalizedWires[392] , 
    \normalizedWires[391] , \normalizedWires[390] , uc_865, uc_866, uc_867, uc_868, 
    uc_869, uc_870, uc_871, uc_872, uc_873, uc_874, uc_875, uc_876, uc_877, uc_878, 
    uc_879, uc_880, uc_881, uc_882, uc_883, uc_884, uc_885, uc_886, uc_887, uc_888, 
    uc_889, uc_890, uc_891, uc_892, uc_893, uc_894, uc_895, uc_896, uc_897, uc_898, 
    \normalizedWires[355] , \normalizedWires[354] , \normalizedWires[353] , \normalizedWires[352] , 
    \normalizedWires[351] , \normalizedWires[350] , \normalizedWires[349] , \normalizedWires[348] , 
    \normalizedWires[347] , \normalizedWires[346] , \normalizedWires[345] , \normalizedWires[344] , 
    \normalizedWires[343] , \normalizedWires[342] , \normalizedWires[341] , \normalizedWires[340] , 
    \normalizedWires[339] , \normalizedWires[338] , \normalizedWires[337] , \normalizedWires[336] , 
    \normalizedWires[335] , \normalizedWires[334] , \normalizedWires[333] , \normalizedWires[332] , 
    \normalizedWires[331] , \normalizedWires[330] , \normalizedWires[329] , \normalizedWires[328] , 
    \normalizedWires[327] , \normalizedWires[326] , \normalizedWires[325] , uc_899, 
    uc_900, uc_901, uc_902, uc_903, uc_904, uc_905, uc_906, uc_907, uc_908, uc_909, 
    uc_910, uc_911, uc_912, uc_913, uc_914, uc_915, uc_916, uc_917, uc_918, uc_919, 
    uc_920, uc_921, uc_922, uc_923, uc_924, uc_925, uc_926, uc_927, uc_928, uc_929, 
    uc_930, uc_931, uc_932, \normalizedWires[290] , \normalizedWires[289] , \normalizedWires[288] , 
    \normalizedWires[287] , \normalizedWires[286] , \normalizedWires[285] , \normalizedWires[284] , 
    \normalizedWires[283] , \normalizedWires[282] , \normalizedWires[281] , \normalizedWires[280] , 
    \normalizedWires[279] , \normalizedWires[278] , \normalizedWires[277] , \normalizedWires[276] , 
    \normalizedWires[275] , \normalizedWires[274] , \normalizedWires[273] , \normalizedWires[272] , 
    \normalizedWires[271] , \normalizedWires[270] , \normalizedWires[269] , \normalizedWires[268] , 
    \normalizedWires[267] , \normalizedWires[266] , \normalizedWires[265] , \normalizedWires[264] , 
    \normalizedWires[263] , \normalizedWires[262] , \normalizedWires[261] , \normalizedWires[260] , 
    uc_933, uc_934, uc_935, uc_936, uc_937, uc_938, uc_939, uc_940, uc_941, uc_942, 
    uc_943, uc_944, uc_945, uc_946, uc_947, uc_948, uc_949, uc_950, uc_951, uc_952, 
    uc_953, uc_954, uc_955, uc_956, uc_957, uc_958, uc_959, uc_960, uc_961, uc_962, 
    uc_963, uc_964, uc_965, uc_966, \normalizedWires[225] , \normalizedWires[224] , 
    \normalizedWires[223] , \normalizedWires[222] , \normalizedWires[221] , \normalizedWires[220] , 
    \normalizedWires[219] , \normalizedWires[218] , \normalizedWires[217] , \normalizedWires[216] , 
    \normalizedWires[215] , \normalizedWires[214] , \normalizedWires[213] , \normalizedWires[212] , 
    \normalizedWires[211] , \normalizedWires[210] , \normalizedWires[209] , \normalizedWires[208] , 
    \normalizedWires[207] , \normalizedWires[206] , \normalizedWires[205] , \normalizedWires[204] , 
    \normalizedWires[203] , \normalizedWires[202] , \normalizedWires[201] , \normalizedWires[200] , 
    \normalizedWires[199] , \normalizedWires[198] , \normalizedWires[197] , \normalizedWires[196] , 
    \normalizedWires[195] , uc_967, uc_968, uc_969, uc_970, uc_971, uc_972, uc_973, 
    uc_974, uc_975, uc_976, uc_977, uc_978, uc_979, uc_980, uc_981, uc_982, uc_983, 
    uc_984, uc_985, uc_986, uc_987, uc_988, uc_989, uc_990, uc_991, uc_992, uc_993, 
    uc_994, uc_995, uc_996, uc_997, uc_998, uc_999, uc_1000, \normalizedWires[160] , 
    \normalizedWires[159] , \normalizedWires[158] , \normalizedWires[157] , \normalizedWires[156] , 
    \normalizedWires[155] , \normalizedWires[154] , \normalizedWires[153] , \normalizedWires[152] , 
    \normalizedWires[151] , \normalizedWires[150] , \normalizedWires[149] , \normalizedWires[148] , 
    \normalizedWires[147] , \normalizedWires[146] , \normalizedWires[145] , \normalizedWires[144] , 
    \normalizedWires[143] , \normalizedWires[142] , \normalizedWires[141] , \normalizedWires[140] , 
    \normalizedWires[139] , \normalizedWires[138] , \normalizedWires[137] , \normalizedWires[136] , 
    \normalizedWires[135] , \normalizedWires[134] , \normalizedWires[133] , \normalizedWires[132] , 
    \normalizedWires[131] , \normalizedWires[130] , uc_1001, uc_1002, uc_1003, uc_1004, 
    uc_1005, uc_1006, uc_1007, uc_1008, uc_1009, uc_1010, uc_1011, uc_1012, uc_1013, 
    uc_1014, uc_1015, uc_1016, uc_1017, uc_1018, uc_1019, uc_1020, uc_1021, uc_1022, 
    uc_1023, uc_1024, uc_1025, uc_1026, uc_1027, uc_1028, uc_1029, uc_1030, uc_1031, 
    uc_1032, uc_1033, uc_1034, \normalizedWires[95] , \normalizedWires[94] , \normalizedWires[93] , 
    \normalizedWires[92] , \normalizedWires[91] , \normalizedWires[90] , \normalizedWires[89] , 
    \normalizedWires[88] , \normalizedWires[87] , \normalizedWires[86] , \normalizedWires[85] , 
    \normalizedWires[84] , \normalizedWires[83] , \normalizedWires[82] , \normalizedWires[81] , 
    \normalizedWires[80] , \normalizedWires[79] , \normalizedWires[78] , \normalizedWires[77] , 
    \normalizedWires[76] , \normalizedWires[75] , \normalizedWires[74] , \normalizedWires[73] , 
    \normalizedWires[72] , \normalizedWires[71] , \normalizedWires[70] , \normalizedWires[69] , 
    \normalizedWires[68] , \normalizedWires[67] , \normalizedWires[66] , \normalizedWires[65] , 
    uc_1035, uc_1036, uc_1037, uc_1038, uc_1039, uc_1040, uc_1041, uc_1042, uc_1043, 
    uc_1044, uc_1045, uc_1046, uc_1047, uc_1048, uc_1049, uc_1050, uc_1051, uc_1052, 
    uc_1053, uc_1054, uc_1055, uc_1056, uc_1057, uc_1058, uc_1059, uc_1060, uc_1061, 
    uc_1062, uc_1063, uc_1064, uc_1065, uc_1066, uc_1067, uc_1068, \normalizedWires[30] , 
    \normalizedWires[29] , \normalizedWires[28] , \normalizedWires[27] , \normalizedWires[26] , 
    \normalizedWires[25] , \normalizedWires[24] , \normalizedWires[23] , \normalizedWires[22] , 
    \normalizedWires[21] , \normalizedWires[20] , \normalizedWires[19] , \normalizedWires[18] , 
    \normalizedWires[17] , \normalizedWires[16] , \normalizedWires[15] , \normalizedWires[14] , 
    \normalizedWires[13] , \normalizedWires[12] , \normalizedWires[11] , \normalizedWires[10] , 
    \normalizedWires[9] , \normalizedWires[8] , \normalizedWires[7] , \normalizedWires[6] , 
    \normalizedWires[5] , \normalizedWires[4] , \normalizedWires[3] , \normalizedWires[2] , 
    \normalizedWires[1] , uc_1069}));
INV_X1 slo__sro_c1238 (.ZN (slo__sro_n1029), .A (drc_ipo_n26));
NOR2_X1 CLOCK_sgo__sro_c2229 (.ZN (CLOCK_sgo__sro_n1964), .A1 (\Res_imm[43] ), .A2 (\Res_imm[46] ));
BUF_X8 hfn_ipo_c25 (.Z (hfn_ipo_n25), .A (CLOCK_slo__sro_n2662));
BUF_X32 drc_ipo_c26 (.Z (drc_ipo_n26), .A (A_in));
NOR2_X1 sgo__sro_c39 (.ZN (sgo__sro_n34), .A1 (sgo__sro_n35), .A2 (slo__n881));
AOI21_X2 sgo__sro_c40 (.ZN (n_0_1_6), .A (sgo__sro_n34), .B1 (opt_ipo_n1555), .B2 (opt_ipo_n1344));
BUF_X8 sgo__c28 (.Z (opt_ipo_n1380), .A (sgo__n28));
BUF_X16 drc_ipo_c27 (.Z (drc_ipo_n27), .A (B_in));
NOR3_X1 sgo__sro_c333 (.ZN (n_0_1_28), .A1 (sgo__sro_n246), .A2 (\Res_imm[36] ), .A3 (\Res_imm[39] ));
NOR2_X4 sgo__sro_c62 (.ZN (sgo__sro_n53), .A1 (n_0_1_69), .A2 (n_0_1_19));
NAND2_X1 slo__sro_c547 (.ZN (slo__sro_n406), .A1 (n_0_98), .A2 (slo__sro_n408));
NOR2_X4 sgo__sro_c64 (.ZN (sgo__sro_n51), .A1 (slo__mro_n391), .A2 (n_0_1_75));
AND2_X1 sgo__sro_c200 (.ZN (sgo__sro_n146), .A1 (n_0_1_74), .A2 (n_0_1_73));
AND2_X1 sgo__sro_c201 (.ZN (sgo__sro_n145), .A1 (n_0_1_70), .A2 (sgo__sro_n146));
NAND2_X2 slo__sro_c546 (.ZN (slo__sro_n407), .A1 (n_0_147), .A2 (drc_ipo_n26));
INV_X4 slo__xsl_c417 (.ZN (slo__xsl_n298), .A (CLOCK_slo__sro_n2662));
AND2_X2 sgo__sro_c178 (.ZN (sgo__sro_n130), .A1 (n_0_1_144), .A2 (n_0_1_143));
NAND3_X2 sgo__sro_c179 (.ZN (n_0_1_75), .A1 (sgo__sro_n130), .A2 (n_0_1_76), .A3 (n_0_1_142));
INV_X1 slo__sro_c521 (.ZN (slo__sro_n384), .A (drc_ipo_n26));
NAND2_X2 slo__sro_c522 (.ZN (slo__sro_n383), .A1 (n_0_141), .A2 (drc_ipo_n26));
NAND2_X1 slo__sro_c523 (.ZN (slo__sro_n382), .A1 (n_0_104), .A2 (slo__sro_n384));
NAND2_X4 slo__sro_c524 (.ZN (slo__sro_n381), .A1 (slo__sro_n383), .A2 (slo__sro_n382));
NOR4_X4 slo__mro_c532 (.ZN (slo__mro_n393), .A1 (\Res_imm[58] ), .A2 (\Res_imm[60] )
    , .A3 (\Res_imm[57] ), .A4 (\Res_imm[63] ));
AND2_X4 slo__mro_c533 (.ZN (slo__mro_n392), .A1 (n_0_1_26), .A2 (slo__mro_n393));
NAND3_X4 slo__mro_c534 (.ZN (slo__mro_n391), .A1 (slo__mro_n392), .A2 (slo__mro_n394), .A3 (sgo__sro_n53));
NAND2_X4 slo__sro_c548 (.ZN (slo__sro_n405), .A1 (slo__sro_n407), .A2 (slo__sro_n406));
NAND2_X1 slo__sro_c564 (.ZN (slo__sro_n422), .A1 (n_0_162), .A2 (drc_ipo_n27));
NAND2_X1 slo__sro_c565 (.ZN (slo__sro_n421), .A1 (n_0_83), .A2 (slo__sro_n423));
NAND2_X4 slo__sro_c566 (.ZN (slo__sro_n420), .A1 (slo__sro_n422), .A2 (slo__sro_n421));
NAND2_X2 slo__sro_c674 (.ZN (slo__sro_n515), .A1 (n_0_174), .A2 (drc_ipo_n27));
NAND2_X4 CLOCK_slo__mro_c2662 (.ZN (CLOCK_slo__mro_n2310), .A1 (slo__sro_n1000), .A2 (slo__sro_n999));
INV_X1 CLOCK_sgo__sro_c2231 (.ZN (n_0_1_68), .A (CLOCK_sgo__sro_n1963));
NAND2_X1 slo__sro_c675 (.ZN (slo__sro_n514), .A1 (n_0_71), .A2 (slo__sro_n516));
NAND2_X4 slo__sro_c676 (.ZN (slo__sro_n513), .A1 (slo__sro_n515), .A2 (slo__sro_n514));
NOR2_X1 slo__sro_c698 (.ZN (slo__sro_n534), .A1 (\Res_imm[27] ), .A2 (\Res_imm[30] ));
AND2_X1 slo__sro_c699 (.ZN (n_0_1_21), .A1 (slo__sro_n534), .A2 (slo__sro_n535));
NAND2_X1 slo__mro_c626 (.ZN (slo__mro_n474), .A1 (n_0_62), .A2 (slo__xsl_n298));
NAND2_X1 slo__mro_c627 (.ZN (n_0_248), .A1 (n_0_1_2), .A2 (slo__mro_n474));
NAND2_X4 slo__sro_c708 (.ZN (slo__sro_n538), .A1 (slo__sro_n540), .A2 (slo__sro_n539));
NAND2_X2 CLOCK_slo__sro_c3800 (.ZN (CLOCK_slo__sro_n3371), .A1 (n_0_145), .A2 (drc_ipo_n26));
NAND2_X1 slo__sro_c717 (.ZN (slo__sro_n549), .A1 (n_0_97), .A2 (slo__sro_n551));
INV_X2 CLOCK_slo__c3686 (.ZN (CLOCK_slo__n3265), .A (CLOCK_slo__n2403));
NAND2_X2 slo__sro_c726 (.ZN (slo__sro_n560), .A1 (opt_ipo_n1428), .A2 (drc_ipo_n26));
NAND2_X1 slo__sro_c727 (.ZN (slo__sro_n559), .A1 (opt_ipo_n1363), .A2 (slo__sro_n561));
NAND2_X4 slo__sro_c728 (.ZN (slo__sro_n558), .A1 (slo__sro_n560), .A2 (slo__sro_n559));
NAND2_X2 slo__sro_c845 (.ZN (slo__sro_n669), .A1 (n_0_143), .A2 (drc_ipo_n26));
CLKBUF_X2 slo__c796 (.Z (slo__n619), .A (slo__n345));
NAND2_X1 slo__sro_c846 (.ZN (slo__sro_n668), .A1 (n_0_102), .A2 (slo__sro_n670));
NAND2_X4 slo__sro_c847 (.ZN (slo__sro_n667), .A1 (slo__sro_n669), .A2 (slo__sro_n668));
NAND2_X2 slo__sro_c876 (.ZN (slo__sro_n702), .A1 (n_0_177), .A2 (drc_ipo_n27));
NAND2_X1 slo__sro_c877 (.ZN (slo__sro_n701), .A1 (n_0_68), .A2 (slo__sro_n703));
NAND2_X4 slo__sro_c878 (.ZN (slo__sro_n700), .A1 (slo__sro_n702), .A2 (slo__sro_n701));
OAI22_X2 slo__sro_c1048 (.ZN (n_0_230), .A1 (hfn_ipo_n25), .A2 (n_0_1_125), .B1 (slo__n453), .B2 (n_0_1_126));
INV_X8 CLOCK_slo__c2764 (.ZN (CLOCK_slo__n2403), .A (CLOCK_slo__sro_n2424));
OR2_X1 slo__sro_c1095 (.ZN (slo__sro_n905), .A1 (n_0_1_17), .A2 (reset));
OR2_X4 slo__sro_c1096 (.ZN (slo__n798), .A1 (sgo__sro_n51), .A2 (slo__sro_n905));
OR3_X1 slo__c1065 (.ZN (slo__n881), .A1 (sgo__sro_n51), .A2 (n_0_1_17), .A3 (reset));
BUF_X4 CLOCK_slo__c2820 (.Z (CLOCK_slo__n2449), .A (slo__n798));
NAND2_X1 slo__sro_c1200 (.ZN (slo__sro_n999), .A1 (n_0_109), .A2 (slo__sro_n1001));
NAND2_X1 CLOCK_slo__sro_c2540 (.ZN (CLOCK_slo__sro_n2213), .A1 (opt_ipo_n1540), .A2 (CLOCK_slo__sro_n2215));
NOR2_X2 slo__c1173 (.ZN (slo__n980), .A1 (sgo__sro_n51), .A2 (n_0_1_17));
NOR2_X1 CLOCK_sgo__sro_c2228 (.ZN (CLOCK_sgo__sro_n1965), .A1 (\Res_imm[40] ), .A2 (\Res_imm[45] ));
NAND2_X1 slo__sro_c1291 (.ZN (slo__sro_n1080), .A1 (n_0_107), .A2 (slo__sro_n1082));
NAND2_X2 slo__sro_c1239 (.ZN (slo__sro_n1028), .A1 (n_0_137), .A2 (drc_ipo_n26));
NAND2_X1 slo__sro_c1240 (.ZN (slo__sro_n1027), .A1 (n_0_108), .A2 (slo__sro_n1029));
NAND2_X4 slo__sro_c1241 (.ZN (slo__sro_n1026), .A1 (slo__sro_n1028), .A2 (slo__sro_n1027));
NAND2_X4 slo__sro_c1292 (.ZN (slo__sro_n1079), .A1 (slo__sro_n1081), .A2 (slo__sro_n1080));
NAND2_X2 slo__sro_c1327 (.ZN (slo__sro_n1122), .A1 (n_0_135), .A2 (drc_ipo_n26));
NAND2_X1 slo__sro_c1328 (.ZN (slo__sro_n1121), .A1 (n_0_110), .A2 (slo__sro_n1123));
NAND2_X4 slo__sro_c1329 (.ZN (slo__sro_n1120), .A1 (slo__sro_n1122), .A2 (slo__sro_n1121));
NAND2_X4 CLOCK_slo__sro_c2649 (.ZN (CLOCK_slo__sro_n2298), .A1 (CLOCK_slo__sro_n2300), .A2 (CLOCK_slo__sro_n2299));
NAND2_X1 slo__sro_c1338 (.ZN (slo__sro_n1131), .A1 (slo__sro_n1133), .A2 (n_0_106));
NAND2_X1 CLOCK_slo__sro_c3056 (.ZN (CLOCK_slo__sro_n2684), .A1 (drc_ipo_n27), .A2 (n_0_168));
NAND2_X2 slo__sro_c1351 (.ZN (slo__sro_n1152), .A1 (n_0_173), .A2 (drc_ipo_n27));
NAND2_X1 slo__sro_c1352 (.ZN (slo__sro_n1151), .A1 (n_0_72), .A2 (slo__sro_n1153));
NAND2_X4 slo__sro_c1353 (.ZN (slo__sro_n1150), .A1 (slo__sro_n1152), .A2 (slo__sro_n1151));
NAND2_X2 slo__sro_c1402 (.ZN (slo__sro_n1188), .A1 (n_0_161), .A2 (drc_ipo_n27));
NAND2_X1 slo__sro_c1403 (.ZN (slo__sro_n1187), .A1 (n_0_84), .A2 (slo__sro_n1189));
NAND2_X4 slo__sro_c1404 (.ZN (slo__sro_n1186), .A1 (slo__sro_n1188), .A2 (slo__sro_n1187));
INV_X2 CLOCK_slo__mro_c3589 (.ZN (CLOCK_slo__mro_n3164), .A (slo__sro_n549));
NAND2_X4 CLOCK_slo__sro_c2541 (.ZN (CLOCK_slo__sro_n2212), .A1 (CLOCK_slo__sro_n2213), .A2 (CLOCK_slo__sro_n2214));
INV_X16 CLOCK_opt_ipo_c1940 (.ZN (CLOCK_opt_ipo_n1683), .A (A[31]));
NAND2_X4 CLOCK_slo__sro_c3480 (.ZN (CLOCK_slo__sro_n3065), .A1 (CLOCK_slo__sro_n3067), .A2 (CLOCK_slo__sro_n3066));
INV_X4 CLOCK_slo__sro_c3477 (.ZN (CLOCK_slo__sro_n3068), .A (drc_ipo_n26));
CLKBUF_X2 opt_ipo_c1602 (.Z (opt_ipo_n1344), .A (\Res_imm[50] ));
NOR3_X4 CLOCK_sgo__sro_c2218 (.ZN (n_0_1_26), .A1 (CLOCK_sgo__sro_n1959), .A2 (\Res_imm[51] ), .A3 (\Res_imm[48] ));
NAND2_X2 CLOCK_slo__sro_c3478 (.ZN (CLOCK_slo__sro_n3067), .A1 (n_0_146), .A2 (drc_ipo_n26));
INV_X1 opt_ipo_c1797 (.ZN (opt_ipo_n1540), .A (opt_ipo_n1541));
INV_X2 opt_ipo_c1798 (.ZN (opt_ipo_n1541), .A (n_0_86));
INV_X1 CLOCK_slo__mro_c2636 (.ZN (slo__sro_n1132), .A (drc_ipo_n26));
NAND2_X4 CLOCK_slo__sro_c3479 (.ZN (CLOCK_slo__sro_n3066), .A1 (n_0_99), .A2 (CLOCK_slo__sro_n3068));
INV_X2 opt_ipo_c1804 (.ZN (opt_ipo_n1547), .A (n_0_1_24));
INV_X8 opt_ipo_c1808 (.ZN (opt_ipo_n1551), .A (slo__n453));
CLKBUF_X1 opt_ipo_c1619 (.Z (opt_ipo_n1361), .A (\Res_imm[48] ));
NAND2_X1 CLOCK_slo__sro_c2648 (.ZN (CLOCK_slo__sro_n2299), .A1 (n_0_78), .A2 (CLOCK_slo__sro_n2301));
INV_X1 opt_ipo_c1621 (.ZN (opt_ipo_n1363), .A (opt_ipo_n1364));
INV_X1 opt_ipo_c1622 (.ZN (opt_ipo_n1364), .A (n_0_113));
CLKBUF_X2 opt_ipo_c1623 (.Z (opt_ipo_n1365), .A (\Res_imm[62] ));
NAND2_X2 CLOCK_slo__mro_c2661 (.ZN (slo__sro_n1000), .A1 (n_0_136), .A2 (drc_ipo_n26));
INV_X8 opt_ipo_c1812 (.ZN (opt_ipo_n1555), .A (CLOCK_slo__n2403));
OR2_X4 CLOCK_slo__sro_c3036 (.ZN (CLOCK_slo__sro_n2662), .A1 (sgo__sro_n51), .A2 (CLOCK_slo__sro_n2663));
NAND2_X4 CLOCK_slo__sro_c2788 (.ZN (CLOCK_slo__sro_n2425), .A1 (opt_ipo_n1652), .A2 (hfn_ipo_n23));
INV_X8 CLOCK_slo__sro_c2789 (.ZN (CLOCK_slo__sro_n2424), .A (CLOCK_slo__sro_n2425));
INV_X1 CLOCK_slo__sro_c3055 (.ZN (CLOCK_slo__sro_n2685), .A (drc_ipo_n27));
CLKBUF_X3 opt_ipo_c1637 (.Z (Res[63]), .A (opt_ipo_n1380));
BUF_X4 CLOCK_slo__c2998 (.Z (CLOCK_slo__n2626), .A (slo__n798));
INV_X1 opt_ipo_c1826 (.ZN (opt_ipo_n1569), .A (n_0_1_9));
INV_X16 CLOCK_sgo__c2073 (.ZN (slo__n453), .A (CLOCK_slo__sro_n2424));
NAND2_X4 CLOCK_slo__sro_c3058 (.ZN (CLOCK_slo__sro_n2682), .A1 (CLOCK_slo__sro_n2684), .A2 (CLOCK_slo__sro_n2683));
INV_X1 CLOCK_slo__sro_c3169 (.ZN (CLOCK_slo__sro_n2796), .A (drc_ipo_n27));
NAND2_X2 CLOCK_slo__sro_c3170 (.ZN (CLOCK_slo__sro_n2795), .A1 (n_0_176), .A2 (drc_ipo_n27));
NAND2_X1 CLOCK_slo__sro_c3171 (.ZN (CLOCK_slo__sro_n2794), .A1 (n_0_69), .A2 (CLOCK_slo__sro_n2796));
NAND2_X4 CLOCK_slo__sro_c3172 (.ZN (CLOCK_slo__sro_n2793), .A1 (CLOCK_slo__sro_n2795), .A2 (CLOCK_slo__sro_n2794));
NAND2_X2 CLOCK_slo__sro_c3218 (.ZN (CLOCK_slo__sro_n2843), .A1 (n_0_158), .A2 (drc_ipo_n27));
NAND2_X4 CLOCK_slo__sro_c3220 (.ZN (CLOCK_slo__sro_n2841), .A1 (CLOCK_slo__sro_n2843), .A2 (CLOCK_slo__sro_n2842));
INV_X8 CLOCK_slo__mro_c3591 (.ZN (CLOCK_slo__mro_n3162), .A (CLOCK_slo__mro_n3163));
NAND2_X4 CLOCK_slo__sro_c3801 (.ZN (CLOCK_slo__sro_n3370), .A1 (n_0_100), .A2 (CLOCK_slo__sro_n3372));
NAND2_X4 CLOCK_slo__sro_c3802 (.ZN (CLOCK_slo__sro_n3369), .A1 (CLOCK_slo__sro_n3371), .A2 (CLOCK_slo__sro_n3370));
INV_X1 opt_ipo_c1855 (.ZN (opt_ipo_n1598), .A (n_0_126));
CLKBUF_X1 CLOCK_slh__c3970 (.Z (CLOCK_slh__n3500), .A (CLOCK_slh__n3499));
CLKBUF_X1 CLOCK_slh__c3971 (.Z (CLOCK_slh__n3501), .A (CLOCK_slh__n3500));
CLKBUF_X1 CLOCK_slh__c3972 (.Z (CLOCK_slh__n3509), .A (CLOCK_slh__n3501));
INV_X8 CLOCK_slo__sro_c3799 (.ZN (CLOCK_slo__sro_n3372), .A (drc_ipo_n26));
CLKBUF_X1 CLOCK_slh__c3980 (.Z (CLOCK_slh__n3510), .A (CLOCK_slh__n3509));
CLKBUF_X1 CLOCK_slh__c3981 (.Z (CLOCK_slh__n3511), .A (CLOCK_slh__n3510));
INV_X2 opt_ipo_c1685 (.ZN (opt_ipo_n1428), .A (n_0_132));
CLKBUF_X1 CLOCK_slh__c3982 (.Z (CLOCK_slh__n3519), .A (CLOCK_slh__n3511));
CLKBUF_X1 CLOCK_slh__c3990 (.Z (CLOCK_slh__n3520), .A (CLOCK_slh__n3519));
CLKBUF_X1 CLOCK_slh__c3991 (.Z (CLOCK_slh__n3521), .A (CLOCK_slh__n3520));
CLKBUF_X1 CLOCK_slh__c3992 (.Z (CLOCK_slh__n3529), .A (CLOCK_slh__n3521));
CLKBUF_X1 CLOCK_slh__c4000 (.Z (CLOCK_slh__n3530), .A (CLOCK_slh__n3529));
CLKBUF_X1 CLOCK_slh__c4001 (.Z (CLOCK_slh__n3531), .A (CLOCK_slh__n3530));
CLKBUF_X1 CLOCK_slh__c4002 (.Z (CLOCK_slh__n3535), .A (CLOCK_slh__n3531));
CLKBUF_X1 CLOCK_slh__c4006 (.Z (CLOCK_slh__n3536), .A (CLOCK_slh__n3535));
CLKBUF_X1 CLOCK_slh__c4007 (.Z (CLOCK_slh__n3537), .A (CLOCK_slh__n3536));
CLKBUF_X1 CLOCK_slh__c4008 (.Z (CLOCK_slh__n3541), .A (CLOCK_slh__n3537));
CLKBUF_X1 CLOCK_slh__c4012 (.Z (CLOCK_slh__n3542), .A (CLOCK_slh__n3541));
CLKBUF_X1 CLOCK_slh__c4013 (.Z (CLOCK_slh__n3543), .A (CLOCK_slh__n3542));
CLKBUF_X1 CLOCK_slh__c4014 (.Z (CLOCK_slh__n3547), .A (CLOCK_slh__n3543));
CLKBUF_X1 CLOCK_slh__c4018 (.Z (CLOCK_slh__n3548), .A (CLOCK_slh__n3547));
CLKBUF_X1 CLOCK_slh__c4019 (.Z (CLOCK_slh__n3549), .A (CLOCK_slh__n3548));
CLKBUF_X1 CLOCK_slh__c4020 (.Z (CLOCK_slh__n3553), .A (CLOCK_slh__n3549));
CLKBUF_X1 CLOCK_slh__c4024 (.Z (CLOCK_slh__n3554), .A (CLOCK_slh__n3553));
CLKBUF_X1 CLOCK_slh__c4025 (.Z (CLOCK_slh__n3555), .A (CLOCK_slh__n3554));
CLKBUF_X1 CLOCK_slh__c4026 (.Z (sph__n4211), .A (CLOCK_slh__n3555));
CLKBUF_X1 sph__c4660 (.Z (sph__n4212), .A (sph__n4211));
CLKBUF_X1 sph__c4661 (.Z (CLOCK_slh_n3498), .A (sph__n4212));

endmodule //multiplierTree


