/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 16 23:47:43 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 747355786 */

module datapath__0_0(A_imm, A_imm_2s_complement);
   input [31:0]A_imm;
   output [31:0]A_imm_2s_complement;

   AOI21_X1 i_0 (.A(n_43), .B1(A_imm[2]), .B2(n_38), .ZN(A_imm_2s_complement[2]));
   AOI21_X1 i_1 (.A(n_5), .B1(A_imm[4]), .B2(n_45), .ZN(A_imm_2s_complement[4]));
   AOI21_X1 i_2 (.A(n_3), .B1(A_imm[5]), .B2(n_4), .ZN(A_imm_2s_complement[5]));
   AOI21_X1 i_3 (.A(n_1), .B1(A_imm[6]), .B2(n_2), .ZN(A_imm_2s_complement[6]));
   AOI21_X1 i_4 (.A(n_40), .B1(A_imm[7]), .B2(n_0), .ZN(A_imm_2s_complement[7]));
   INV_X1 i_5 (.A(n_1), .ZN(n_0));
   NOR2_X1 i_6 (.A1(n_45), .A2(n_50), .ZN(n_1));
   INV_X1 i_7 (.A(n_3), .ZN(n_2));
   NOR2_X1 i_8 (.A1(A_imm[5]), .A2(n_4), .ZN(n_3));
   INV_X1 i_9 (.A(n_5), .ZN(n_4));
   NOR2_X1 i_10 (.A1(A_imm[4]), .A2(n_45), .ZN(n_5));
   AOI21_X1 i_11 (.A(n_9), .B1(A_imm[9]), .B2(n_10), .ZN(A_imm_2s_complement[9]));
   AOI21_X1 i_12 (.A(n_7), .B1(A_imm[10]), .B2(n_8), .ZN(A_imm_2s_complement[10]));
   AOI21_X1 i_13 (.A(n_37), .B1(A_imm[11]), .B2(n_6), .ZN(
      A_imm_2s_complement[11]));
   INV_X1 i_14 (.A(n_7), .ZN(n_6));
   NOR2_X1 i_15 (.A1(n_47), .A2(n_56), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   NOR2_X1 i_17 (.A1(A_imm[9]), .A2(n_10), .ZN(n_9));
   INV_X1 i_18 (.A(n_46), .ZN(n_10));
   AOI21_X1 i_19 (.A(n_17), .B1(A_imm[12]), .B2(n_36), .ZN(
      A_imm_2s_complement[12]));
   AOI21_X1 i_20 (.A(n_15), .B1(A_imm[13]), .B2(n_16), .ZN(
      A_imm_2s_complement[13]));
   AOI21_X1 i_21 (.A(n_13), .B1(A_imm[14]), .B2(n_14), .ZN(
      A_imm_2s_complement[14]));
   AOI21_X1 i_22 (.A(n_34), .B1(A_imm[15]), .B2(n_12), .ZN(
      A_imm_2s_complement[15]));
   INV_X1 i_23 (.A(n_13), .ZN(n_12));
   NOR2_X1 i_24 (.A1(n_36), .A2(n_54), .ZN(n_13));
   INV_X1 i_25 (.A(n_15), .ZN(n_14));
   NOR2_X1 i_26 (.A1(A_imm[13]), .A2(n_16), .ZN(n_15));
   INV_X1 i_27 (.A(n_17), .ZN(n_16));
   NOR2_X1 i_28 (.A1(A_imm[12]), .A2(n_36), .ZN(n_17));
   AOI21_X1 i_29 (.A(n_23), .B1(A_imm[16]), .B2(n_33), .ZN(
      A_imm_2s_complement[16]));
   AOI21_X1 i_30 (.A(n_21), .B1(A_imm[17]), .B2(n_22), .ZN(
      A_imm_2s_complement[17]));
   AOI21_X1 i_31 (.A(n_19), .B1(A_imm[18]), .B2(n_20), .ZN(
      A_imm_2s_complement[18]));
   AOI21_X1 i_32 (.A(n_31), .B1(A_imm[19]), .B2(n_18), .ZN(
      A_imm_2s_complement[19]));
   INV_X1 i_33 (.A(n_19), .ZN(n_18));
   NOR2_X1 i_34 (.A1(n_33), .A2(n_52), .ZN(n_19));
   INV_X1 i_35 (.A(n_21), .ZN(n_20));
   NOR2_X1 i_36 (.A1(A_imm[17]), .A2(n_22), .ZN(n_21));
   INV_X1 i_37 (.A(n_23), .ZN(n_22));
   NOR2_X1 i_38 (.A1(A_imm[16]), .A2(n_33), .ZN(n_23));
   AOI21_X1 i_39 (.A(n_25), .B1(A_imm[20]), .B2(n_30), .ZN(
      A_imm_2s_complement[20]));
   NOR2_X1 i_40 (.A1(A_imm[20]), .A2(n_30), .ZN(n_25));
   AOI21_X1 i_41 (.A(n_24), .B1(n_26), .B2(A_imm[21]), .ZN(
      A_imm_2s_complement[21]));
   INV_X1 i_42 (.A(n_27), .ZN(n_24));
   INV_X1 i_43 (.A(n_25), .ZN(n_26));
   AOI21_X1 i_44 (.A(n_28), .B1(n_27), .B2(A_imm[22]), .ZN(
      A_imm_2s_complement[22]));
   NAND3_X1 i_45 (.A1(n_31), .A2(n_32), .A3(n_11), .ZN(n_27));
   INV_X1 i_46 (.A(n_48), .ZN(n_28));
   INV_X1 i_47 (.A(n_29), .ZN(A_imm_2s_complement[23]));
   XNOR2_X1 i_48 (.A(n_48), .B(A_imm[23]), .ZN(n_29));
   OR2_X1 i_49 (.A1(n_48), .A2(A_imm[23]), .ZN(A_imm_2s_complement[27]));
   NAND4_X1 i_50 (.A1(n_31), .A2(n_35), .A3(n_32), .A4(n_11), .ZN(n_48));
   INV_X1 i_51 (.A(n_30), .ZN(n_31));
   NAND2_X1 i_52 (.A1(n_34), .A2(n_51), .ZN(n_30));
   INV_X1 i_53 (.A(n_33), .ZN(n_34));
   NAND2_X1 i_54 (.A1(n_37), .A2(n_53), .ZN(n_33));
   INV_X1 i_55 (.A(n_36), .ZN(n_37));
   NAND2_X1 i_56 (.A1(n_40), .A2(n_55), .ZN(n_36));
   INV_X1 i_57 (.A(n_47), .ZN(n_40));
   INV_X1 i_58 (.A(A_imm[20]), .ZN(n_11));
   INV_X1 i_59 (.A(A_imm[21]), .ZN(n_32));
   INV_X1 i_60 (.A(A_imm[22]), .ZN(n_35));
   AOI21_X1 i_61 (.A(n_39), .B1(A_imm[1]), .B2(A_imm[0]), .ZN(
      A_imm_2s_complement[1]));
   INV_X1 i_62 (.A(n_39), .ZN(n_38));
   NOR2_X1 i_63 (.A1(A_imm[1]), .A2(A_imm[0]), .ZN(n_39));
   INV_X1 i_64 (.A(A_imm[2]), .ZN(n_41));
   NAND2_X1 i_65 (.A1(n_41), .A2(n_39), .ZN(n_42));
   INV_X1 i_66 (.A(n_42), .ZN(n_43));
   NOR2_X1 i_67 (.A1(n_42), .A2(A_imm[3]), .ZN(n_44));
   INV_X1 i_68 (.A(n_44), .ZN(n_45));
   AOI21_X1 i_69 (.A(n_44), .B1(A_imm[3]), .B2(n_42), .ZN(A_imm_2s_complement[3]));
   AOI21_X1 i_70 (.A(n_46), .B1(A_imm[8]), .B2(n_47), .ZN(A_imm_2s_complement[8]));
   NOR2_X1 i_71 (.A1(A_imm[8]), .A2(n_47), .ZN(n_46));
   NAND2_X1 i_72 (.A1(n_44), .A2(n_49), .ZN(n_47));
   NOR2_X1 i_73 (.A1(A_imm[7]), .A2(n_50), .ZN(n_49));
   OR3_X1 i_74 (.A1(A_imm[5]), .A2(A_imm[4]), .A3(A_imm[6]), .ZN(n_50));
   NOR2_X1 i_75 (.A1(A_imm[19]), .A2(n_52), .ZN(n_51));
   OR3_X1 i_76 (.A1(A_imm[17]), .A2(A_imm[16]), .A3(A_imm[18]), .ZN(n_52));
   NOR2_X1 i_77 (.A1(A_imm[15]), .A2(n_54), .ZN(n_53));
   OR3_X1 i_78 (.A1(A_imm[13]), .A2(A_imm[12]), .A3(A_imm[14]), .ZN(n_54));
   NOR2_X1 i_79 (.A1(A_imm[11]), .A2(n_56), .ZN(n_55));
   OR3_X1 i_80 (.A1(A_imm[9]), .A2(A_imm[8]), .A3(A_imm[10]), .ZN(n_56));
endmodule

module datapath__0_67(p_0, p_1, p_2, p_3, p_4, p_5, p_6, p_7, p_8, p_9, p_10, 
      p_11, p_12, p_13, p_14, p_15, \aggregated_res[14] );
   input [63:0]p_0;
   input [63:0]p_1;
   input [63:0]p_2;
   input [63:0]p_3;
   input [63:0]p_4;
   input [63:0]p_5;
   input [63:0]p_6;
   input [63:0]p_7;
   input [63:0]p_8;
   input [63:0]p_9;
   input [63:0]p_10;
   input [63:0]p_11;
   input [63:0]p_12;
   input [63:0]p_13;
   input [63:0]p_14;
   input [63:0]p_15;
   output [63:0]\aggregated_res[14] ;

   FA_X1 i_58 (.A(p_6[18]), .B(p_7[18]), .CI(p_8[18]), .CO(n_117), .S(n_116));
   XOR2_X1 i_0 (.A(p_3[40]), .B(p_4[33]), .Z(n_179));
   OAI21_X1 i_1 (.A(n_661), .B1(n_665), .B2(n_662), .ZN(n_198));
   XOR2_X1 i_290 (.A(p_2[38]), .B(p_3[31]), .Z(n_201));
   OAI222_X1 i_2 (.A1(p_2[38]), .A2(n_209), .B1(p_2[38]), .B2(n_786), .C1(n_786), 
      .C2(n_209), .ZN(n_203));
   XOR2_X1 i_3 (.A(n_567), .B(n_563), .Z(\aggregated_res[14] [24]));
   AOI21_X1 i_4 (.A(n_489), .B1(n_269), .B2(n_405), .ZN(n_563));
   XOR2_X1 i_5 (.A(n_570), .B(n_564), .Z(\aggregated_res[14] [25]));
   AOI21_X1 i_6 (.A(n_489), .B1(n_485), .B2(n_566), .ZN(n_564));
   INV_X1 i_7 (.A(n_567), .ZN(n_566));
   AOI21_X1 i_8 (.A(n_277), .B1(n_491), .B2(n_281), .ZN(n_567));
   AOI21_X1 i_9 (.A(n_487), .B1(n_407), .B2(n_409), .ZN(n_570));
   XOR2_X1 i_10 (.A(n_552), .B(n_573), .Z(\aggregated_res[14] [27]));
   XOR2_X1 i_11 (.A(n_545), .B(n_571), .Z(\aggregated_res[14] [28]));
   NOR2_X1 i_12 (.A1(n_574), .A2(n_568), .ZN(n_571));
   NOR2_X1 i_13 (.A1(n_565), .A2(n_557), .ZN(n_573));
   XOR2_X1 i_14 (.A(n_581), .B(n_580), .Z(\aggregated_res[14] [32]));
   OAI21_X1 i_15 (.A(n_626), .B1(n_627), .B2(n_624), .ZN(n_580));
   OAI21_X1 i_16 (.A(n_652), .B1(n_621), .B2(n_633), .ZN(n_581));
   XOR2_X1 i_17 (.A(n_593), .B(n_582), .Z(\aggregated_res[14] [33]));
   OAI21_X1 i_18 (.A(n_652), .B1(n_739), .B2(n_630), .ZN(n_582));
   AOI21_X1 i_19 (.A(n_660), .B1(n_634), .B2(n_631), .ZN(n_593));
   XOR2_X1 i_20 (.A(n_685), .B(n_596), .Z(\aggregated_res[14] [35]));
   XOR2_X1 i_21 (.A(n_684), .B(n_594), .Z(\aggregated_res[14] [36]));
   NOR2_X1 i_22 (.A1(n_708), .A2(n_690), .ZN(n_594));
   AOI21_X1 i_23 (.A(n_689), .B1(n_643), .B2(n_675), .ZN(n_596));
   XOR2_X1 i_24 (.A(n_732), .B(n_604), .Z(\aggregated_res[14] [39]));
   XOR2_X1 i_25 (.A(n_731), .B(n_602), .Z(\aggregated_res[14] [40]));
   NOR2_X1 i_26 (.A1(n_754), .A2(n_737), .ZN(n_602));
   AOI21_X1 i_27 (.A(n_736), .B1(n_703), .B2(n_722), .ZN(n_604));
   XOR2_X1 i_28 (.A(n_781), .B(n_775), .Z(\aggregated_res[14] [43]));
   XNOR2_X1 i_29 (.A(n_611), .B(n_610), .ZN(\aggregated_res[14] [44]));
   OAI22_X1 i_30 (.A1(n_749), .A2(n_765), .B1(n_777), .B2(n_781), .ZN(n_610));
   NOR2_X1 i_31 (.A1(n_774), .A2(n_779), .ZN(n_611));
   AND2_X1 i_455 (.A1(p_0[3]), .A2(p_15[3]), .ZN(n_205));
   AND2_X1 i_456 (.A1(p_0[2]), .A2(p_15[2]), .ZN(n_207));
   INV_X1 i_32 (.A(p_4[31]), .ZN(n_209));
   INV_X1 i_33 (.A(p_3[31]), .ZN(n_786));
   OAI21_X1 i_34 (.A(n_626), .B1(n_621), .B2(n_633), .ZN(n_739));
   XNOR2_X1 i_35 (.A(p_1[27]), .B(p_0[34]), .ZN(n_211));
   FA_X1 i_36 (.A(p_3[19]), .B(p_4[19]), .CI(p_5[19]), .CO(n_131), .S(n_130));
   FA_X1 i_37 (.A(p_0[19]), .B(p_1[19]), .CI(p_2[19]), .CO(n_129), .S(n_128));
   FA_X1 i_38 (.A(p_15[19]), .B(n_117), .CI(n_115), .CO(n_135), .S(n_134));
   FA_X1 i_39 (.A(n_130), .B(n_128), .CI(n_134), .CO(n_139), .S(n_138));
   FA_X1 i_40 (.A(n_102), .B(n_100), .CI(n_98), .CO(n_107), .S(n_106));
   FA_X1 i_41 (.A(n_99), .B(n_105), .CI(n_116), .CO(n_121), .S(n_120));
   FA_X1 i_42 (.A(n_91), .B(n_104), .CI(n_93), .CO(n_109), .S(n_108));
   FA_X1 i_43 (.A(n_107), .B(n_120), .CI(n_109), .CO(n_125), .S(n_124));
   FA_X1 i_44 (.A(n_113), .B(n_119), .CI(n_132), .CO(n_137), .S(n_136));
   FA_X1 i_45 (.A(n_114), .B(n_112), .CI(n_118), .CO(n_123), .S(n_122));
   FA_X1 i_46 (.A(n_121), .B(n_136), .CI(n_123), .CO(n_141), .S(n_140));
   FA_X1 i_47 (.A(n_138), .B(n_125), .CI(n_140), .CO(n_143), .S(n_142));
   FA_X1 i_48 (.A(p_0[20]), .B(p_1[20]), .CI(p_2[20]), .CO(n_145), .S(n_144));
   FA_X1 i_49 (.A(n_131), .B(n_129), .CI(n_135), .CO(n_153), .S(n_152));
   FA_X1 i_50 (.A(n_144), .B(n_152), .CI(n_137), .CO(n_157), .S(n_156));
   FA_X1 i_51 (.A(n_150), .B(n_148), .CI(n_146), .CO(n_155), .S(n_154));
   FA_X1 i_52 (.A(n_139), .B(n_154), .CI(n_141), .CO(n_159), .S(n_158));
   HA_X1 i_53 (.A(n_156), .B(n_158), .CO(n_161), .S(n_160));
   FA_X1 i_54 (.A(p_0[21]), .B(p_1[21]), .CI(p_2[21]), .CO(n_163), .S(n_162));
   FA_X1 i_55 (.A(n_147), .B(n_145), .CI(n_151), .CO(n_171), .S(n_170));
   FA_X1 i_56 (.A(n_162), .B(n_153), .CI(n_170), .CO(n_175), .S(n_174));
   FA_X1 i_57 (.A(n_168), .B(n_166), .CI(n_164), .CO(n_173), .S(n_172));
   FA_X1 i_59 (.A(n_155), .B(n_157), .CI(n_172), .CO(n_177), .S(n_176));
   FA_X1 i_60 (.A(n_174), .B(n_159), .CI(n_176), .CO(n_213), .S(n_178));
   FA_X1 i_61 (.A(p_3[18]), .B(p_4[18]), .CI(p_5[18]), .CO(n_115), .S(n_114));
   FA_X1 i_62 (.A(p_0[18]), .B(p_1[18]), .CI(p_2[18]), .CO(n_113), .S(n_112));
   FA_X1 i_63 (.A(p_15[18]), .B(n_103), .CI(n_101), .CO(n_119), .S(n_118));
   HA_X1 i_64 (.A(n_122), .B(n_124), .CO(n_127), .S(n_126));
   FA_X1 i_65 (.A(p_6[17]), .B(p_7[17]), .CI(p_15[17]), .CO(n_103), .S(n_102));
   FA_X1 i_66 (.A(p_3[17]), .B(p_4[17]), .CI(p_5[17]), .CO(n_101), .S(n_100));
   FA_X1 i_67 (.A(p_0[17]), .B(p_1[17]), .CI(p_2[17]), .CO(n_99), .S(n_98));
   FA_X1 i_68 (.A(n_75), .B(n_73), .CI(n_77), .CO(n_91), .S(n_90));
   FA_X1 i_69 (.A(n_61), .B(n_65), .CI(n_76), .CO(n_79), .S(n_78));
   FA_X1 i_70 (.A(n_74), .B(n_72), .CI(n_67), .CO(n_81), .S(n_80));
   FA_X1 i_71 (.A(n_90), .B(n_79), .CI(n_81), .CO(n_95), .S(n_94));
   FA_X1 i_72 (.A(n_89), .B(n_87), .CI(n_85), .CO(n_105), .S(n_104));
   FA_X1 i_73 (.A(n_88), .B(n_86), .CI(n_84), .CO(n_93), .S(n_92));
   FA_X1 i_74 (.A(n_106), .B(n_95), .CI(n_108), .CO(n_111), .S(n_110));
   FA_X1 i_75 (.A(p_0[14]), .B(p_1[14]), .CI(p_2[14]), .CO(n_61), .S(n_60));
   FA_X1 i_76 (.A(p_3[13]), .B(p_4[13]), .CI(p_5[13]), .CO(n_53), .S(n_52));
   FA_X1 i_77 (.A(p_6[14]), .B(p_15[14]), .CI(n_53), .CO(n_65), .S(n_64));
   FA_X1 i_78 (.A(p_3[14]), .B(p_4[14]), .CI(p_5[14]), .CO(n_63), .S(n_62));
   FA_X1 i_79 (.A(p_6[15]), .B(p_15[15]), .CI(n_63), .CO(n_77), .S(n_76));
   FA_X1 i_80 (.A(p_15[12]), .B(n_35), .CI(n_33), .CO(n_45), .S(n_44));
   FA_X1 i_81 (.A(p_0[13]), .B(p_1[13]), .CI(p_2[13]), .CO(n_51), .S(n_50));
   FA_X1 i_82 (.A(n_45), .B(n_52), .CI(n_50), .CO(n_57), .S(n_56));
   FA_X1 i_83 (.A(n_62), .B(n_60), .CI(n_57), .CO(n_69), .S(n_68));
   FA_X1 i_84 (.A(p_3[15]), .B(p_4[15]), .CI(p_5[15]), .CO(n_75), .S(n_74));
   FA_X1 i_85 (.A(p_0[15]), .B(p_1[15]), .CI(p_2[15]), .CO(n_73), .S(n_72));
   FA_X1 i_86 (.A(p_15[13]), .B(n_43), .CI(n_41), .CO(n_55), .S(n_54));
   FA_X1 i_87 (.A(n_51), .B(n_55), .CI(n_64), .CO(n_67), .S(n_66));
   FA_X1 i_88 (.A(n_78), .B(n_69), .CI(n_80), .CO(n_83), .S(n_82));
   FA_X1 i_89 (.A(p_6[16]), .B(p_7[16]), .CI(p_15[16]), .CO(n_89), .S(n_88));
   FA_X1 i_90 (.A(p_3[16]), .B(p_4[16]), .CI(p_5[16]), .CO(n_87), .S(n_86));
   FA_X1 i_91 (.A(p_0[16]), .B(p_1[16]), .CI(p_2[16]), .CO(n_85), .S(n_84));
   HA_X1 i_92 (.A(n_92), .B(n_94), .CO(n_97), .S(n_96));
   HA_X1 i_93 (.A(n_66), .B(n_68), .CO(n_71), .S(n_70));
   FA_X1 i_94 (.A(p_3[12]), .B(p_4[12]), .CI(p_5[12]), .CO(n_43), .S(n_42));
   FA_X1 i_95 (.A(p_0[12]), .B(p_1[12]), .CI(p_2[12]), .CO(n_41), .S(n_40));
   FA_X1 i_96 (.A(p_3[11]), .B(p_4[11]), .CI(p_15[11]), .CO(n_35), .S(n_34));
   FA_X1 i_97 (.A(p_0[11]), .B(p_1[11]), .CI(p_2[11]), .CO(n_33), .S(n_32));
   FA_X1 i_98 (.A(n_42), .B(n_40), .CI(n_44), .CO(n_47), .S(n_46));
   FA_X1 i_99 (.A(n_54), .B(n_47), .CI(n_56), .CO(n_59), .S(n_58));
   FA_X1 i_100 (.A(n_27), .B(n_25), .CI(n_34), .CO(n_37), .S(n_36));
   FA_X1 i_101 (.A(n_32), .B(n_29), .CI(n_36), .CO(n_39), .S(n_38));
   HA_X1 i_102 (.A(n_37), .B(n_39), .CO(n_49), .S(n_48));
   FA_X1 i_103 (.A(p_0[10]), .B(p_1[10]), .CI(p_2[10]), .CO(n_25), .S(n_24));
   FA_X1 i_104 (.A(n_15), .B(n_20), .CI(n_18), .CO(n_23), .S(n_22));
   HA_X1 i_105 (.A(n_24), .B(n_23), .CO(n_31), .S(n_30));
   FA_X1 i_106 (.A(n_19), .B(n_21), .CI(n_26), .CO(n_29), .S(n_28));
   FA_X1 i_107 (.A(p_0[9]), .B(p_1[9]), .CI(p_2[9]), .CO(n_19), .S(n_18));
   FA_X1 i_108 (.A(p_3[9]), .B(p_15[9]), .CI(n_13), .CO(n_21), .S(n_20));
   FA_X1 i_109 (.A(p_3[10]), .B(p_4[10]), .CI(p_15[10]), .CO(n_27), .S(n_26));
   FA_X1 i_110 (.A(p_0[8]), .B(p_1[8]), .CI(p_2[8]), .CO(n_13), .S(n_12));
   FA_X1 i_111 (.A(p_15[7]), .B(n_5), .CI(n_7), .CO(n_11), .S(n_10));
   FA_X1 i_112 (.A(p_3[8]), .B(p_15[8]), .CI(n_9), .CO(n_15), .S(n_14));
   HA_X1 i_113 (.A(n_11), .B(n_14), .CO(n_17), .S(n_16));
   FA_X1 i_114 (.A(p_0[7]), .B(p_1[7]), .CI(p_2[7]), .CO(n_9), .S(n_8));
   FA_X1 i_115 (.A(p_0[6]), .B(p_1[6]), .CI(p_2[6]), .CO(n_5), .S(n_4));
   HA_X1 i_116 (.A(p_15[6]), .B(n_3), .CO(n_7), .S(n_6));
   FA_X1 i_117 (.A(p_0[5]), .B(p_1[5]), .CI(p_15[5]), .CO(n_3), .S(n_2));
   HA_X1 i_118 (.A(p_0[4]), .B(p_1[4]), .CO(n_1), .S(n_0));
   FA_X1 i_119 (.A(p_3[22]), .B(p_4[22]), .CI(p_5[22]), .CO(n_183), .S(n_182));
   FA_X1 i_120 (.A(p_0[22]), .B(p_1[22]), .CI(p_2[22]), .CO(n_181), .S(n_180));
   FA_X1 i_121 (.A(p_3[20]), .B(p_4[20]), .CI(p_5[20]), .CO(n_147), .S(n_146));
   FA_X1 i_122 (.A(p_6[19]), .B(p_7[19]), .CI(p_8[19]), .CO(n_133), .S(n_132));
   FA_X1 i_123 (.A(p_9[20]), .B(p_15[20]), .CI(n_133), .CO(n_151), .S(n_150));
   FA_X1 i_124 (.A(n_182), .B(n_180), .CI(n_171), .CO(n_193), .S(n_192));
   FA_X1 i_125 (.A(p_6[20]), .B(p_7[20]), .CI(p_8[20]), .CO(n_149), .S(n_148));
   FA_X1 i_126 (.A(p_9[21]), .B(p_15[21]), .CI(n_149), .CO(n_169), .S(n_168));
   FA_X1 i_127 (.A(p_9[22]), .B(p_10[22]), .CI(p_15[22]), .CO(n_187), .S(n_186));
   FA_X1 i_128 (.A(p_6[22]), .B(p_7[22]), .CI(p_8[22]), .CO(n_185), .S(n_184));
   FA_X1 i_129 (.A(n_169), .B(n_186), .CI(n_184), .CO(n_191), .S(n_190));
   FA_X1 i_130 (.A(p_6[21]), .B(p_7[21]), .CI(p_8[21]), .CO(n_167), .S(n_166));
   FA_X1 i_131 (.A(p_3[21]), .B(p_4[21]), .CI(p_5[21]), .CO(n_165), .S(n_164));
   FA_X1 i_132 (.A(n_167), .B(n_165), .CI(n_163), .CO(n_189), .S(n_188));
   FA_X1 i_133 (.A(n_188), .B(n_173), .CI(n_175), .CO(n_195), .S(n_194));
   FA_X1 i_134 (.A(n_192), .B(n_190), .CI(n_194), .CO(n_197), .S(n_196));
   HA_X1 i_135 (.A(n_177), .B(n_196), .CO(n_199), .S(n_215));
   FA_X1 i_136 (.A(n_187), .B(n_185), .CI(n_183), .CO(n_217), .S(n_208));
   FA_X1 i_137 (.A(n_208), .B(n_191), .CI(n_193), .CO(n_219), .S(n_214));
   FA_X1 i_138 (.A(p_9[23]), .B(p_10[23]), .CI(p_15[23]), .CO(n_240), .S(n_206));
   FA_X1 i_139 (.A(n_181), .B(n_189), .CI(n_206), .CO(n_241), .S(n_210));
   FA_X1 i_140 (.A(p_6[23]), .B(p_7[23]), .CI(p_8[23]), .CO(n_260), .S(n_204));
   FA_X1 i_141 (.A(p_3[23]), .B(p_4[23]), .CI(p_5[23]), .CO(n_261), .S(n_202));
   FA_X1 i_142 (.A(p_0[23]), .B(p_1[23]), .CI(p_2[23]), .CO(n_263), .S(n_200));
   FA_X1 i_143 (.A(n_204), .B(n_202), .CI(n_200), .CO(n_265), .S(n_212));
   FA_X1 i_144 (.A(n_210), .B(n_212), .CI(n_195), .CO(n_267), .S(n_216));
   FA_X1 i_145 (.A(n_214), .B(n_197), .CI(n_216), .CO(n_269), .S(n_218));
   XNOR2_X1 i_146 (.A(n_273), .B(n_271), .ZN(\aggregated_res[14] [23]));
   NOR2_X1 i_147 (.A1(n_277), .A2(n_275), .ZN(n_271));
   AOI21_X1 i_148 (.A(n_279), .B1(n_213), .B2(n_215), .ZN(n_273));
   AND2_X1 i_149 (.A1(n_199), .A2(n_218), .ZN(n_275));
   NOR2_X1 i_150 (.A1(n_199), .A2(n_218), .ZN(n_277));
   INV_X1 i_151 (.A(n_281), .ZN(n_279));
   OAI21_X1 i_152 (.A(n_282), .B1(n_213), .B2(n_215), .ZN(n_281));
   NAND3_X1 i_153 (.A1(n_369), .A2(n_367), .A3(n_283), .ZN(n_282));
   OAI211_X1 i_154 (.A(n_323), .B(n_390), .C1(n_126), .C2(n_111), .ZN(n_283));
   OAI222_X1 i_155 (.A1(n_331), .A2(n_327), .B1(n_333), .B2(n_325), .C1(n_331), 
      .C2(n_329), .ZN(n_323));
   AOI22_X1 i_156 (.A1(n_110), .A2(n_97), .B1(n_83), .B2(n_96), .ZN(n_325));
   AOI22_X1 i_157 (.A1(n_70), .A2(n_59), .B1(n_82), .B2(n_71), .ZN(n_327));
   OAI22_X1 i_158 (.A1(n_339), .A2(n_335), .B1(n_70), .B2(n_59), .ZN(n_329));
   OAI222_X1 i_159 (.A1(n_83), .A2(n_96), .B1(n_110), .B2(n_97), .C1(n_82), 
      .C2(n_71), .ZN(n_331));
   NOR2_X1 i_160 (.A1(n_110), .A2(n_97), .ZN(n_333));
   NOR2_X1 i_161 (.A1(n_362), .A2(n_337), .ZN(n_335));
   AOI22_X1 i_162 (.A1(n_58), .A2(n_49), .B1(n_46), .B2(n_48), .ZN(n_337));
   AOI211_X1 i_163 (.A(n_365), .B(n_361), .C1(n_359), .C2(n_340), .ZN(n_339));
   OAI21_X1 i_164 (.A(n_341), .B1(n_30), .B2(n_28), .ZN(n_340));
   OAI222_X1 i_165 (.A1(n_351), .A2(n_345), .B1(n_353), .B2(n_343), .C1(n_355), 
      .C2(n_347), .ZN(n_341));
   AOI22_X1 i_166 (.A1(n_12), .A2(n_16), .B1(n_22), .B2(n_17), .ZN(n_343));
   AOI22_X1 i_167 (.A1(n_4), .A2(n_6), .B1(n_10), .B2(n_8), .ZN(n_345));
   OAI221_X1 i_168 (.A(n_349), .B1(n_4), .B2(n_6), .C1(n_2), .C2(n_1), .ZN(n_347));
   INV_X1 i_169 (.A(n_351), .ZN(n_349));
   OAI222_X1 i_170 (.A1(n_10), .A2(n_8), .B1(n_12), .B2(n_16), .C1(n_22), 
      .C2(n_17), .ZN(n_351));
   NOR2_X1 i_171 (.A1(n_22), .A2(n_17), .ZN(n_353));
   AOI221_X1 i_172 (.A(n_357), .B1(p_15[4]), .B2(n_0), .C1(n_2), .C2(n_1), 
      .ZN(n_355));
   INV_X1 i_173 (.A(n_358), .ZN(n_357));
   OAI222_X1 i_174 (.A1(p_0[3]), .A2(p_15[3]), .B1(p_15[4]), .B2(n_0), .C1(n_207), 
      .C2(n_205), .ZN(n_358));
   AOI22_X1 i_175 (.A1(n_30), .A2(n_28), .B1(n_38), .B2(n_31), .ZN(n_359));
   OAI22_X1 i_176 (.A1(n_58), .A2(n_49), .B1(n_38), .B2(n_31), .ZN(n_361));
   NOR2_X1 i_177 (.A1(n_58), .A2(n_49), .ZN(n_362));
   NOR2_X1 i_178 (.A1(n_46), .A2(n_48), .ZN(n_365));
   NAND2_X1 i_179 (.A1(n_161), .A2(n_178), .ZN(n_367));
   INV_X1 i_180 (.A(n_371), .ZN(n_369));
   OAI22_X1 i_181 (.A1(n_391), .A2(n_375), .B1(n_404), .B2(n_373), .ZN(n_371));
   OAI21_X1 i_182 (.A(n_160), .B1(n_161), .B2(n_178), .ZN(n_373));
   AOI22_X1 i_183 (.A1(n_126), .A2(n_111), .B1(n_142), .B2(n_127), .ZN(n_375));
   INV_X1 i_184 (.A(n_391), .ZN(n_390));
   OAI222_X1 i_185 (.A1(n_143), .A2(n_160), .B1(n_161), .B2(n_178), .C1(n_142), 
      .C2(n_127), .ZN(n_391));
   INV_X1 i_186 (.A(n_143), .ZN(n_404));
   FA_X1 i_187 (.A(n_226), .B(n_224), .CI(n_222), .CO(n_233), .S(n_232));
   FA_X1 i_188 (.A(n_265), .B(n_241), .CI(n_219), .CO(n_237), .S(n_236));
   FA_X1 i_189 (.A(n_220), .B(n_230), .CI(n_228), .CO(n_235), .S(n_234));
   FA_X1 i_190 (.A(n_232), .B(n_236), .CI(n_234), .CO(n_239), .S(n_238));
   HA_X1 i_191 (.A(n_267), .B(n_238), .CO(n_407), .S(n_405));
   FA_X1 i_192 (.A(p_0[24]), .B(p_1[24]), .CI(p_2[24]), .CO(n_221), .S(n_220));
   FA_X1 i_193 (.A(n_261), .B(n_263), .CI(n_217), .CO(n_231), .S(n_230));
   FA_X1 i_194 (.A(p_15[24]), .B(n_240), .CI(n_260), .CO(n_229), .S(n_228));
   FA_X1 i_195 (.A(p_5[25]), .B(p_6[25]), .CI(p_7[25]), .CO(n_245), .S(n_244));
   FA_X1 i_196 (.A(p_2[25]), .B(p_3[25]), .CI(p_4[25]), .CO(n_243), .S(n_242));
   FA_X1 i_197 (.A(n_244), .B(n_242), .CI(n_561), .CO(n_253), .S(n_252));
   FA_X1 i_198 (.A(p_8[25]), .B(p_9[25]), .CI(p_10[25]), .CO(n_247), .S(n_246));
   FA_X1 i_199 (.A(n_229), .B(n_558), .CI(n_246), .CO(n_251), .S(n_250));
   FA_X1 i_200 (.A(n_235), .B(n_252), .CI(n_250), .CO(n_257), .S(n_256));
   FA_X1 i_201 (.A(p_6[24]), .B(p_7[24]), .CI(p_8[24]), .CO(n_225), .S(n_224));
   FA_X1 i_202 (.A(p_3[24]), .B(p_4[24]), .CI(p_5[24]), .CO(n_223), .S(n_222));
   FA_X1 i_203 (.A(n_225), .B(n_223), .CI(n_221), .CO(n_249), .S(n_248));
   FA_X1 i_204 (.A(p_9[24]), .B(p_10[24]), .CI(p_11[24]), .CO(n_227), .S(n_226));
   FA_X1 i_205 (.A(n_231), .B(n_248), .CI(n_233), .CO(n_255), .S(n_254));
   FA_X1 i_206 (.A(n_237), .B(n_254), .CI(n_239), .CO(n_259), .S(n_258));
   HA_X1 i_207 (.A(n_256), .B(n_258), .CO(n_411), .S(n_409));
   FA_X1 i_208 (.A(p_11[26]), .B(n_247), .CI(n_245), .CO(n_413), .S(n_268));
   FA_X1 i_209 (.A(n_268), .B(n_253), .CI(n_251), .CO(n_415), .S(n_276));
   FA_X1 i_210 (.A(p_2[26]), .B(p_3[26]), .CI(p_4[26]), .CO(n_417), .S(n_262));
   FA_X1 i_211 (.A(n_243), .B(n_562), .CI(n_249), .CO(n_418), .S(n_270));
   FA_X1 i_212 (.A(n_262), .B(n_554), .CI(n_270), .CO(n_419), .S(n_274));
   FA_X1 i_213 (.A(p_8[26]), .B(p_9[26]), .CI(p_10[26]), .CO(n_430), .S(n_266));
   FA_X1 i_214 (.A(p_5[26]), .B(p_6[26]), .CI(p_7[26]), .CO(n_431), .S(n_264));
   FA_X1 i_215 (.A(n_556), .B(n_266), .CI(n_264), .CO(n_442), .S(n_272));
   FA_X1 i_216 (.A(n_255), .B(n_274), .CI(n_272), .CO(n_445), .S(n_278));
   FA_X1 i_217 (.A(n_276), .B(n_257), .CI(n_278), .CO(n_447), .S(n_280));
   HA_X1 i_218 (.A(n_259), .B(n_280), .CO(n_451), .S(n_449));
   OAI21_X1 i_219 (.A(n_462), .B1(n_505), .B2(n_502), .ZN(n_554));
   XNOR2_X1 i_220 (.A(p_11[25]), .B(n_453), .ZN(n_558));
   OAI22_X1 i_221 (.A1(p_15[32]), .A2(n_494), .B1(n_500), .B2(n_455), .ZN(n_556));
   OAI21_X1 i_222 (.A(n_457), .B1(p_15[32]), .B2(n_494), .ZN(n_453));
   INV_X1 i_223 (.A(n_457), .ZN(n_455));
   NAND2_X1 i_224 (.A1(p_15[32]), .A2(n_494), .ZN(n_457));
   OAI21_X1 i_225 (.A(n_562), .B1(n_503), .B2(n_501), .ZN(n_561));
   NAND2_X1 i_226 (.A1(n_503), .A2(n_501), .ZN(n_562));
   XNOR2_X1 i_227 (.A(n_470), .B(n_459), .ZN(\aggregated_res[14] [26]));
   OAI21_X1 i_228 (.A(n_461), .B1(n_411), .B2(n_449), .ZN(n_459));
   NAND2_X1 i_229 (.A1(n_411), .A2(n_449), .ZN(n_461));
   NAND2_X1 i_230 (.A1(n_505), .A2(n_502), .ZN(n_462));
   INV_X1 i_231 (.A(n_470), .ZN(n_463));
   OAI21_X1 i_232 (.A(n_478), .B1(n_499), .B2(n_471), .ZN(n_470));
   OAI21_X1 i_233 (.A(n_483), .B1(n_213), .B2(n_215), .ZN(n_471));
   AOI221_X1 i_234 (.A(n_481), .B1(n_407), .B2(n_409), .C1(n_490), .C2(n_483), 
      .ZN(n_478));
   NOR2_X1 i_235 (.A1(n_487), .A2(n_485), .ZN(n_481));
   NOR3_X1 i_236 (.A1(n_277), .A2(n_487), .A3(n_489), .ZN(n_483));
   NAND2_X1 i_237 (.A1(n_405), .A2(n_269), .ZN(n_485));
   NOR2_X1 i_238 (.A1(n_407), .A2(n_409), .ZN(n_487));
   NOR2_X1 i_239 (.A1(n_405), .A2(n_269), .ZN(n_489));
   INV_X1 i_240 (.A(n_491), .ZN(n_490));
   AOI21_X1 i_241 (.A(n_275), .B1(n_213), .B2(n_215), .ZN(n_491));
   INV_X1 i_242 (.A(n_227), .ZN(n_494));
   INV_X1 i_243 (.A(n_282), .ZN(n_499));
   INV_X1 i_244 (.A(p_11[25]), .ZN(n_500));
   INV_X1 i_245 (.A(p_1[25]), .ZN(n_501));
   INV_X1 i_246 (.A(p_1[26]), .ZN(n_502));
   INV_X1 i_247 (.A(p_0[25]), .ZN(n_503));
   INV_X1 i_248 (.A(p_0[26]), .ZN(n_505));
   FA_X1 i_249 (.A(n_430), .B(n_431), .CI(n_417), .CO(n_291), .S(n_290));
   FA_X1 i_250 (.A(p_9[28]), .B(p_10[28]), .CI(p_11[28]), .CO(n_309), .S(n_308));
   FA_X1 i_251 (.A(n_553), .B(n_291), .CI(n_308), .CO(n_313), .S(n_312));
   FA_X1 i_252 (.A(n_418), .B(n_290), .CI(n_442), .CO(n_297), .S(n_296));
   FA_X1 i_253 (.A(p_6[28]), .B(p_7[28]), .CI(p_8[28]), .CO(n_307), .S(n_306));
   FA_X1 i_254 (.A(p_3[28]), .B(p_4[28]), .CI(p_5[28]), .CO(n_305), .S(n_304));
   FA_X1 i_255 (.A(n_306), .B(n_304), .CI(n_549), .CO(n_315), .S(n_314));
   FA_X1 i_256 (.A(n_312), .B(n_297), .CI(n_314), .CO(n_319), .S(n_318));
   FA_X1 i_257 (.A(p_4[29]), .B(p_5[29]), .CI(p_6[29]), .CO(n_507), .S(n_324));
   FA_X1 i_258 (.A(n_307), .B(n_305), .CI(n_550), .CO(n_512), .S(n_330));
   FA_X1 i_259 (.A(n_324), .B(n_546), .CI(n_330), .CO(n_515), .S(n_334));
   FA_X1 i_260 (.A(p_9[27]), .B(p_10[27]), .CI(p_11[27]), .CO(n_289), .S(n_288));
   FA_X1 i_261 (.A(p_6[27]), .B(p_7[27]), .CI(p_8[27]), .CO(n_287), .S(n_286));
   FA_X1 i_262 (.A(p_3[27]), .B(p_4[27]), .CI(p_5[27]), .CO(n_285), .S(n_284));
   FA_X1 i_263 (.A(n_289), .B(n_287), .CI(n_285), .CO(n_311), .S(n_310));
   FA_X1 i_264 (.A(p_10[29]), .B(p_11[29]), .CI(n_309), .CO(n_517), .S(n_328));
   FA_X1 i_265 (.A(p_7[29]), .B(p_8[29]), .CI(p_9[29]), .CO(n_522), .S(n_326));
   FA_X1 i_266 (.A(n_311), .B(n_328), .CI(n_326), .CO(n_525), .S(n_332));
   FA_X1 i_267 (.A(n_286), .B(n_284), .CI(n_551), .CO(n_295), .S(n_294));
   FA_X1 i_268 (.A(n_462), .B(n_413), .CI(n_288), .CO(n_293), .S(n_292));
   FA_X1 i_269 (.A(n_310), .B(n_295), .CI(n_293), .CO(n_317), .S(n_316));
   FA_X1 i_270 (.A(n_315), .B(n_313), .CI(n_317), .CO(n_527), .S(n_336));
   FA_X1 i_271 (.A(n_334), .B(n_332), .CI(n_336), .CO(n_532), .S(n_338));
   FA_X1 i_272 (.A(n_292), .B(n_415), .CI(n_419), .CO(n_299), .S(n_298));
   FA_X1 i_273 (.A(n_299), .B(n_316), .CI(n_318), .CO(n_321), .S(n_320));
   FA_X1 i_274 (.A(n_319), .B(n_338), .CI(n_321), .CO(n_537), .S(n_535));
   FA_X1 i_275 (.A(n_294), .B(n_296), .CI(n_445), .CO(n_301), .S(n_300));
   HA_X1 i_276 (.A(n_301), .B(n_320), .CO(n_539), .S(n_322));
   FA_X1 i_277 (.A(n_298), .B(n_300), .CI(n_447), .CO(n_303), .S(n_302));
   XOR2_X1 i_278 (.A(p_2[27]), .B(n_211), .Z(n_551));
   XNOR2_X1 i_279 (.A(p_3[29]), .B(n_540), .ZN(n_546));
   XOR2_X1 i_280 (.A(p_2[29]), .B(p_1[36]), .Z(n_540));
   OAI21_X1 i_281 (.A(n_550), .B1(n_583), .B2(n_578), .ZN(n_549));
   NAND2_X1 i_282 (.A1(n_583), .A2(n_578), .ZN(n_550));
   OAI222_X1 i_283 (.A1(n_577), .A2(p_0[34]), .B1(n_579), .B2(p_0[34]), .C1(
      n_579), .C2(n_577), .ZN(n_553));
   XOR2_X1 i_284 (.A(n_543), .B(n_542), .Z(\aggregated_res[14] [29]));
   AOI21_X1 i_285 (.A(n_574), .B1(n_569), .B2(n_547), .ZN(n_542));
   AOI21_X1 i_286 (.A(n_576), .B1(n_535), .B2(n_539), .ZN(n_543));
   INV_X1 i_287 (.A(n_547), .ZN(n_545));
   OAI21_X1 i_288 (.A(n_560), .B1(n_557), .B2(n_552), .ZN(n_547));
   AOI21_X1 i_289 (.A(n_555), .B1(n_461), .B2(n_463), .ZN(n_552));
   NOR2_X1 i_291 (.A1(n_411), .A2(n_449), .ZN(n_555));
   INV_X1 i_292 (.A(n_559), .ZN(n_557));
   NAND2_X1 i_293 (.A1(n_451), .A2(n_302), .ZN(n_559));
   INV_X1 i_294 (.A(n_565), .ZN(n_560));
   NOR2_X1 i_295 (.A1(n_451), .A2(n_302), .ZN(n_565));
   INV_X1 i_296 (.A(n_569), .ZN(n_568));
   NAND2_X1 i_297 (.A1(n_322), .A2(n_303), .ZN(n_569));
   INV_X1 i_298 (.A(n_574), .ZN(n_572));
   NOR2_X1 i_299 (.A1(n_322), .A2(n_303), .ZN(n_574));
   INV_X1 i_300 (.A(n_576), .ZN(n_575));
   NOR2_X1 i_301 (.A1(n_535), .A2(n_539), .ZN(n_576));
   INV_X1 i_302 (.A(p_1[27]), .ZN(n_577));
   INV_X1 i_303 (.A(p_1[28]), .ZN(n_578));
   INV_X1 i_304 (.A(p_2[27]), .ZN(n_579));
   INV_X1 i_305 (.A(p_2[28]), .ZN(n_583));
   FA_X1 i_306 (.A(p_10[30]), .B(p_11[30]), .CI(n_522), .CO(n_584), .S(n_346));
   FA_X1 i_307 (.A(p_7[30]), .B(p_8[30]), .CI(p_9[30]), .CO(n_585), .S(n_344));
   FA_X1 i_308 (.A(n_517), .B(n_346), .CI(n_344), .CO(n_586), .S(n_350));
   FA_X1 i_309 (.A(p_4[30]), .B(p_5[30]), .CI(p_6[30]), .CO(n_587), .S(n_342));
   FA_X1 i_310 (.A(n_507), .B(n_548), .CI(n_512), .CO(n_588), .S(n_348));
   FA_X1 i_311 (.A(n_342), .B(n_544), .CI(n_348), .CO(n_589), .S(n_352));
   FA_X1 i_312 (.A(n_525), .B(n_515), .CI(n_352), .CO(n_590), .S(n_354));
   FA_X1 i_313 (.A(n_350), .B(n_527), .CI(n_354), .CO(n_591), .S(n_356));
   HA_X1 i_314 (.A(n_532), .B(n_356), .CO(n_595), .S(n_592));
   AOI21_X1 i_315 (.A(n_598), .B1(p_1[36]), .B2(n_597), .ZN(n_548));
   NAND2_X1 i_316 (.A1(p_2[29]), .A2(p_3[29]), .ZN(n_597));
   NOR2_X1 i_317 (.A1(p_2[29]), .A2(p_3[29]), .ZN(n_598));
   OAI21_X1 i_318 (.A(n_601), .B1(n_614), .B2(n_613), .ZN(n_544));
   XNOR2_X1 i_319 (.A(n_603), .B(n_599), .ZN(\aggregated_res[14] [30]));
   OAI21_X1 i_320 (.A(n_600), .B1(n_592), .B2(n_537), .ZN(n_599));
   NAND2_X1 i_321 (.A1(n_592), .A2(n_537), .ZN(n_600));
   NAND2_X1 i_322 (.A1(n_614), .A2(n_613), .ZN(n_601));
   OAI21_X1 i_323 (.A(n_607), .B1(n_463), .B2(n_605), .ZN(n_603));
   OR2_X1 i_324 (.A1(n_555), .A2(n_612), .ZN(n_605));
   INV_X1 i_325 (.A(n_607), .ZN(n_606));
   AOI211_X1 i_326 (.A(n_608), .B(n_609), .C1(n_535), .C2(n_539), .ZN(n_607));
   NOR2_X1 i_327 (.A1(n_576), .A2(n_569), .ZN(n_608));
   AOI21_X1 i_328 (.A(n_612), .B1(n_559), .B2(n_461), .ZN(n_609));
   NAND3_X1 i_329 (.A1(n_560), .A2(n_572), .A3(n_575), .ZN(n_612));
   INV_X1 i_330 (.A(p_3[30]), .ZN(n_613));
   INV_X1 i_331 (.A(p_2[30]), .ZN(n_614));
   FA_X1 i_332 (.A(p_5[31]), .B(p_6[31]), .CI(p_7[31]), .CO(n_615), .S(n_360));
   FA_X1 i_333 (.A(n_360), .B(n_541), .CI(n_588), .CO(n_616), .S(n_368));
   FA_X1 i_334 (.A(p_11[31]), .B(n_585), .CI(n_587), .CO(n_617), .S(n_364));
   FA_X1 i_335 (.A(n_601), .B(n_584), .CI(n_639), .CO(n_618), .S(n_366));
   FA_X1 i_336 (.A(n_364), .B(n_586), .CI(n_366), .CO(n_619), .S(n_370));
   FA_X1 i_337 (.A(n_589), .B(n_368), .CI(n_370), .CO(n_620), .S(n_372));
   FA_X1 i_338 (.A(n_590), .B(n_372), .CI(n_591), .CO(n_621), .S(n_374));
   XOR2_X1 i_339 (.A(n_209), .B(n_201), .Z(n_541));
   INV_X1 i_340 (.A(n_600), .ZN(n_622));
   OAI22_X1 i_341 (.A1(n_622), .A2(n_603), .B1(n_537), .B2(n_592), .ZN(n_623));
   INV_X1 i_342 (.A(n_623), .ZN(n_624));
   NOR2_X1 i_343 (.A1(n_595), .A2(n_374), .ZN(n_625));
   INV_X1 i_344 (.A(n_625), .ZN(n_626));
   AND2_X1 i_345 (.A1(n_595), .A2(n_374), .ZN(n_627));
   NOR2_X1 i_346 (.A1(n_627), .A2(n_625), .ZN(n_628));
   NAND2_X1 i_347 (.A1(n_628), .A2(n_623), .ZN(n_629));
   INV_X1 i_348 (.A(n_629), .ZN(n_630));
   OAI21_X1 i_349 (.A(n_629), .B1(n_623), .B2(n_628), .ZN(
      \aggregated_res[14] [31]));
   FA_X1 i_350 (.A(n_379), .B(n_377), .CI(n_661), .CO(n_397), .S(n_396));
   FA_X1 i_351 (.A(n_203), .B(n_617), .CI(n_378), .CO(n_383), .S(n_382));
   FA_X1 i_352 (.A(n_536), .B(n_396), .CI(n_383), .CO(n_401), .S(n_400));
   FA_X1 i_353 (.A(n_376), .B(n_198), .CI(n_380), .CO(n_385), .S(n_384));
   FA_X1 i_354 (.A(n_618), .B(n_616), .CI(n_382), .CO(n_387), .S(n_386));
   FA_X1 i_355 (.A(n_384), .B(n_619), .CI(n_386), .CO(n_389), .S(n_388));
   FA_X1 i_356 (.A(n_381), .B(n_394), .CI(n_392), .CO(n_399), .S(n_398));
   FA_X1 i_357 (.A(n_385), .B(n_398), .CI(n_387), .CO(n_403), .S(n_402));
   FA_X1 i_358 (.A(n_400), .B(n_389), .CI(n_402), .CO(n_632), .S(n_631));
   HA_X1 i_359 (.A(n_620), .B(n_388), .CO(n_634), .S(n_633));
   FA_X1 i_360 (.A(p_8[32]), .B(p_9[32]), .CI(p_10[32]), .CO(n_379), .S(n_378));
   FA_X1 i_361 (.A(p_5[32]), .B(p_6[32]), .CI(p_7[32]), .CO(n_377), .S(n_376));
   FA_X1 i_362 (.A(p_9[34]), .B(p_10[34]), .CI(p_11[34]), .CO(n_635), .S(n_408));
   FA_X1 i_363 (.A(p_6[34]), .B(p_7[34]), .CI(p_8[34]), .CO(n_636), .S(n_406));
   FA_X1 i_364 (.A(n_397), .B(n_408), .CI(n_406), .CO(n_637), .S(n_412));
   FA_X1 i_365 (.A(p_9[33]), .B(p_10[33]), .CI(p_11[33]), .CO(n_395), .S(n_394));
   FA_X1 i_366 (.A(p_6[33]), .B(p_7[33]), .CI(p_8[33]), .CO(n_393), .S(n_392));
   FA_X1 i_367 (.A(n_395), .B(n_393), .CI(n_538), .CO(n_638), .S(n_410));
   FA_X1 i_368 (.A(p_8[31]), .B(p_9[31]), .CI(p_10[31]), .CO(n_363), .S(n_639));
   FA_X1 i_369 (.A(p_11[32]), .B(n_363), .CI(n_615), .CO(n_381), .S(n_380));
   FA_X1 i_370 (.A(n_534), .B(n_410), .CI(n_399), .CO(n_640), .S(n_414));
   FA_X1 i_371 (.A(n_401), .B(n_412), .CI(n_414), .CO(n_641), .S(n_416));
   HA_X1 i_372 (.A(n_403), .B(n_416), .CO(n_643), .S(n_642));
   OAI222_X1 i_373 (.A1(p_3[40]), .A2(n_663), .B1(n_666), .B2(p_3[40]), .C1(
      n_666), .C2(n_663), .ZN(n_538));
   OAI21_X1 i_374 (.A(n_646), .B1(n_667), .B2(n_664), .ZN(n_534));
   XOR2_X1 i_375 (.A(n_179), .B(n_666), .Z(n_536));
   XOR2_X1 i_376 (.A(n_647), .B(n_644), .Z(\aggregated_res[14] [34]));
   OAI21_X1 i_377 (.A(n_645), .B1(n_632), .B2(n_642), .ZN(n_644));
   NAND2_X1 i_378 (.A1(n_632), .A2(n_642), .ZN(n_645));
   NAND2_X1 i_379 (.A1(n_667), .A2(n_664), .ZN(n_646));
   AND2_X1 i_380 (.A1(n_653), .A2(n_648), .ZN(n_647));
   AOI21_X1 i_381 (.A(n_649), .B1(n_606), .B2(n_654), .ZN(n_648));
   OAI211_X1 i_382 (.A(n_650), .B(n_651), .C1(n_660), .C2(n_652), .ZN(n_649));
   NAND2_X1 i_383 (.A1(n_631), .A2(n_634), .ZN(n_650));
   OAI21_X1 i_384 (.A(n_656), .B1(n_622), .B2(n_627), .ZN(n_651));
   NAND2_X1 i_385 (.A1(n_633), .A2(n_621), .ZN(n_652));
   NAND3_X1 i_386 (.A1(n_668), .A2(n_658), .A3(n_654), .ZN(n_653));
   INV_X1 i_387 (.A(n_655), .ZN(n_654));
   OAI21_X1 i_388 (.A(n_656), .B1(n_592), .B2(n_537), .ZN(n_655));
   NOR2_X1 i_389 (.A1(n_660), .A2(n_657), .ZN(n_656));
   OAI21_X1 i_390 (.A(n_626), .B1(n_633), .B2(n_621), .ZN(n_657));
   OAI21_X1 i_391 (.A(n_478), .B1(n_471), .B2(n_659), .ZN(n_658));
   AND3_X1 i_392 (.A1(n_369), .A2(n_367), .A3(n_283), .ZN(n_659));
   NOR2_X1 i_393 (.A1(n_631), .A2(n_634), .ZN(n_660));
   NAND2_X1 i_394 (.A1(n_665), .A2(n_662), .ZN(n_661));
   INV_X1 i_395 (.A(p_4[32]), .ZN(n_662));
   INV_X1 i_396 (.A(p_4[33]), .ZN(n_663));
   INV_X1 i_397 (.A(p_4[34]), .ZN(n_664));
   INV_X1 i_398 (.A(p_3[32]), .ZN(n_665));
   INV_X1 i_399 (.A(p_5[33]), .ZN(n_666));
   INV_X1 i_400 (.A(p_5[34]), .ZN(n_667));
   INV_X1 i_401 (.A(n_605), .ZN(n_668));
   FA_X1 i_402 (.A(n_636), .B(n_646), .CI(n_638), .CO(n_425), .S(n_424));
   FA_X1 i_403 (.A(n_424), .B(n_637), .CI(n_640), .CO(n_429), .S(n_428));
   FA_X1 i_404 (.A(p_10[35]), .B(p_11[35]), .CI(n_635), .CO(n_423), .S(n_422));
   FA_X1 i_405 (.A(p_7[35]), .B(p_8[35]), .CI(p_9[35]), .CO(n_421), .S(n_420));
   FA_X1 i_406 (.A(n_422), .B(n_420), .CI(n_531), .CO(n_427), .S(n_426));
   FA_X1 i_407 (.A(p_10[36]), .B(p_11[36]), .CI(n_421), .CO(n_435), .S(n_434));
   FA_X1 i_408 (.A(n_533), .B(n_423), .CI(n_434), .CO(n_437), .S(n_436));
   FA_X1 i_409 (.A(p_7[36]), .B(p_8[36]), .CI(p_9[36]), .CO(n_433), .S(n_432));
   FA_X1 i_410 (.A(n_432), .B(n_529), .CI(n_425), .CO(n_439), .S(n_438));
   FA_X1 i_411 (.A(n_427), .B(n_436), .CI(n_438), .CO(n_441), .S(n_440));
   HA_X1 i_412 (.A(n_429), .B(n_440), .CO(n_443), .S(n_669));
   FA_X1 i_413 (.A(p_8[37]), .B(p_9[37]), .CI(p_10[37]), .CO(n_670), .S(n_444));
   FA_X1 i_414 (.A(n_435), .B(n_444), .CI(n_526), .CO(n_671), .S(n_448));
   FA_X1 i_415 (.A(p_11[37]), .B(n_433), .CI(n_530), .CO(n_672), .S(n_446));
   FA_X1 i_416 (.A(n_446), .B(n_437), .CI(n_439), .CO(n_673), .S(n_450));
   FA_X1 i_417 (.A(n_448), .B(n_450), .CI(n_441), .CO(n_674), .S(n_452));
   FA_X1 i_418 (.A(n_426), .B(n_428), .CI(n_641), .CO(n_676), .S(n_675));
   XNOR2_X1 i_419 (.A(p_7[37]), .B(n_677), .ZN(n_526));
   XOR2_X1 i_420 (.A(p_6[37]), .B(p_5[43]), .Z(n_677));
   OAI21_X1 i_421 (.A(n_530), .B1(n_696), .B2(n_694), .ZN(n_529));
   NAND2_X1 i_422 (.A1(n_696), .A2(n_694), .ZN(n_530));
   NAND2_X1 i_423 (.A1(n_681), .A2(n_678), .ZN(n_533));
   NAND2_X1 i_424 (.A1(p_6[35]), .A2(n_680), .ZN(n_678));
   XNOR2_X1 i_425 (.A(p_6[35]), .B(n_679), .ZN(n_531));
   NAND2_X1 i_426 (.A1(n_681), .A2(n_680), .ZN(n_679));
   OR2_X1 i_427 (.A1(n_695), .A2(p_5[35]), .ZN(n_680));
   NAND2_X1 i_428 (.A1(n_695), .A2(p_5[35]), .ZN(n_681));
   XOR2_X1 i_429 (.A(n_683), .B(n_682), .Z(\aggregated_res[14] [37]));
   OAI22_X1 i_430 (.A1(n_669), .A2(n_676), .B1(n_690), .B2(n_684), .ZN(n_682));
   OAI21_X1 i_431 (.A(n_692), .B1(n_443), .B2(n_452), .ZN(n_683));
   AOI21_X1 i_432 (.A(n_689), .B1(n_688), .B2(n_686), .ZN(n_684));
   INV_X1 i_433 (.A(n_686), .ZN(n_685));
   OAI21_X1 i_434 (.A(n_687), .B1(n_632), .B2(n_642), .ZN(n_686));
   NAND2_X1 i_435 (.A1(n_647), .A2(n_645), .ZN(n_687));
   NAND2_X1 i_436 (.A1(n_675), .A2(n_643), .ZN(n_688));
   NOR2_X1 i_437 (.A1(n_675), .A2(n_643), .ZN(n_689));
   INV_X1 i_438 (.A(n_691), .ZN(n_690));
   NAND2_X1 i_439 (.A1(n_669), .A2(n_676), .ZN(n_691));
   NAND2_X1 i_440 (.A1(n_443), .A2(n_452), .ZN(n_692));
   NOR2_X1 i_441 (.A1(n_443), .A2(n_452), .ZN(n_693));
   INV_X1 i_442 (.A(p_5[36]), .ZN(n_694));
   INV_X1 i_443 (.A(p_4[42]), .ZN(n_695));
   INV_X1 i_444 (.A(p_6[36]), .ZN(n_696));
   INV_X1 i_445 (.A(p_7[37]), .ZN(n_697));
   FA_X1 i_446 (.A(p_8[38]), .B(p_9[38]), .CI(p_10[38]), .CO(n_698), .S(n_454));
   FA_X1 i_447 (.A(n_672), .B(n_454), .CI(n_524), .CO(n_699), .S(n_458));
   FA_X1 i_448 (.A(p_11[38]), .B(n_670), .CI(n_528), .CO(n_700), .S(n_456));
   FA_X1 i_449 (.A(n_456), .B(n_671), .CI(n_673), .CO(n_701), .S(n_460));
   HA_X1 i_450 (.A(n_458), .B(n_460), .CO(n_703), .S(n_702));
   INV_X1 i_451 (.A(p_6[37]), .ZN(n_704));
   OAI222_X1 i_452 (.A1(n_704), .A2(n_697), .B1(n_704), .B2(p_5[43]), .C1(
      p_5[43]), .C2(n_697), .ZN(n_528));
   INV_X1 i_453 (.A(p_6[38]), .ZN(n_705));
   INV_X1 i_454 (.A(p_7[38]), .ZN(n_706));
   NAND2_X1 i_457 (.A1(n_705), .A2(n_706), .ZN(n_707));
   OAI21_X1 i_458 (.A(n_707), .B1(n_705), .B2(n_706), .ZN(n_524));
   NOR2_X1 i_459 (.A1(n_676), .A2(n_669), .ZN(n_708));
   NOR3_X1 i_460 (.A1(n_708), .A2(n_689), .A3(n_693), .ZN(n_709));
   OAI21_X1 i_461 (.A(n_709), .B1(n_632), .B2(n_642), .ZN(n_710));
   AOI21_X1 i_462 (.A(n_710), .B1(n_653), .B2(n_648), .ZN(n_711));
   INV_X1 i_463 (.A(n_709), .ZN(n_712));
   AND2_X1 i_464 (.A1(n_645), .A2(n_688), .ZN(n_713));
   OAI221_X1 i_465 (.A(n_692), .B1(n_693), .B2(n_691), .C1(n_712), .C2(n_713), 
      .ZN(n_714));
   NOR2_X1 i_466 (.A1(n_714), .A2(n_711), .ZN(n_715));
   NAND2_X1 i_467 (.A1(n_702), .A2(n_674), .ZN(n_716));
   OAI21_X1 i_468 (.A(n_716), .B1(n_702), .B2(n_674), .ZN(n_717));
   XOR2_X1 i_469 (.A(n_715), .B(n_717), .Z(\aggregated_res[14] [38]));
   FA_X1 i_470 (.A(p_9[39]), .B(p_10[39]), .CI(p_11[39]), .CO(n_465), .S(n_464));
   FA_X1 i_471 (.A(n_698), .B(n_707), .CI(n_700), .CO(n_467), .S(n_466));
   FA_X1 i_472 (.A(n_464), .B(n_521), .CI(n_466), .CO(n_469), .S(n_468));
   FA_X1 i_473 (.A(p_9[40]), .B(p_10[40]), .CI(p_11[40]), .CO(n_473), .S(n_472));
   FA_X1 i_474 (.A(n_465), .B(n_523), .CI(n_472), .CO(n_475), .S(n_474));
   FA_X1 i_475 (.A(n_519), .B(n_467), .CI(n_474), .CO(n_477), .S(n_476));
   HA_X1 i_476 (.A(n_469), .B(n_476), .CO(n_479), .S(n_718));
   FA_X1 i_477 (.A(p_10[41]), .B(p_11[41]), .CI(n_473), .CO(n_719), .S(n_480));
   FA_X1 i_478 (.A(n_520), .B(n_480), .CI(n_516), .CO(n_720), .S(n_482));
   FA_X1 i_479 (.A(n_475), .B(n_477), .CI(n_482), .CO(n_721), .S(n_484));
   FA_X1 i_480 (.A(n_699), .B(n_468), .CI(n_701), .CO(n_723), .S(n_722));
   XNOR2_X1 i_481 (.A(p_9[41]), .B(n_724), .ZN(n_516));
   XOR2_X1 i_482 (.A(p_8[41]), .B(p_7[45]), .Z(n_724));
   NAND2_X1 i_483 (.A1(n_728), .A2(n_725), .ZN(n_523));
   NAND2_X1 i_484 (.A1(p_8[39]), .A2(n_727), .ZN(n_725));
   OAI21_X1 i_485 (.A(n_520), .B1(n_744), .B2(n_742), .ZN(n_519));
   NAND2_X1 i_486 (.A1(n_744), .A2(n_742), .ZN(n_520));
   XNOR2_X1 i_487 (.A(p_8[39]), .B(n_726), .ZN(n_521));
   NAND2_X1 i_488 (.A1(n_728), .A2(n_727), .ZN(n_726));
   OR2_X1 i_489 (.A1(n_743), .A2(p_7[39]), .ZN(n_727));
   NAND2_X1 i_490 (.A1(n_743), .A2(p_7[39]), .ZN(n_728));
   XOR2_X1 i_491 (.A(n_730), .B(n_729), .Z(\aggregated_res[14] [41]));
   OAI22_X1 i_492 (.A1(n_718), .A2(n_723), .B1(n_737), .B2(n_731), .ZN(n_729));
   OAI21_X1 i_493 (.A(n_740), .B1(n_479), .B2(n_484), .ZN(n_730));
   AOI21_X1 i_494 (.A(n_736), .B1(n_735), .B2(n_733), .ZN(n_731));
   INV_X1 i_495 (.A(n_733), .ZN(n_732));
   OAI21_X1 i_496 (.A(n_734), .B1(n_702), .B2(n_674), .ZN(n_733));
   NAND2_X1 i_497 (.A1(n_715), .A2(n_716), .ZN(n_734));
   NAND2_X1 i_498 (.A1(n_722), .A2(n_703), .ZN(n_735));
   NOR2_X1 i_499 (.A1(n_722), .A2(n_703), .ZN(n_736));
   INV_X1 i_500 (.A(n_738), .ZN(n_737));
   NAND2_X1 i_501 (.A1(n_718), .A2(n_723), .ZN(n_738));
   NAND2_X1 i_502 (.A1(n_479), .A2(n_484), .ZN(n_740));
   NOR2_X1 i_503 (.A1(n_479), .A2(n_484), .ZN(n_741));
   INV_X1 i_504 (.A(p_7[40]), .ZN(n_742));
   INV_X1 i_505 (.A(p_6[45]), .ZN(n_743));
   INV_X1 i_506 (.A(p_8[40]), .ZN(n_744));
   INV_X1 i_507 (.A(p_9[41]), .ZN(n_745));
   FA_X1 i_508 (.A(p_10[42]), .B(p_11[42]), .CI(n_518), .CO(n_746), .S(n_486));
   FA_X1 i_509 (.A(n_719), .B(n_486), .CI(n_514), .CO(n_747), .S(n_488));
   HA_X1 i_510 (.A(n_720), .B(n_488), .CO(n_749), .S(n_748));
   INV_X1 i_511 (.A(p_8[42]), .ZN(n_750));
   INV_X1 i_512 (.A(p_9[42]), .ZN(n_751));
   NAND2_X1 i_513 (.A1(n_750), .A2(n_751), .ZN(n_752));
   OAI21_X1 i_514 (.A(n_752), .B1(n_750), .B2(n_751), .ZN(n_514));
   INV_X1 i_515 (.A(p_8[41]), .ZN(n_753));
   OAI222_X1 i_516 (.A1(n_753), .A2(n_745), .B1(n_753), .B2(p_7[45]), .C1(
      p_7[45]), .C2(n_745), .ZN(n_518));
   NOR2_X1 i_517 (.A1(n_723), .A2(n_718), .ZN(n_754));
   OR3_X1 i_518 (.A1(n_754), .A2(n_736), .A3(n_741), .ZN(n_755));
   OAI22_X1 i_519 (.A1(n_711), .A2(n_714), .B1(n_674), .B2(n_702), .ZN(n_756));
   AND3_X1 i_520 (.A1(n_756), .A2(n_735), .A3(n_716), .ZN(n_757));
   OAI221_X1 i_521 (.A(n_740), .B1(n_741), .B2(n_738), .C1(n_755), .C2(n_757), 
      .ZN(n_758));
   NAND2_X1 i_522 (.A1(n_748), .A2(n_721), .ZN(n_759));
   OAI21_X1 i_523 (.A(n_759), .B1(n_748), .B2(n_721), .ZN(n_760));
   XNOR2_X1 i_524 (.A(n_758), .B(n_760), .ZN(\aggregated_res[14] [42]));
   INV_X1 i_525 (.A(n_758), .ZN(n_761));
   FA_X1 i_526 (.A(p_11[43]), .B(n_752), .CI(n_746), .CO(n_493), .S(n_492));
   FA_X1 i_527 (.A(p_11[44]), .B(n_513), .CI(n_509), .CO(n_497), .S(n_496));
   HA_X1 i_528 (.A(n_493), .B(n_496), .CO(n_762), .S(n_498));
   FA_X1 i_529 (.A(n_510), .B(n_506), .CI(n_497), .CO(n_764), .S(n_763));
   FA_X1 i_530 (.A(n_511), .B(n_492), .CI(n_747), .CO(n_495), .S(n_765));
   XNOR2_X1 i_531 (.A(n_788), .B(n_766), .ZN(n_511));
   AOI21_X1 i_532 (.A(n_769), .B1(n_785), .B2(p_8[45]), .ZN(n_766));
   XNOR2_X1 i_533 (.A(p_11[45]), .B(n_767), .ZN(n_506));
   XOR2_X1 i_534 (.A(p_10[45]), .B(p_9[45]), .Z(n_767));
   OAI21_X1 i_535 (.A(n_510), .B1(n_789), .B2(n_787), .ZN(n_509));
   NAND2_X1 i_536 (.A1(n_789), .A2(n_787), .ZN(n_510));
   AOI22_X1 i_537 (.A1(n_785), .A2(p_8[45]), .B1(n_788), .B2(n_768), .ZN(n_513));
   INV_X1 i_538 (.A(n_769), .ZN(n_768));
   NOR2_X1 i_539 (.A1(n_785), .A2(p_8[45]), .ZN(n_769));
   XNOR2_X1 i_540 (.A(n_772), .B(n_770), .ZN(\aggregated_res[14] [45]));
   NAND2_X1 i_541 (.A1(n_780), .A2(n_771), .ZN(n_770));
   OAI21_X1 i_542 (.A(n_773), .B1(n_781), .B2(n_777), .ZN(n_771));
   OAI21_X1 i_543 (.A(n_783), .B1(n_762), .B2(n_763), .ZN(n_772));
   NOR2_X1 i_544 (.A1(n_776), .A2(n_774), .ZN(n_773));
   NOR2_X1 i_545 (.A1(n_498), .A2(n_495), .ZN(n_774));
   NOR2_X1 i_546 (.A1(n_777), .A2(n_776), .ZN(n_775));
   NOR2_X1 i_547 (.A1(n_765), .A2(n_749), .ZN(n_776));
   INV_X1 i_548 (.A(n_778), .ZN(n_777));
   NAND2_X1 i_549 (.A1(n_765), .A2(n_749), .ZN(n_778));
   INV_X1 i_550 (.A(n_780), .ZN(n_779));
   NAND2_X1 i_551 (.A1(n_498), .A2(n_495), .ZN(n_780));
   AOI21_X1 i_552 (.A(n_782), .B1(n_761), .B2(n_759), .ZN(n_781));
   NOR2_X1 i_553 (.A1(n_721), .A2(n_748), .ZN(n_782));
   NAND2_X1 i_554 (.A1(n_762), .A2(n_763), .ZN(n_783));
   NOR2_X1 i_555 (.A1(n_762), .A2(n_763), .ZN(n_784));
   INV_X1 i_556 (.A(p_9[43]), .ZN(n_785));
   INV_X1 i_557 (.A(p_9[44]), .ZN(n_787));
   INV_X1 i_558 (.A(p_10[43]), .ZN(n_788));
   INV_X1 i_559 (.A(p_10[44]), .ZN(n_789));
   INV_X1 i_560 (.A(p_11[45]), .ZN(n_790));
   HA_X1 i_561 (.A(n_508), .B(n_504), .CO(n_792), .S(n_791));
   INV_X1 i_562 (.A(n_793), .ZN(n_504));
   AOI21_X1 i_563 (.A(n_796), .B1(p_10[46]), .B2(p_11[46]), .ZN(n_793));
   OAI222_X1 i_564 (.A1(p_9[45]), .A2(n_790), .B1(n_804), .B2(p_9[45]), .C1(
      n_804), .C2(n_790), .ZN(n_508));
   XNOR2_X1 i_565 (.A(n_795), .B(n_794), .ZN(\aggregated_res[14] [46]));
   OAI22_X1 i_566 (.A1(n_805), .A2(n_764), .B1(n_791), .B2(n_803), .ZN(n_794));
   AOI21_X1 i_567 (.A(n_799), .B1(n_758), .B2(n_797), .ZN(n_795));
   NOR2_X1 i_568 (.A1(p_10[46]), .A2(p_11[46]), .ZN(n_796));
   NOR2_X1 i_569 (.A1(n_802), .A2(n_798), .ZN(n_797));
   NOR2_X1 i_570 (.A1(n_721), .A2(n_748), .ZN(n_798));
   OAI211_X1 i_571 (.A(n_783), .B(n_800), .C1(n_780), .C2(n_784), .ZN(n_799));
   INV_X1 i_572 (.A(n_801), .ZN(n_800));
   AOI21_X1 i_573 (.A(n_802), .B1(n_759), .B2(n_778), .ZN(n_801));
   OAI21_X1 i_574 (.A(n_773), .B1(n_762), .B2(n_763), .ZN(n_802));
   INV_X1 i_575 (.A(n_764), .ZN(n_803));
   INV_X1 i_576 (.A(p_10[45]), .ZN(n_804));
   INV_X1 i_577 (.A(n_791), .ZN(n_805));
   XOR2_X1 i_578 (.A(n_809), .B(n_806), .Z(\aggregated_res[14] [47]));
   XOR2_X1 i_579 (.A(n_792), .B(n_807), .Z(n_806));
   XOR2_X1 i_580 (.A(n_796), .B(n_808), .Z(n_807));
   XOR2_X1 i_581 (.A(p_10[47]), .B(p_11[47]), .Z(n_808));
   NOR2_X1 i_582 (.A1(n_812), .A2(n_810), .ZN(n_809));
   AOI211_X1 i_583 (.A(n_811), .B(n_799), .C1(n_758), .C2(n_797), .ZN(n_810));
   NOR2_X1 i_584 (.A1(n_805), .A2(n_803), .ZN(n_811));
   NOR2_X1 i_585 (.A1(n_791), .A2(n_764), .ZN(n_812));
endmodule

module boothAlgoR4(Res, OVF, A, B, clk, reset, enable);
   output [63:0]Res;
   output OVF;
   input [31:0]A;
   input [31:0]B;
   input clk;
   input reset;
   input enable;

   wire [31:0]A_imm_2s_complement;
   wire [63:0]\aggregated_res[14] ;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_32;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_58;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_89;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_122;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_153;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_184;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_215;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_246;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_277;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_302;
   wire n_0_303;
   wire n_0_308;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_335;
   wire n_0_339;
   wire n_0_344;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_363;
   wire n_0_365;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_386;
   wire n_0_388;
   wire n_0_391;
   wire n_0_385;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_33;
   wire n_0_34;
   wire n_0_57;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_88;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_202;
   wire n_0_206;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_268;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_301;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_330;
   wire n_0_334;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_345;
   wire n_0_358;
   wire n_0_362;
   wire n_0_364;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_381;
   wire n_0_387;
   wire n_0_389;
   wire n_0_390;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_1_0__0;
   wire n_1_0__1;

   datapath__0_0 i_2 (.A_imm({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, 
      n_46, n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, 
      n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22}), 
      .A_imm_2s_complement({uc_8, uc_9, uc_10, uc_11, A_imm_2s_complement[27], 
      uc_12, uc_13, uc_14, A_imm_2s_complement[23], A_imm_2s_complement[22], 
      A_imm_2s_complement[21], A_imm_2s_complement[20], A_imm_2s_complement[19], 
      A_imm_2s_complement[18], A_imm_2s_complement[17], A_imm_2s_complement[16], 
      A_imm_2s_complement[15], A_imm_2s_complement[14], A_imm_2s_complement[13], 
      A_imm_2s_complement[12], A_imm_2s_complement[11], A_imm_2s_complement[10], 
      A_imm_2s_complement[9], A_imm_2s_complement[8], A_imm_2s_complement[7], 
      A_imm_2s_complement[6], A_imm_2s_complement[5], A_imm_2s_complement[4], 
      A_imm_2s_complement[3], A_imm_2s_complement[2], A_imm_2s_complement[1], 
      uc_15}));
   datapath__0_67 i_53 (.p_0({uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, 
      uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, uc_32, 
      uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, 
      uc_43, uc_44, n_361, uc_45, uc_46, uc_47, uc_48, uc_49, uc_50, uc_51, 
      n_360, n_359, n_379, n_358, n_357, n_356, n_378, n_355, n_354, n_353, 
      n_352, n_351, n_350, n_349, n_348, n_347, n_346, n_345, n_344, n_343, 
      n_342, n_341, n_340, n_377, n_339, uc_52, uc_53}), .p_1({uc_54, uc_55, 
      uc_56, uc_57, uc_58, uc_59, uc_60, uc_61, uc_62, uc_63, uc_64, uc_65, 
      uc_66, uc_67, uc_68, uc_69, uc_70, uc_71, uc_72, uc_73, uc_74, uc_75, 
      uc_76, uc_77, uc_78, uc_79, uc_80, n_338, uc_81, uc_82, uc_83, uc_84, 
      uc_85, uc_86, uc_87, n_337, n_376, n_336, n_335, n_375, n_334, n_333, 
      n_332, n_331, n_330, n_329, n_328, n_327, n_326, n_325, n_324, n_323, 
      n_322, n_321, n_320, n_319, n_318, n_317, n_374, n_316, uc_88, uc_89, 
      uc_90, uc_91}), .p_2({uc_92, uc_93, uc_94, uc_95, uc_96, uc_97, uc_98, 
      uc_99, uc_100, uc_101, uc_102, uc_103, uc_104, uc_105, uc_106, uc_107, 
      uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, uc_114, uc_115, uc_116, 
      n_315, uc_117, uc_118, uc_119, uc_120, uc_121, uc_122, uc_123, n_314, 
      n_313, n_312, n_311, n_310, n_309, n_373, n_308, n_307, n_306, n_305, 
      n_304, n_303, n_302, n_301, n_300, n_299, n_298, n_297, n_296, n_295, 
      n_294, n_293, n_372, n_292, uc_124, uc_125, uc_126, uc_127, uc_128, uc_129}), 
      .p_3({uc_130, uc_131, uc_132, uc_133, uc_134, uc_135, uc_136, uc_137, 
      uc_138, uc_139, uc_140, uc_141, uc_142, uc_143, uc_144, uc_145, uc_146, 
      uc_147, uc_148, uc_149, uc_150, uc_151, uc_152, n_291, uc_153, uc_154, 
      uc_155, uc_156, uc_157, uc_158, uc_159, n_290, n_289, n_288, n_287, n_286, 
      n_285, n_284, n_283, n_282, n_281, n_280, n_279, n_278, n_277, n_276, 
      n_275, n_274, n_273, n_272, n_271, n_270, n_269, n_268, n_371, n_267, 
      uc_160, uc_161, uc_162, uc_163, uc_164, uc_165, uc_166, uc_167}), .p_4({
      uc_168, uc_169, uc_170, uc_171, uc_172, uc_173, uc_174, uc_175, uc_176, 
      uc_177, uc_178, uc_179, uc_180, uc_181, uc_182, uc_183, uc_184, uc_185, 
      uc_186, uc_187, uc_188, n_266, uc_189, uc_190, uc_191, uc_192, uc_193, 
      uc_194, uc_195, n_265, n_264, n_263, n_262, n_261, n_260, n_370, n_259, 
      n_258, n_257, n_369, n_256, n_255, n_254, n_253, n_252, n_251, n_250, 
      n_249, n_248, n_247, n_246, n_245, n_368, n_244, uc_196, uc_197, uc_198, 
      uc_199, uc_200, uc_201, uc_202, uc_203, uc_204, uc_205}), .p_5({uc_206, 
      uc_207, uc_208, uc_209, uc_210, uc_211, uc_212, uc_213, uc_214, uc_215, 
      uc_216, uc_217, uc_218, uc_219, uc_220, uc_221, uc_222, uc_223, uc_224, 
      uc_225, n_243, uc_226, uc_227, uc_228, uc_229, uc_230, uc_231, n_242, 
      n_241, n_240, n_239, n_238, n_237, n_236, n_235, n_234, n_233, n_232, 
      n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, n_222, 
      n_221, n_220, n_367, n_219, uc_232, uc_233, uc_234, uc_235, uc_236, uc_237, 
      uc_238, uc_239, uc_240, uc_241, uc_242, uc_243}), .p_6({uc_244, uc_245, 
      uc_246, uc_247, uc_248, uc_249, uc_250, uc_251, uc_252, uc_253, uc_254, 
      uc_255, uc_256, uc_257, uc_258, uc_259, uc_260, uc_261, n_218, uc_262, 
      uc_263, uc_264, uc_265, uc_266, uc_267, n_217, n_216, n_215, n_214, n_213, 
      n_212, n_211, n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, 
      n_202, n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_366, n_194, 
      uc_268, uc_269, uc_270, uc_271, uc_272, uc_273, uc_274, uc_275, uc_276, 
      uc_277, uc_278, uc_279, uc_280, uc_281}), .p_7({uc_282, uc_283, uc_284, 
      uc_285, uc_286, uc_287, uc_288, uc_289, uc_290, uc_291, uc_292, uc_293, 
      uc_294, uc_295, uc_296, uc_297, uc_298, uc_299, n_193, uc_300, uc_301, 
      uc_302, uc_303, n_192, n_191, n_190, n_189, n_188, n_187, n_186, n_185, 
      n_184, n_183, n_182, n_181, n_180, n_179, n_178, n_177, n_176, n_175, 
      n_174, n_173, n_172, n_171, n_170, n_365, n_169, uc_304, uc_305, uc_306, 
      uc_307, uc_308, uc_309, uc_310, uc_311, uc_312, uc_313, uc_314, uc_315, 
      uc_316, uc_317, uc_318, uc_319}), .p_8({uc_320, uc_321, uc_322, uc_323, 
      uc_324, uc_325, uc_326, uc_327, uc_328, uc_329, uc_330, uc_331, uc_332, 
      uc_333, uc_334, uc_335, uc_336, uc_337, n_168, uc_338, uc_339, n_167, 
      n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, n_157, 
      n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, n_147, 
      n_146, n_145, n_364, n_144, uc_340, uc_341, uc_342, uc_343, uc_344, uc_345, 
      uc_346, uc_347, uc_348, uc_349, uc_350, uc_351, uc_352, uc_353, uc_354, 
      uc_355, uc_356, uc_357}), .p_9({uc_358, uc_359, uc_360, uc_361, uc_362, 
      uc_363, uc_364, uc_365, uc_366, uc_367, uc_368, uc_369, uc_370, uc_371, 
      uc_372, uc_373, uc_374, uc_375, n_143, n_142, n_141, n_140, n_139, n_138, 
      n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, n_129, n_128, 
      n_127, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_363, n_119, 
      uc_376, uc_377, uc_378, uc_379, uc_380, uc_381, uc_382, uc_383, uc_384, 
      uc_385, uc_386, uc_387, uc_388, uc_389, uc_390, uc_391, uc_392, uc_393, 
      uc_394, uc_395}), .p_10({uc_396, uc_397, uc_398, uc_399, uc_400, uc_401, 
      uc_402, uc_403, uc_404, uc_405, uc_406, uc_407, uc_408, uc_409, uc_410, 
      uc_411, n_118, n_117, n_362, n_116, n_115, n_114, n_113, n_112, n_111, 
      n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, 
      n_100, n_99, n_98, n_97, n_96, n_95, n_94, uc_412, uc_413, uc_414, uc_415, 
      uc_416, uc_417, uc_418, uc_419, uc_420, uc_421, uc_422, uc_423, uc_424, 
      uc_425, uc_426, uc_427, uc_428, uc_429, uc_430, uc_431, uc_432, uc_433}), 
      .p_11({uc_434, uc_435, uc_436, uc_437, uc_438, uc_439, uc_440, uc_441, 
      uc_442, uc_443, uc_444, uc_445, uc_446, uc_447, uc_448, uc_449, n_46, n_93, 
      n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, 
      n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, uc_450, uc_451, 
      uc_452, uc_453, uc_454, uc_455, uc_456, uc_457, uc_458, uc_459, uc_460, 
      uc_461, uc_462, uc_463, uc_464, uc_465, uc_466, uc_467, uc_468, uc_469, 
      uc_470, uc_471, uc_472, uc_473}), .p_12(), .p_13(), .p_14(), .p_15({uc_474, 
      uc_475, uc_476, uc_477, uc_478, uc_479, uc_480, uc_481, uc_482, uc_483, 
      uc_484, uc_485, uc_486, uc_487, uc_488, uc_489, uc_490, uc_491, uc_492, 
      uc_493, uc_494, uc_495, uc_496, uc_497, uc_498, uc_499, uc_500, uc_501, 
      uc_502, uc_503, uc_504, n_70, uc_505, uc_506, uc_507, uc_508, uc_509, 
      uc_510, uc_511, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, 
      n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, 
      n_47, uc_512, uc_513}), .\aggregated_res[14] ({uc_514, uc_515, uc_516, 
      uc_517, uc_518, uc_519, uc_520, uc_521, uc_522, uc_523, uc_524, uc_525, 
      uc_526, uc_527, uc_528, uc_529, \aggregated_res[14] [47], 
      \aggregated_res[14] [46], \aggregated_res[14] [45], 
      \aggregated_res[14] [44], \aggregated_res[14] [43], 
      \aggregated_res[14] [42], \aggregated_res[14] [41], 
      \aggregated_res[14] [40], \aggregated_res[14] [39], 
      \aggregated_res[14] [38], \aggregated_res[14] [37], 
      \aggregated_res[14] [36], \aggregated_res[14] [35], 
      \aggregated_res[14] [34], \aggregated_res[14] [33], 
      \aggregated_res[14] [32], \aggregated_res[14] [31], 
      \aggregated_res[14] [30], \aggregated_res[14] [29], 
      \aggregated_res[14] [28], \aggregated_res[14] [27], 
      \aggregated_res[14] [26], \aggregated_res[14] [25], 
      \aggregated_res[14] [24], \aggregated_res[14] [23], uc_530, uc_531, uc_532, 
      uc_533, uc_534, uc_535, uc_536, uc_537, uc_538, uc_539, uc_540, uc_541, 
      uc_542, uc_543, uc_544, uc_545, uc_546, uc_547, uc_548, uc_549, uc_550, 
      uc_551, uc_552}));
   DLH_X1 \Res_reg[47]  (.D(n_404), .G(n_452), .Q(Res[47]));
   DLH_X1 \Res_reg[46]  (.D(n_403), .G(n_452), .Q(Res[46]));
   DLH_X1 \Res_reg[45]  (.D(n_402), .G(n_452), .Q(Res[45]));
   DLH_X1 \Res_reg[44]  (.D(n_401), .G(n_452), .Q(Res[44]));
   DLH_X1 \Res_reg[43]  (.D(n_400), .G(n_452), .Q(Res[43]));
   DLH_X1 \Res_reg[42]  (.D(n_399), .G(n_452), .Q(Res[42]));
   DLH_X1 \Res_reg[41]  (.D(n_398), .G(n_452), .Q(Res[41]));
   DLH_X1 \Res_reg[40]  (.D(n_397), .G(n_452), .Q(Res[40]));
   DLH_X1 \Res_reg[39]  (.D(n_396), .G(n_452), .Q(Res[39]));
   DLH_X1 \Res_reg[38]  (.D(n_395), .G(n_452), .Q(Res[38]));
   DLH_X1 \Res_reg[37]  (.D(n_394), .G(n_452), .Q(Res[37]));
   DLH_X1 \Res_reg[36]  (.D(n_393), .G(n_452), .Q(Res[36]));
   DLH_X1 \Res_reg[35]  (.D(n_392), .G(n_452), .Q(Res[35]));
   DLH_X1 \Res_reg[34]  (.D(n_391), .G(n_452), .Q(Res[34]));
   DLH_X1 \Res_reg[33]  (.D(n_390), .G(n_452), .Q(Res[33]));
   DLH_X1 \Res_reg[32]  (.D(n_389), .G(n_452), .Q(Res[32]));
   DLH_X1 \Res_reg[31]  (.D(n_388), .G(n_452), .Q(Res[31]));
   DLH_X1 \Res_reg[30]  (.D(n_387), .G(n_452), .Q(Res[30]));
   DLH_X1 \Res_reg[29]  (.D(n_386), .G(n_452), .Q(Res[29]));
   DLH_X1 \Res_reg[28]  (.D(n_385), .G(n_452), .Q(Res[28]));
   DLH_X1 \Res_reg[27]  (.D(n_384), .G(n_452), .Q(Res[27]));
   DLH_X1 \Res_reg[26]  (.D(n_383), .G(n_452), .Q(Res[26]));
   DLH_X1 \Res_reg[25]  (.D(n_382), .G(n_452), .Q(Res[25]));
   DLH_X1 \Res_reg[24]  (.D(n_381), .G(n_452), .Q(Res[24]));
   DLH_X1 \Res_reg[23]  (.D(n_380), .G(n_452), .Q(Res[23]));
   DLH_X1 \A_in_reg[22]  (.D(n_451), .G(n_428), .Q(n_0));
   DLH_X1 \A_in_reg[21]  (.D(n_450), .G(n_428), .Q(n_1));
   DLH_X1 \A_in_reg[20]  (.D(n_449), .G(n_428), .Q(n_2));
   DLH_X1 \A_in_reg[19]  (.D(n_448), .G(n_428), .Q(n_3));
   DLH_X1 \A_in_reg[18]  (.D(n_447), .G(n_428), .Q(n_4));
   DLH_X1 \A_in_reg[17]  (.D(n_446), .G(n_428), .Q(n_5));
   DLH_X1 \A_in_reg[16]  (.D(n_445), .G(n_428), .Q(n_6));
   DLH_X1 \A_in_reg[15]  (.D(n_444), .G(n_428), .Q(n_7));
   DLH_X1 \A_in_reg[14]  (.D(n_443), .G(n_428), .Q(n_8));
   DLH_X1 \A_in_reg[13]  (.D(n_442), .G(n_428), .Q(n_9));
   DLH_X1 \A_in_reg[12]  (.D(n_441), .G(n_428), .Q(n_10));
   DLH_X1 \A_in_reg[11]  (.D(n_440), .G(n_428), .Q(n_11));
   DLH_X1 \A_in_reg[10]  (.D(n_439), .G(n_428), .Q(n_12));
   DLH_X1 \A_in_reg[9]  (.D(n_438), .G(n_428), .Q(n_13));
   DLH_X1 \A_in_reg[8]  (.D(n_437), .G(n_428), .Q(n_14));
   DLH_X1 \A_in_reg[7]  (.D(n_436), .G(n_428), .Q(n_15));
   DLH_X1 \A_in_reg[6]  (.D(n_435), .G(n_428), .Q(n_16));
   DLH_X1 \A_in_reg[5]  (.D(n_434), .G(n_428), .Q(n_17));
   DLH_X1 \A_in_reg[4]  (.D(n_433), .G(n_428), .Q(n_18));
   DLH_X1 \A_in_reg[3]  (.D(n_432), .G(n_428), .Q(n_19));
   DLH_X1 \A_in_reg[2]  (.D(n_431), .G(n_428), .Q(n_20));
   DLH_X1 \A_in_reg[1]  (.D(n_430), .G(n_428), .Q(n_21));
   DLH_X1 \A_in_reg[0]  (.D(n_429), .G(n_428), .Q(n_22));
   DLH_X1 \B_in_reg[22]  (.D(n_427), .G(n_428), .Q(n_23));
   DLH_X1 \B_in_reg[21]  (.D(n_426), .G(n_428), .Q(n_24));
   DLH_X1 \B_in_reg[20]  (.D(n_425), .G(n_428), .Q(n_25));
   DLH_X1 \B_in_reg[19]  (.D(n_424), .G(n_428), .Q(n_26));
   DLH_X1 \B_in_reg[18]  (.D(n_423), .G(n_428), .Q(n_27));
   DLH_X1 \B_in_reg[17]  (.D(n_422), .G(n_428), .Q(n_28));
   DLH_X1 \B_in_reg[16]  (.D(n_421), .G(n_428), .Q(n_29));
   DLH_X1 \B_in_reg[15]  (.D(n_420), .G(n_428), .Q(n_30));
   DLH_X1 \B_in_reg[14]  (.D(n_419), .G(n_428), .Q(n_31));
   DLH_X1 \B_in_reg[13]  (.D(n_418), .G(n_428), .Q(n_32));
   DLH_X1 \B_in_reg[12]  (.D(n_417), .G(n_428), .Q(n_33));
   DLH_X1 \B_in_reg[11]  (.D(n_416), .G(n_428), .Q(n_34));
   DLH_X1 \B_in_reg[10]  (.D(n_415), .G(n_428), .Q(n_35));
   DLH_X1 \B_in_reg[9]  (.D(n_414), .G(n_428), .Q(n_36));
   DLH_X1 \B_in_reg[8]  (.D(n_413), .G(n_428), .Q(n_37));
   DLH_X1 \B_in_reg[7]  (.D(n_412), .G(n_428), .Q(n_38));
   DLH_X1 \B_in_reg[6]  (.D(n_411), .G(n_428), .Q(n_39));
   DLH_X1 \B_in_reg[5]  (.D(n_410), .G(n_428), .Q(n_40));
   DLH_X1 \B_in_reg[4]  (.D(n_409), .G(n_428), .Q(n_41));
   DLH_X1 \B_in_reg[3]  (.D(n_408), .G(n_428), .Q(n_42));
   DLH_X1 \B_in_reg[2]  (.D(n_407), .G(n_428), .Q(n_43));
   DLH_X1 \B_in_reg[1]  (.D(n_406), .G(n_428), .Q(n_44));
   DLH_X1 \B_in_reg[0]  (.D(n_405), .G(n_428), .Q(n_45));
   DLH_X1 \A_in_reg[23]  (.D(n_1_0__1), .G(n_428), .Q(n_46));
   OAI222_X1 i_0_0 (.A1(n_0_346), .A2(n_0_0), .B1(n_0_92), .B2(n_0_2), .C1(
      n_0_369), .C2(n_0_1), .ZN(n_47));
   OAI222_X1 i_0_1 (.A1(n_0_347), .A2(n_0_0), .B1(n_0_369), .B2(n_0_2), .C1(
      n_0_370), .C2(n_0_1), .ZN(n_48));
   OAI222_X1 i_0_2 (.A1(n_0_348), .A2(n_0_0), .B1(n_0_370), .B2(n_0_2), .C1(
      n_0_371), .C2(n_0_1), .ZN(n_49));
   OAI222_X1 i_0_3 (.A1(n_0_349), .A2(n_0_0), .B1(n_0_371), .B2(n_0_2), .C1(
      n_0_372), .C2(n_0_1), .ZN(n_50));
   OAI222_X1 i_0_4 (.A1(n_0_350), .A2(n_0_0), .B1(n_0_372), .B2(n_0_2), .C1(
      n_0_373), .C2(n_0_1), .ZN(n_51));
   OAI222_X1 i_0_5 (.A1(n_0_351), .A2(n_0_0), .B1(n_0_373), .B2(n_0_2), .C1(
      n_0_374), .C2(n_0_1), .ZN(n_52));
   OAI222_X1 i_0_6 (.A1(n_0_352), .A2(n_0_0), .B1(n_0_374), .B2(n_0_2), .C1(
      n_0_375), .C2(n_0_1), .ZN(n_53));
   OAI222_X1 i_0_7 (.A1(n_0_353), .A2(n_0_0), .B1(n_0_375), .B2(n_0_2), .C1(
      n_0_376), .C2(n_0_1), .ZN(n_54));
   OAI222_X1 i_0_8 (.A1(n_0_354), .A2(n_0_0), .B1(n_0_376), .B2(n_0_2), .C1(
      n_0_377), .C2(n_0_1), .ZN(n_55));
   OAI222_X1 i_0_9 (.A1(n_0_355), .A2(n_0_0), .B1(n_0_377), .B2(n_0_2), .C1(
      n_0_378), .C2(n_0_1), .ZN(n_56));
   OAI222_X1 i_0_10 (.A1(n_0_356), .A2(n_0_0), .B1(n_0_378), .B2(n_0_2), 
      .C1(n_0_379), .C2(n_0_1), .ZN(n_57));
   OAI222_X1 i_0_11 (.A1(n_0_357), .A2(n_0_0), .B1(n_0_379), .B2(n_0_2), 
      .C1(n_0_380), .C2(n_0_1), .ZN(n_58));
   OAI222_X1 i_0_12 (.A1(n_0_306), .A2(n_0_0), .B1(n_0_380), .B2(n_0_2), 
      .C1(n_0_305), .C2(n_0_1), .ZN(n_59));
   OAI222_X1 i_0_13 (.A1(n_0_359), .A2(n_0_0), .B1(n_0_305), .B2(n_0_2), 
      .C1(n_0_382), .C2(n_0_1), .ZN(n_60));
   OAI222_X1 i_0_14 (.A1(n_0_360), .A2(n_0_0), .B1(n_0_382), .B2(n_0_2), 
      .C1(n_0_383), .C2(n_0_1), .ZN(n_61));
   OAI222_X1 i_0_15 (.A1(n_0_361), .A2(n_0_0), .B1(n_0_383), .B2(n_0_2), 
      .C1(n_0_384), .C2(n_0_1), .ZN(n_62));
   OAI222_X1 i_0_16 (.A1(n_0_310), .A2(n_0_0), .B1(n_0_384), .B2(n_0_2), 
      .C1(n_0_385), .C2(n_0_1), .ZN(n_63));
   OAI222_X1 i_0_17 (.A1(n_0_363), .A2(n_0_0), .B1(n_0_385), .B2(n_0_2), 
      .C1(n_0_386), .C2(n_0_1), .ZN(n_64));
   OAI222_X1 i_0_18 (.A1(n_0_404), .A2(n_0_0), .B1(n_0_386), .B2(n_0_2), 
      .C1(n_0_403), .C2(n_0_1), .ZN(n_65));
   OAI222_X1 i_0_19 (.A1(n_0_365), .A2(n_0_0), .B1(n_0_403), .B2(n_0_2), 
      .C1(n_0_388), .C2(n_0_1), .ZN(n_66));
   OAI222_X1 i_0_20 (.A1(n_0_31), .A2(n_0_0), .B1(n_0_388), .B2(n_0_2), .C1(
      n_0_27), .C2(n_0_1), .ZN(n_67));
   OAI222_X1 i_0_21 (.A1(n_0_28), .A2(n_0_0), .B1(n_0_27), .B2(n_0_2), .C1(
      n_0_60), .C2(n_0_1), .ZN(n_68));
   NAND2_X1 i_0_22 (.A1(n_0_407), .A2(n_45), .ZN(n_0_0));
   OAI22_X1 i_0_23 (.A1(n_0_60), .A2(n_0_2), .B1(n_0_391), .B2(n_0_1), .ZN(n_69));
   NAND2_X1 i_0_24 (.A1(n_44), .A2(n_45), .ZN(n_0_1));
   OR2_X1 i_0_25 (.A1(n_0_407), .A2(n_45), .ZN(n_0_2));
   NOR2_X1 i_0_26 (.A1(n_0_407), .A2(n_0_391), .ZN(n_70));
   NOR2_X1 i_0_27 (.A1(n_0_28), .A2(n_0_344), .ZN(n_71));
   NOR2_X1 i_0_28 (.A1(n_0_28), .A2(n_0_95), .ZN(n_72));
   NOR2_X1 i_0_29 (.A1(n_0_28), .A2(n_0_346), .ZN(n_73));
   NOR2_X1 i_0_30 (.A1(n_0_28), .A2(n_0_347), .ZN(n_74));
   NOR2_X1 i_0_31 (.A1(n_0_28), .A2(n_0_348), .ZN(n_75));
   NOR2_X1 i_0_32 (.A1(n_0_28), .A2(n_0_349), .ZN(n_76));
   NOR2_X1 i_0_33 (.A1(n_0_28), .A2(n_0_350), .ZN(n_77));
   NOR2_X1 i_0_34 (.A1(n_0_28), .A2(n_0_351), .ZN(n_78));
   NOR2_X1 i_0_35 (.A1(n_0_28), .A2(n_0_352), .ZN(n_79));
   NOR2_X1 i_0_36 (.A1(n_0_28), .A2(n_0_353), .ZN(n_80));
   NOR2_X1 i_0_37 (.A1(n_0_28), .A2(n_0_354), .ZN(n_81));
   NOR2_X1 i_0_38 (.A1(n_0_28), .A2(n_0_355), .ZN(n_82));
   NOR2_X1 i_0_39 (.A1(n_0_28), .A2(n_0_356), .ZN(n_83));
   NOR2_X1 i_0_40 (.A1(n_0_28), .A2(n_0_357), .ZN(n_84));
   NOR2_X1 i_0_41 (.A1(n_0_28), .A2(n_0_306), .ZN(n_85));
   NOR2_X1 i_0_42 (.A1(n_0_28), .A2(n_0_359), .ZN(n_86));
   NOR2_X1 i_0_43 (.A1(n_0_28), .A2(n_0_360), .ZN(n_87));
   NOR2_X1 i_0_44 (.A1(n_0_28), .A2(n_0_361), .ZN(n_88));
   NOR2_X1 i_0_45 (.A1(n_0_28), .A2(n_0_310), .ZN(n_89));
   NOR2_X1 i_0_46 (.A1(n_0_28), .A2(n_0_363), .ZN(n_90));
   NOR2_X1 i_0_47 (.A1(n_0_28), .A2(n_0_404), .ZN(n_91));
   NOR2_X1 i_0_48 (.A1(n_0_28), .A2(n_0_365), .ZN(n_92));
   NOR2_X1 i_0_49 (.A1(n_0_28), .A2(n_0_31), .ZN(n_93));
   NOR2_X1 i_0_50 (.A1(n_0_344), .A2(n_0_61), .ZN(n_94));
   OAI221_X1 i_0_51 (.A(n_0_3), .B1(n_0_95), .B2(n_0_25), .C1(n_0_92), .C2(
      n_0_62), .ZN(n_95));
   OAI21_X1 i_0_52 (.A(n_22), .B1(n_0_29), .B2(n_0_26), .ZN(n_0_3));
   OAI221_X1 i_0_53 (.A(n_0_4), .B1(n_0_346), .B2(n_0_25), .C1(n_0_369), 
      .C2(n_0_62), .ZN(n_96));
   AOI22_X1 i_0_54 (.A1(n_21), .A2(n_0_26), .B1(A_imm_2s_complement[1]), 
      .B2(n_0_29), .ZN(n_0_4));
   OAI221_X1 i_0_55 (.A(n_0_5), .B1(n_0_347), .B2(n_0_25), .C1(n_0_370), 
      .C2(n_0_62), .ZN(n_97));
   AOI22_X1 i_0_56 (.A1(n_20), .A2(n_0_26), .B1(A_imm_2s_complement[2]), 
      .B2(n_0_29), .ZN(n_0_5));
   OAI221_X1 i_0_57 (.A(n_0_6), .B1(n_0_348), .B2(n_0_25), .C1(n_0_371), 
      .C2(n_0_62), .ZN(n_98));
   AOI22_X1 i_0_58 (.A1(n_19), .A2(n_0_26), .B1(A_imm_2s_complement[3]), 
      .B2(n_0_29), .ZN(n_0_6));
   OAI221_X1 i_0_59 (.A(n_0_7), .B1(n_0_349), .B2(n_0_25), .C1(n_0_372), 
      .C2(n_0_62), .ZN(n_99));
   AOI22_X1 i_0_60 (.A1(n_18), .A2(n_0_26), .B1(A_imm_2s_complement[4]), 
      .B2(n_0_29), .ZN(n_0_7));
   OAI221_X1 i_0_61 (.A(n_0_8), .B1(n_0_350), .B2(n_0_25), .C1(n_0_373), 
      .C2(n_0_62), .ZN(n_100));
   AOI22_X1 i_0_62 (.A1(n_17), .A2(n_0_26), .B1(A_imm_2s_complement[5]), 
      .B2(n_0_29), .ZN(n_0_8));
   OAI221_X1 i_0_63 (.A(n_0_9), .B1(n_0_351), .B2(n_0_25), .C1(n_0_374), 
      .C2(n_0_62), .ZN(n_101));
   AOI22_X1 i_0_64 (.A1(n_16), .A2(n_0_26), .B1(A_imm_2s_complement[6]), 
      .B2(n_0_29), .ZN(n_0_9));
   OAI221_X1 i_0_65 (.A(n_0_10), .B1(n_0_352), .B2(n_0_25), .C1(n_0_375), 
      .C2(n_0_62), .ZN(n_102));
   AOI22_X1 i_0_66 (.A1(n_15), .A2(n_0_26), .B1(A_imm_2s_complement[7]), 
      .B2(n_0_29), .ZN(n_0_10));
   OAI221_X1 i_0_67 (.A(n_0_11), .B1(n_0_353), .B2(n_0_25), .C1(n_0_376), 
      .C2(n_0_62), .ZN(n_103));
   AOI22_X1 i_0_68 (.A1(n_14), .A2(n_0_26), .B1(A_imm_2s_complement[8]), 
      .B2(n_0_29), .ZN(n_0_11));
   OAI221_X1 i_0_69 (.A(n_0_12), .B1(n_0_354), .B2(n_0_25), .C1(n_0_377), 
      .C2(n_0_62), .ZN(n_104));
   AOI22_X1 i_0_70 (.A1(n_13), .A2(n_0_26), .B1(A_imm_2s_complement[9]), 
      .B2(n_0_29), .ZN(n_0_12));
   OAI221_X1 i_0_71 (.A(n_0_13), .B1(n_0_355), .B2(n_0_25), .C1(n_0_378), 
      .C2(n_0_62), .ZN(n_105));
   AOI22_X1 i_0_72 (.A1(n_12), .A2(n_0_26), .B1(A_imm_2s_complement[10]), 
      .B2(n_0_29), .ZN(n_0_13));
   OAI221_X1 i_0_73 (.A(n_0_14), .B1(n_0_356), .B2(n_0_25), .C1(n_0_379), 
      .C2(n_0_62), .ZN(n_106));
   AOI22_X1 i_0_74 (.A1(n_11), .A2(n_0_26), .B1(A_imm_2s_complement[11]), 
      .B2(n_0_29), .ZN(n_0_14));
   OAI221_X1 i_0_75 (.A(n_0_15), .B1(n_0_357), .B2(n_0_25), .C1(n_0_380), 
      .C2(n_0_62), .ZN(n_107));
   AOI22_X1 i_0_76 (.A1(n_10), .A2(n_0_26), .B1(A_imm_2s_complement[12]), 
      .B2(n_0_29), .ZN(n_0_15));
   OAI221_X1 i_0_77 (.A(n_0_16), .B1(n_0_306), .B2(n_0_25), .C1(n_0_305), 
      .C2(n_0_62), .ZN(n_108));
   AOI22_X1 i_0_78 (.A1(n_9), .A2(n_0_26), .B1(A_imm_2s_complement[13]), 
      .B2(n_0_29), .ZN(n_0_16));
   OAI221_X1 i_0_79 (.A(n_0_17), .B1(n_0_359), .B2(n_0_25), .C1(n_0_382), 
      .C2(n_0_62), .ZN(n_109));
   AOI22_X1 i_0_80 (.A1(n_8), .A2(n_0_26), .B1(A_imm_2s_complement[14]), 
      .B2(n_0_29), .ZN(n_0_17));
   OAI221_X1 i_0_81 (.A(n_0_18), .B1(n_0_360), .B2(n_0_25), .C1(n_0_383), 
      .C2(n_0_62), .ZN(n_110));
   AOI22_X1 i_0_82 (.A1(n_7), .A2(n_0_26), .B1(A_imm_2s_complement[15]), 
      .B2(n_0_29), .ZN(n_0_18));
   OAI221_X1 i_0_83 (.A(n_0_19), .B1(n_0_361), .B2(n_0_25), .C1(n_0_384), 
      .C2(n_0_62), .ZN(n_111));
   AOI22_X1 i_0_84 (.A1(n_6), .A2(n_0_26), .B1(A_imm_2s_complement[16]), 
      .B2(n_0_29), .ZN(n_0_19));
   OAI221_X1 i_0_85 (.A(n_0_20), .B1(n_0_310), .B2(n_0_25), .C1(n_0_385), 
      .C2(n_0_62), .ZN(n_112));
   AOI22_X1 i_0_86 (.A1(n_5), .A2(n_0_26), .B1(A_imm_2s_complement[17]), 
      .B2(n_0_29), .ZN(n_0_20));
   OAI221_X1 i_0_87 (.A(n_0_21), .B1(n_0_363), .B2(n_0_25), .C1(n_0_386), 
      .C2(n_0_62), .ZN(n_113));
   AOI22_X1 i_0_88 (.A1(n_4), .A2(n_0_26), .B1(A_imm_2s_complement[18]), 
      .B2(n_0_29), .ZN(n_0_21));
   OAI221_X1 i_0_89 (.A(n_0_22), .B1(n_0_404), .B2(n_0_25), .C1(n_0_403), 
      .C2(n_0_62), .ZN(n_114));
   AOI22_X1 i_0_90 (.A1(n_3), .A2(n_0_26), .B1(A_imm_2s_complement[19]), 
      .B2(n_0_29), .ZN(n_0_22));
   OAI221_X1 i_0_91 (.A(n_0_23), .B1(n_0_365), .B2(n_0_25), .C1(n_0_388), 
      .C2(n_0_62), .ZN(n_115));
   AOI22_X1 i_0_92 (.A1(n_2), .A2(n_0_26), .B1(A_imm_2s_complement[20]), 
      .B2(n_0_29), .ZN(n_0_23));
   OAI221_X1 i_0_93 (.A(n_0_24), .B1(n_0_31), .B2(n_0_25), .C1(n_0_27), .C2(
      n_0_62), .ZN(n_116));
   AOI22_X1 i_0_94 (.A1(n_1), .A2(n_0_26), .B1(A_imm_2s_complement[21]), 
      .B2(n_0_29), .ZN(n_0_24));
   OR2_X1 i_0_95 (.A1(n_46), .A2(n_0_61), .ZN(n_0_25));
   INV_X1 i_0_96 (.A(n_0_59), .ZN(n_0_26));
   OAI22_X1 i_0_97 (.A1(n_0_60), .A2(n_0_30), .B1(n_0_32), .B2(n_0_61), .ZN(
      n_117));
   NOR2_X1 i_0_98 (.A1(n_0_57), .A2(n_0_32), .ZN(n_118));
   NAND2_X1 i_0_99 (.A1(A_imm_2s_complement[27]), .A2(n_46), .ZN(n_0_32));
   NOR2_X1 i_0_107 (.A1(n_0_344), .A2(n_0_93), .ZN(n_119));
   OAI221_X1 i_0_100 (.A(n_0_35), .B1(n_0_346), .B2(n_0_96), .C1(n_0_369), 
      .C2(n_0_94), .ZN(n_120));
   AOI22_X1 i_0_101 (.A1(A_imm_2s_complement[1]), .A2(n_0_91), .B1(n_21), 
      .B2(n_0_90), .ZN(n_0_35));
   OAI221_X1 i_0_112 (.A(n_0_36), .B1(n_0_347), .B2(n_0_96), .C1(n_0_370), 
      .C2(n_0_94), .ZN(n_121));
   AOI22_X1 i_0_113 (.A1(A_imm_2s_complement[2]), .A2(n_0_91), .B1(n_20), 
      .B2(n_0_90), .ZN(n_0_36));
   OAI221_X1 i_0_114 (.A(n_0_37), .B1(n_0_348), .B2(n_0_96), .C1(n_0_371), 
      .C2(n_0_94), .ZN(n_122));
   AOI22_X1 i_0_115 (.A1(A_imm_2s_complement[3]), .A2(n_0_91), .B1(n_19), 
      .B2(n_0_90), .ZN(n_0_37));
   OAI221_X1 i_0_116 (.A(n_0_38), .B1(n_0_349), .B2(n_0_96), .C1(n_0_372), 
      .C2(n_0_94), .ZN(n_123));
   AOI22_X1 i_0_117 (.A1(A_imm_2s_complement[4]), .A2(n_0_91), .B1(n_18), 
      .B2(n_0_90), .ZN(n_0_38));
   OAI221_X1 i_0_118 (.A(n_0_39), .B1(n_0_350), .B2(n_0_96), .C1(n_0_373), 
      .C2(n_0_94), .ZN(n_124));
   AOI22_X1 i_0_119 (.A1(A_imm_2s_complement[5]), .A2(n_0_91), .B1(n_17), 
      .B2(n_0_90), .ZN(n_0_39));
   OAI221_X1 i_0_120 (.A(n_0_40), .B1(n_0_351), .B2(n_0_96), .C1(n_0_374), 
      .C2(n_0_94), .ZN(n_125));
   AOI22_X1 i_0_121 (.A1(A_imm_2s_complement[6]), .A2(n_0_91), .B1(n_16), 
      .B2(n_0_90), .ZN(n_0_40));
   OAI221_X1 i_0_122 (.A(n_0_41), .B1(n_0_352), .B2(n_0_96), .C1(n_0_375), 
      .C2(n_0_94), .ZN(n_126));
   AOI22_X1 i_0_123 (.A1(A_imm_2s_complement[7]), .A2(n_0_91), .B1(n_15), 
      .B2(n_0_90), .ZN(n_0_41));
   OAI221_X1 i_0_124 (.A(n_0_42), .B1(n_0_353), .B2(n_0_96), .C1(n_0_376), 
      .C2(n_0_94), .ZN(n_127));
   AOI22_X1 i_0_125 (.A1(A_imm_2s_complement[8]), .A2(n_0_91), .B1(n_14), 
      .B2(n_0_90), .ZN(n_0_42));
   OAI221_X1 i_0_126 (.A(n_0_43), .B1(n_0_354), .B2(n_0_96), .C1(n_0_377), 
      .C2(n_0_94), .ZN(n_128));
   AOI22_X1 i_0_127 (.A1(A_imm_2s_complement[9]), .A2(n_0_91), .B1(n_13), 
      .B2(n_0_90), .ZN(n_0_43));
   OAI221_X1 i_0_128 (.A(n_0_44), .B1(n_0_355), .B2(n_0_96), .C1(n_0_378), 
      .C2(n_0_94), .ZN(n_129));
   AOI22_X1 i_0_129 (.A1(A_imm_2s_complement[10]), .A2(n_0_91), .B1(n_12), 
      .B2(n_0_90), .ZN(n_0_44));
   OAI221_X1 i_0_130 (.A(n_0_45), .B1(n_0_356), .B2(n_0_96), .C1(n_0_379), 
      .C2(n_0_94), .ZN(n_130));
   AOI22_X1 i_0_131 (.A1(A_imm_2s_complement[11]), .A2(n_0_91), .B1(n_11), 
      .B2(n_0_90), .ZN(n_0_45));
   OAI221_X1 i_0_132 (.A(n_0_46), .B1(n_0_357), .B2(n_0_96), .C1(n_0_380), 
      .C2(n_0_94), .ZN(n_131));
   AOI22_X1 i_0_133 (.A1(A_imm_2s_complement[12]), .A2(n_0_91), .B1(n_10), 
      .B2(n_0_90), .ZN(n_0_46));
   OAI221_X1 i_0_134 (.A(n_0_47), .B1(n_0_306), .B2(n_0_96), .C1(n_0_305), 
      .C2(n_0_94), .ZN(n_132));
   AOI22_X1 i_0_135 (.A1(A_imm_2s_complement[13]), .A2(n_0_91), .B1(n_9), 
      .B2(n_0_90), .ZN(n_0_47));
   OAI221_X1 i_0_136 (.A(n_0_48), .B1(n_0_359), .B2(n_0_96), .C1(n_0_382), 
      .C2(n_0_94), .ZN(n_133));
   AOI22_X1 i_0_137 (.A1(A_imm_2s_complement[14]), .A2(n_0_91), .B1(n_8), 
      .B2(n_0_90), .ZN(n_0_48));
   OAI221_X1 i_0_138 (.A(n_0_49), .B1(n_0_360), .B2(n_0_96), .C1(n_0_383), 
      .C2(n_0_94), .ZN(n_134));
   AOI22_X1 i_0_139 (.A1(A_imm_2s_complement[15]), .A2(n_0_91), .B1(n_7), 
      .B2(n_0_90), .ZN(n_0_49));
   OAI221_X1 i_0_140 (.A(n_0_50), .B1(n_0_361), .B2(n_0_96), .C1(n_0_384), 
      .C2(n_0_94), .ZN(n_135));
   AOI22_X1 i_0_141 (.A1(A_imm_2s_complement[16]), .A2(n_0_91), .B1(n_6), 
      .B2(n_0_90), .ZN(n_0_50));
   OAI221_X1 i_0_142 (.A(n_0_51), .B1(n_0_310), .B2(n_0_96), .C1(n_0_385), 
      .C2(n_0_94), .ZN(n_136));
   AOI22_X1 i_0_143 (.A1(A_imm_2s_complement[17]), .A2(n_0_91), .B1(n_5), 
      .B2(n_0_90), .ZN(n_0_51));
   OAI221_X1 i_0_144 (.A(n_0_52), .B1(n_0_363), .B2(n_0_96), .C1(n_0_386), 
      .C2(n_0_94), .ZN(n_137));
   AOI22_X1 i_0_145 (.A1(A_imm_2s_complement[18]), .A2(n_0_91), .B1(n_4), 
      .B2(n_0_90), .ZN(n_0_52));
   OAI221_X1 i_0_146 (.A(n_0_53), .B1(n_0_404), .B2(n_0_96), .C1(n_0_403), 
      .C2(n_0_94), .ZN(n_138));
   AOI22_X1 i_0_147 (.A1(A_imm_2s_complement[19]), .A2(n_0_91), .B1(n_3), 
      .B2(n_0_90), .ZN(n_0_53));
   OAI221_X1 i_0_148 (.A(n_0_54), .B1(n_0_365), .B2(n_0_96), .C1(n_0_388), 
      .C2(n_0_94), .ZN(n_139));
   AOI22_X1 i_0_149 (.A1(A_imm_2s_complement[20]), .A2(n_0_91), .B1(n_2), 
      .B2(n_0_90), .ZN(n_0_54));
   OAI221_X1 i_0_102 (.A(n_0_55), .B1(n_0_31), .B2(n_0_96), .C1(n_0_27), 
      .C2(n_0_94), .ZN(n_140));
   AOI22_X1 i_0_103 (.A1(A_imm_2s_complement[21]), .A2(n_0_91), .B1(n_1), 
      .B2(n_0_90), .ZN(n_0_55));
   OAI221_X1 i_0_152 (.A(n_0_56), .B1(n_0_28), .B2(n_0_96), .C1(n_0_60), 
      .C2(n_0_94), .ZN(n_141));
   AOI22_X1 i_0_153 (.A1(A_imm_2s_complement[22]), .A2(n_0_91), .B1(n_0), 
      .B2(n_0_90), .ZN(n_0_56));
   OAI222_X1 i_0_104 (.A1(n_0_28), .A2(n_0_88), .B1(n_0_60), .B2(n_0_58), 
      .C1(n_0_391), .C2(n_0_94), .ZN(n_142));
   INV_X1 i_0_105 (.A(n_0_91), .ZN(n_0_58));
   NOR3_X1 i_0_106 (.A1(n_0_33), .A2(n_0_391), .A3(n_0_65), .ZN(n_143));
   NOR2_X1 i_0_164 (.A1(n_0_344), .A2(n_0_127), .ZN(n_144));
   OAI221_X1 i_0_167 (.A(n_0_66), .B1(n_0_346), .B2(n_0_151), .C1(n_0_369), 
      .C2(n_0_150), .ZN(n_145));
   AOI22_X1 i_0_168 (.A1(A_imm_2s_complement[1]), .A2(n_0_126), .B1(n_21), 
      .B2(n_0_125), .ZN(n_0_66));
   OAI221_X1 i_0_169 (.A(n_0_67), .B1(n_0_347), .B2(n_0_151), .C1(n_0_370), 
      .C2(n_0_150), .ZN(n_146));
   AOI22_X1 i_0_170 (.A1(A_imm_2s_complement[2]), .A2(n_0_126), .B1(n_20), 
      .B2(n_0_125), .ZN(n_0_67));
   OAI221_X1 i_0_171 (.A(n_0_68), .B1(n_0_348), .B2(n_0_151), .C1(n_0_371), 
      .C2(n_0_150), .ZN(n_147));
   AOI22_X1 i_0_172 (.A1(A_imm_2s_complement[3]), .A2(n_0_126), .B1(n_19), 
      .B2(n_0_125), .ZN(n_0_68));
   OAI221_X1 i_0_173 (.A(n_0_69), .B1(n_0_349), .B2(n_0_151), .C1(n_0_372), 
      .C2(n_0_150), .ZN(n_148));
   AOI22_X1 i_0_174 (.A1(A_imm_2s_complement[4]), .A2(n_0_126), .B1(n_18), 
      .B2(n_0_125), .ZN(n_0_69));
   OAI221_X1 i_0_175 (.A(n_0_70), .B1(n_0_350), .B2(n_0_151), .C1(n_0_373), 
      .C2(n_0_150), .ZN(n_149));
   AOI22_X1 i_0_176 (.A1(A_imm_2s_complement[5]), .A2(n_0_126), .B1(n_17), 
      .B2(n_0_125), .ZN(n_0_70));
   OAI221_X1 i_0_177 (.A(n_0_71), .B1(n_0_351), .B2(n_0_151), .C1(n_0_374), 
      .C2(n_0_150), .ZN(n_150));
   AOI22_X1 i_0_178 (.A1(A_imm_2s_complement[6]), .A2(n_0_126), .B1(n_16), 
      .B2(n_0_125), .ZN(n_0_71));
   OAI221_X1 i_0_179 (.A(n_0_72), .B1(n_0_352), .B2(n_0_151), .C1(n_0_375), 
      .C2(n_0_150), .ZN(n_151));
   AOI22_X1 i_0_180 (.A1(A_imm_2s_complement[7]), .A2(n_0_126), .B1(n_15), 
      .B2(n_0_125), .ZN(n_0_72));
   OAI221_X1 i_0_181 (.A(n_0_73), .B1(n_0_353), .B2(n_0_151), .C1(n_0_376), 
      .C2(n_0_150), .ZN(n_152));
   AOI22_X1 i_0_182 (.A1(A_imm_2s_complement[8]), .A2(n_0_126), .B1(n_14), 
      .B2(n_0_125), .ZN(n_0_73));
   OAI221_X1 i_0_183 (.A(n_0_74), .B1(n_0_354), .B2(n_0_151), .C1(n_0_377), 
      .C2(n_0_150), .ZN(n_153));
   AOI22_X1 i_0_184 (.A1(A_imm_2s_complement[9]), .A2(n_0_126), .B1(n_13), 
      .B2(n_0_125), .ZN(n_0_74));
   OAI221_X1 i_0_185 (.A(n_0_75), .B1(n_0_355), .B2(n_0_151), .C1(n_0_378), 
      .C2(n_0_150), .ZN(n_154));
   AOI22_X1 i_0_186 (.A1(A_imm_2s_complement[10]), .A2(n_0_126), .B1(n_12), 
      .B2(n_0_125), .ZN(n_0_75));
   OAI221_X1 i_0_187 (.A(n_0_76), .B1(n_0_356), .B2(n_0_151), .C1(n_0_379), 
      .C2(n_0_150), .ZN(n_155));
   AOI22_X1 i_0_188 (.A1(A_imm_2s_complement[11]), .A2(n_0_126), .B1(n_11), 
      .B2(n_0_125), .ZN(n_0_76));
   OAI221_X1 i_0_189 (.A(n_0_77), .B1(n_0_357), .B2(n_0_151), .C1(n_0_380), 
      .C2(n_0_150), .ZN(n_156));
   AOI22_X1 i_0_190 (.A1(A_imm_2s_complement[12]), .A2(n_0_126), .B1(n_10), 
      .B2(n_0_125), .ZN(n_0_77));
   OAI221_X1 i_0_191 (.A(n_0_78), .B1(n_0_306), .B2(n_0_151), .C1(n_0_305), 
      .C2(n_0_150), .ZN(n_157));
   AOI22_X1 i_0_192 (.A1(A_imm_2s_complement[13]), .A2(n_0_126), .B1(n_9), 
      .B2(n_0_125), .ZN(n_0_78));
   OAI221_X1 i_0_193 (.A(n_0_79), .B1(n_0_359), .B2(n_0_151), .C1(n_0_382), 
      .C2(n_0_150), .ZN(n_158));
   AOI22_X1 i_0_194 (.A1(A_imm_2s_complement[14]), .A2(n_0_126), .B1(n_8), 
      .B2(n_0_125), .ZN(n_0_79));
   OAI221_X1 i_0_195 (.A(n_0_80), .B1(n_0_360), .B2(n_0_151), .C1(n_0_383), 
      .C2(n_0_150), .ZN(n_159));
   AOI22_X1 i_0_196 (.A1(A_imm_2s_complement[15]), .A2(n_0_126), .B1(n_7), 
      .B2(n_0_125), .ZN(n_0_80));
   OAI221_X1 i_0_197 (.A(n_0_81), .B1(n_0_361), .B2(n_0_151), .C1(n_0_384), 
      .C2(n_0_150), .ZN(n_160));
   AOI22_X1 i_0_198 (.A1(A_imm_2s_complement[16]), .A2(n_0_126), .B1(n_6), 
      .B2(n_0_125), .ZN(n_0_81));
   OAI221_X1 i_0_199 (.A(n_0_82), .B1(n_0_310), .B2(n_0_151), .C1(n_0_385), 
      .C2(n_0_150), .ZN(n_161));
   AOI22_X1 i_0_200 (.A1(A_imm_2s_complement[17]), .A2(n_0_126), .B1(n_5), 
      .B2(n_0_125), .ZN(n_0_82));
   OAI221_X1 i_0_201 (.A(n_0_83), .B1(n_0_363), .B2(n_0_151), .C1(n_0_386), 
      .C2(n_0_150), .ZN(n_162));
   AOI22_X1 i_0_202 (.A1(A_imm_2s_complement[18]), .A2(n_0_126), .B1(n_4), 
      .B2(n_0_125), .ZN(n_0_83));
   OAI221_X1 i_0_203 (.A(n_0_84), .B1(n_0_404), .B2(n_0_151), .C1(n_0_403), 
      .C2(n_0_150), .ZN(n_163));
   AOI22_X1 i_0_204 (.A1(A_imm_2s_complement[19]), .A2(n_0_126), .B1(n_3), 
      .B2(n_0_125), .ZN(n_0_84));
   OAI221_X1 i_0_205 (.A(n_0_85), .B1(n_0_365), .B2(n_0_151), .C1(n_0_388), 
      .C2(n_0_150), .ZN(n_164));
   AOI22_X1 i_0_206 (.A1(A_imm_2s_complement[20]), .A2(n_0_126), .B1(n_2), 
      .B2(n_0_125), .ZN(n_0_85));
   OAI221_X1 i_0_207 (.A(n_0_86), .B1(n_0_31), .B2(n_0_151), .C1(n_0_27), 
      .C2(n_0_150), .ZN(n_165));
   AOI22_X1 i_0_208 (.A1(A_imm_2s_complement[21]), .A2(n_0_126), .B1(n_1), 
      .B2(n_0_125), .ZN(n_0_86));
   OAI221_X1 i_0_209 (.A(n_0_87), .B1(n_0_28), .B2(n_0_151), .C1(n_0_60), 
      .C2(n_0_150), .ZN(n_166));
   AOI22_X1 i_0_210 (.A1(A_imm_2s_complement[22]), .A2(n_0_126), .B1(n_0), 
      .B2(n_0_125), .ZN(n_0_87));
   OAI222_X1 i_0_212 (.A1(n_0_28), .A2(n_0_124), .B1(n_0_60), .B2(n_0_89), 
      .C1(n_0_391), .C2(n_0_150), .ZN(n_167));
   INV_X1 i_0_213 (.A(n_0_126), .ZN(n_0_89));
   NOR3_X1 i_0_219 (.A1(n_0_63), .A2(n_0_391), .A3(n_0_123), .ZN(n_168));
   NOR2_X1 i_0_221 (.A1(n_0_344), .A2(n_0_182), .ZN(n_169));
   OAI221_X1 i_0_224 (.A(n_0_97), .B1(n_0_346), .B2(n_0_183), .C1(n_0_369), 
      .C2(n_0_185), .ZN(n_170));
   AOI22_X1 i_0_225 (.A1(n_21), .A2(n_0_181), .B1(A_imm_2s_complement[1]), 
      .B2(n_0_154), .ZN(n_0_97));
   OAI221_X1 i_0_226 (.A(n_0_98), .B1(n_0_347), .B2(n_0_183), .C1(n_0_370), 
      .C2(n_0_185), .ZN(n_171));
   AOI22_X1 i_0_227 (.A1(n_20), .A2(n_0_181), .B1(A_imm_2s_complement[2]), 
      .B2(n_0_154), .ZN(n_0_98));
   OAI221_X1 i_0_228 (.A(n_0_99), .B1(n_0_348), .B2(n_0_183), .C1(n_0_371), 
      .C2(n_0_185), .ZN(n_172));
   AOI22_X1 i_0_229 (.A1(n_19), .A2(n_0_181), .B1(A_imm_2s_complement[3]), 
      .B2(n_0_154), .ZN(n_0_99));
   OAI221_X1 i_0_230 (.A(n_0_100), .B1(n_0_349), .B2(n_0_183), .C1(n_0_372), 
      .C2(n_0_185), .ZN(n_173));
   AOI22_X1 i_0_231 (.A1(n_18), .A2(n_0_181), .B1(A_imm_2s_complement[4]), 
      .B2(n_0_154), .ZN(n_0_100));
   OAI221_X1 i_0_232 (.A(n_0_101), .B1(n_0_350), .B2(n_0_183), .C1(n_0_373), 
      .C2(n_0_185), .ZN(n_174));
   AOI22_X1 i_0_233 (.A1(n_17), .A2(n_0_181), .B1(A_imm_2s_complement[5]), 
      .B2(n_0_154), .ZN(n_0_101));
   OAI221_X1 i_0_234 (.A(n_0_102), .B1(n_0_351), .B2(n_0_183), .C1(n_0_374), 
      .C2(n_0_185), .ZN(n_175));
   AOI22_X1 i_0_235 (.A1(n_16), .A2(n_0_181), .B1(A_imm_2s_complement[6]), 
      .B2(n_0_154), .ZN(n_0_102));
   OAI221_X1 i_0_236 (.A(n_0_103), .B1(n_0_352), .B2(n_0_183), .C1(n_0_375), 
      .C2(n_0_185), .ZN(n_176));
   AOI22_X1 i_0_237 (.A1(n_15), .A2(n_0_181), .B1(A_imm_2s_complement[7]), 
      .B2(n_0_154), .ZN(n_0_103));
   OAI221_X1 i_0_238 (.A(n_0_104), .B1(n_0_353), .B2(n_0_183), .C1(n_0_376), 
      .C2(n_0_185), .ZN(n_177));
   AOI22_X1 i_0_239 (.A1(n_14), .A2(n_0_181), .B1(A_imm_2s_complement[8]), 
      .B2(n_0_154), .ZN(n_0_104));
   OAI221_X1 i_0_240 (.A(n_0_105), .B1(n_0_354), .B2(n_0_183), .C1(n_0_377), 
      .C2(n_0_185), .ZN(n_178));
   AOI22_X1 i_0_241 (.A1(n_13), .A2(n_0_181), .B1(A_imm_2s_complement[9]), 
      .B2(n_0_154), .ZN(n_0_105));
   OAI221_X1 i_0_242 (.A(n_0_106), .B1(n_0_355), .B2(n_0_183), .C1(n_0_378), 
      .C2(n_0_185), .ZN(n_179));
   AOI22_X1 i_0_243 (.A1(n_12), .A2(n_0_181), .B1(A_imm_2s_complement[10]), 
      .B2(n_0_154), .ZN(n_0_106));
   OAI221_X1 i_0_244 (.A(n_0_107), .B1(n_0_356), .B2(n_0_183), .C1(n_0_379), 
      .C2(n_0_185), .ZN(n_180));
   AOI22_X1 i_0_245 (.A1(n_11), .A2(n_0_181), .B1(A_imm_2s_complement[11]), 
      .B2(n_0_154), .ZN(n_0_107));
   OAI221_X1 i_0_246 (.A(n_0_108), .B1(n_0_357), .B2(n_0_183), .C1(n_0_380), 
      .C2(n_0_185), .ZN(n_181));
   AOI22_X1 i_0_247 (.A1(n_10), .A2(n_0_181), .B1(A_imm_2s_complement[12]), 
      .B2(n_0_154), .ZN(n_0_108));
   OAI221_X1 i_0_248 (.A(n_0_109), .B1(n_0_306), .B2(n_0_183), .C1(n_0_305), 
      .C2(n_0_185), .ZN(n_182));
   AOI22_X1 i_0_249 (.A1(n_9), .A2(n_0_181), .B1(A_imm_2s_complement[13]), 
      .B2(n_0_154), .ZN(n_0_109));
   OAI221_X1 i_0_250 (.A(n_0_110), .B1(n_0_359), .B2(n_0_183), .C1(n_0_382), 
      .C2(n_0_185), .ZN(n_183));
   AOI22_X1 i_0_251 (.A1(n_8), .A2(n_0_181), .B1(A_imm_2s_complement[14]), 
      .B2(n_0_154), .ZN(n_0_110));
   OAI221_X1 i_0_252 (.A(n_0_111), .B1(n_0_360), .B2(n_0_183), .C1(n_0_383), 
      .C2(n_0_185), .ZN(n_184));
   AOI22_X1 i_0_253 (.A1(n_7), .A2(n_0_181), .B1(A_imm_2s_complement[15]), 
      .B2(n_0_154), .ZN(n_0_111));
   OAI221_X1 i_0_254 (.A(n_0_112), .B1(n_0_361), .B2(n_0_183), .C1(n_0_384), 
      .C2(n_0_185), .ZN(n_185));
   AOI22_X1 i_0_255 (.A1(n_6), .A2(n_0_181), .B1(A_imm_2s_complement[16]), 
      .B2(n_0_154), .ZN(n_0_112));
   OAI221_X1 i_0_256 (.A(n_0_113), .B1(n_0_310), .B2(n_0_183), .C1(n_0_385), 
      .C2(n_0_185), .ZN(n_186));
   AOI22_X1 i_0_257 (.A1(n_5), .A2(n_0_181), .B1(A_imm_2s_complement[17]), 
      .B2(n_0_154), .ZN(n_0_113));
   OAI221_X1 i_0_258 (.A(n_0_114), .B1(n_0_363), .B2(n_0_183), .C1(n_0_386), 
      .C2(n_0_185), .ZN(n_187));
   AOI22_X1 i_0_259 (.A1(n_4), .A2(n_0_181), .B1(A_imm_2s_complement[18]), 
      .B2(n_0_154), .ZN(n_0_114));
   OAI221_X1 i_0_260 (.A(n_0_115), .B1(n_0_404), .B2(n_0_183), .C1(n_0_403), 
      .C2(n_0_185), .ZN(n_188));
   AOI22_X1 i_0_261 (.A1(n_3), .A2(n_0_181), .B1(A_imm_2s_complement[19]), 
      .B2(n_0_154), .ZN(n_0_115));
   OAI221_X1 i_0_262 (.A(n_0_116), .B1(n_0_365), .B2(n_0_183), .C1(n_0_388), 
      .C2(n_0_185), .ZN(n_189));
   AOI22_X1 i_0_263 (.A1(n_2), .A2(n_0_181), .B1(A_imm_2s_complement[20]), 
      .B2(n_0_154), .ZN(n_0_116));
   OAI221_X1 i_0_264 (.A(n_0_117), .B1(n_0_31), .B2(n_0_183), .C1(n_0_27), 
      .C2(n_0_185), .ZN(n_190));
   AOI22_X1 i_0_265 (.A1(n_1), .A2(n_0_181), .B1(A_imm_2s_complement[21]), 
      .B2(n_0_154), .ZN(n_0_117));
   OAI221_X1 i_0_266 (.A(n_0_118), .B1(n_0_28), .B2(n_0_183), .C1(n_0_60), 
      .C2(n_0_185), .ZN(n_191));
   AOI22_X1 i_0_267 (.A1(n_0), .A2(n_0_181), .B1(A_imm_2s_complement[22]), 
      .B2(n_0_154), .ZN(n_0_118));
   OAI222_X1 i_0_108 (.A1(n_0_60), .A2(n_0_122), .B1(n_0_28), .B2(n_0_158), 
      .C1(n_0_391), .C2(n_0_185), .ZN(n_192));
   INV_X1 i_0_109 (.A(n_0_154), .ZN(n_0_122));
   NOR3_X1 i_0_276 (.A1(n_0_120), .A2(n_0_391), .A3(n_0_157), .ZN(n_193));
   NOR2_X1 i_0_278 (.A1(n_0_344), .A2(n_0_213), .ZN(n_194));
   OAI221_X1 i_0_281 (.A(n_0_128), .B1(n_0_346), .B2(n_0_214), .C1(n_0_369), 
      .C2(n_0_216), .ZN(n_195));
   AOI22_X1 i_0_282 (.A1(n_21), .A2(n_0_212), .B1(A_imm_2s_complement[1]), 
      .B2(n_0_187), .ZN(n_0_128));
   OAI221_X1 i_0_283 (.A(n_0_129), .B1(n_0_347), .B2(n_0_214), .C1(n_0_370), 
      .C2(n_0_216), .ZN(n_196));
   AOI22_X1 i_0_284 (.A1(n_20), .A2(n_0_212), .B1(A_imm_2s_complement[2]), 
      .B2(n_0_187), .ZN(n_0_129));
   OAI221_X1 i_0_285 (.A(n_0_130), .B1(n_0_348), .B2(n_0_214), .C1(n_0_371), 
      .C2(n_0_216), .ZN(n_197));
   AOI22_X1 i_0_286 (.A1(n_19), .A2(n_0_212), .B1(A_imm_2s_complement[3]), 
      .B2(n_0_187), .ZN(n_0_130));
   OAI221_X1 i_0_287 (.A(n_0_131), .B1(n_0_349), .B2(n_0_214), .C1(n_0_372), 
      .C2(n_0_216), .ZN(n_198));
   AOI22_X1 i_0_288 (.A1(n_18), .A2(n_0_212), .B1(A_imm_2s_complement[4]), 
      .B2(n_0_187), .ZN(n_0_131));
   OAI221_X1 i_0_289 (.A(n_0_132), .B1(n_0_350), .B2(n_0_214), .C1(n_0_373), 
      .C2(n_0_216), .ZN(n_199));
   AOI22_X1 i_0_290 (.A1(n_17), .A2(n_0_212), .B1(A_imm_2s_complement[5]), 
      .B2(n_0_187), .ZN(n_0_132));
   OAI221_X1 i_0_291 (.A(n_0_133), .B1(n_0_351), .B2(n_0_214), .C1(n_0_374), 
      .C2(n_0_216), .ZN(n_200));
   AOI22_X1 i_0_292 (.A1(n_16), .A2(n_0_212), .B1(A_imm_2s_complement[6]), 
      .B2(n_0_187), .ZN(n_0_133));
   OAI221_X1 i_0_293 (.A(n_0_134), .B1(n_0_352), .B2(n_0_214), .C1(n_0_375), 
      .C2(n_0_216), .ZN(n_201));
   AOI22_X1 i_0_294 (.A1(n_15), .A2(n_0_212), .B1(A_imm_2s_complement[7]), 
      .B2(n_0_187), .ZN(n_0_134));
   OAI221_X1 i_0_295 (.A(n_0_135), .B1(n_0_353), .B2(n_0_214), .C1(n_0_376), 
      .C2(n_0_216), .ZN(n_202));
   AOI22_X1 i_0_296 (.A1(n_14), .A2(n_0_212), .B1(A_imm_2s_complement[8]), 
      .B2(n_0_187), .ZN(n_0_135));
   OAI221_X1 i_0_297 (.A(n_0_136), .B1(n_0_354), .B2(n_0_214), .C1(n_0_377), 
      .C2(n_0_216), .ZN(n_203));
   AOI22_X1 i_0_298 (.A1(n_13), .A2(n_0_212), .B1(A_imm_2s_complement[9]), 
      .B2(n_0_187), .ZN(n_0_136));
   OAI221_X1 i_0_299 (.A(n_0_137), .B1(n_0_355), .B2(n_0_214), .C1(n_0_378), 
      .C2(n_0_216), .ZN(n_204));
   AOI22_X1 i_0_300 (.A1(n_12), .A2(n_0_212), .B1(A_imm_2s_complement[10]), 
      .B2(n_0_187), .ZN(n_0_137));
   OAI221_X1 i_0_301 (.A(n_0_138), .B1(n_0_356), .B2(n_0_214), .C1(n_0_379), 
      .C2(n_0_216), .ZN(n_205));
   AOI22_X1 i_0_302 (.A1(n_11), .A2(n_0_212), .B1(A_imm_2s_complement[11]), 
      .B2(n_0_187), .ZN(n_0_138));
   OAI221_X1 i_0_303 (.A(n_0_139), .B1(n_0_357), .B2(n_0_214), .C1(n_0_380), 
      .C2(n_0_216), .ZN(n_206));
   AOI22_X1 i_0_304 (.A1(n_10), .A2(n_0_212), .B1(A_imm_2s_complement[12]), 
      .B2(n_0_187), .ZN(n_0_139));
   OAI221_X1 i_0_305 (.A(n_0_140), .B1(n_0_306), .B2(n_0_214), .C1(n_0_305), 
      .C2(n_0_216), .ZN(n_207));
   AOI22_X1 i_0_306 (.A1(n_9), .A2(n_0_212), .B1(A_imm_2s_complement[13]), 
      .B2(n_0_187), .ZN(n_0_140));
   OAI221_X1 i_0_307 (.A(n_0_141), .B1(n_0_359), .B2(n_0_214), .C1(n_0_382), 
      .C2(n_0_216), .ZN(n_208));
   AOI22_X1 i_0_308 (.A1(n_8), .A2(n_0_212), .B1(A_imm_2s_complement[14]), 
      .B2(n_0_187), .ZN(n_0_141));
   OAI221_X1 i_0_309 (.A(n_0_142), .B1(n_0_360), .B2(n_0_214), .C1(n_0_383), 
      .C2(n_0_216), .ZN(n_209));
   AOI22_X1 i_0_310 (.A1(n_7), .A2(n_0_212), .B1(A_imm_2s_complement[15]), 
      .B2(n_0_187), .ZN(n_0_142));
   OAI221_X1 i_0_311 (.A(n_0_143), .B1(n_0_361), .B2(n_0_214), .C1(n_0_384), 
      .C2(n_0_216), .ZN(n_210));
   AOI22_X1 i_0_312 (.A1(n_6), .A2(n_0_212), .B1(A_imm_2s_complement[16]), 
      .B2(n_0_187), .ZN(n_0_143));
   OAI221_X1 i_0_313 (.A(n_0_144), .B1(n_0_310), .B2(n_0_214), .C1(n_0_385), 
      .C2(n_0_216), .ZN(n_211));
   AOI22_X1 i_0_314 (.A1(n_5), .A2(n_0_212), .B1(A_imm_2s_complement[17]), 
      .B2(n_0_187), .ZN(n_0_144));
   OAI221_X1 i_0_315 (.A(n_0_145), .B1(n_0_363), .B2(n_0_214), .C1(n_0_386), 
      .C2(n_0_216), .ZN(n_212));
   AOI22_X1 i_0_316 (.A1(n_4), .A2(n_0_212), .B1(A_imm_2s_complement[18]), 
      .B2(n_0_187), .ZN(n_0_145));
   OAI221_X1 i_0_317 (.A(n_0_146), .B1(n_0_404), .B2(n_0_214), .C1(n_0_403), 
      .C2(n_0_216), .ZN(n_213));
   AOI22_X1 i_0_318 (.A1(n_3), .A2(n_0_212), .B1(A_imm_2s_complement[19]), 
      .B2(n_0_187), .ZN(n_0_146));
   OAI221_X1 i_0_319 (.A(n_0_147), .B1(n_0_365), .B2(n_0_214), .C1(n_0_388), 
      .C2(n_0_216), .ZN(n_214));
   AOI22_X1 i_0_320 (.A1(n_2), .A2(n_0_212), .B1(A_imm_2s_complement[20]), 
      .B2(n_0_187), .ZN(n_0_147));
   OAI221_X1 i_0_321 (.A(n_0_148), .B1(n_0_31), .B2(n_0_214), .C1(n_0_27), 
      .C2(n_0_216), .ZN(n_215));
   AOI22_X1 i_0_322 (.A1(n_1), .A2(n_0_212), .B1(A_imm_2s_complement[21]), 
      .B2(n_0_187), .ZN(n_0_148));
   OAI221_X1 i_0_323 (.A(n_0_149), .B1(n_0_28), .B2(n_0_214), .C1(n_0_60), 
      .C2(n_0_216), .ZN(n_216));
   AOI22_X1 i_0_324 (.A1(n_0), .A2(n_0_212), .B1(A_imm_2s_complement[22]), 
      .B2(n_0_187), .ZN(n_0_149));
   OAI222_X1 i_0_326 (.A1(n_0_60), .A2(n_0_153), .B1(n_0_28), .B2(n_0_206), 
      .C1(n_0_391), .C2(n_0_216), .ZN(n_217));
   INV_X1 i_0_329 (.A(n_0_187), .ZN(n_0_153));
   NOR3_X1 i_0_333 (.A1(n_0_155), .A2(n_0_391), .A3(n_0_202), .ZN(n_218));
   NOR2_X1 i_0_335 (.A1(n_0_344), .A2(n_0_247), .ZN(n_219));
   OAI221_X1 i_0_338 (.A(n_0_159), .B1(n_0_346), .B2(n_0_248), .C1(n_0_369), 
      .C2(n_0_249), .ZN(n_220));
   AOI22_X1 i_0_339 (.A1(n_21), .A2(n_0_245), .B1(A_imm_2s_complement[1]), 
      .B2(n_0_218), .ZN(n_0_159));
   OAI221_X1 i_0_340 (.A(n_0_160), .B1(n_0_347), .B2(n_0_248), .C1(n_0_370), 
      .C2(n_0_249), .ZN(n_221));
   AOI22_X1 i_0_341 (.A1(n_20), .A2(n_0_245), .B1(A_imm_2s_complement[2]), 
      .B2(n_0_218), .ZN(n_0_160));
   OAI221_X1 i_0_342 (.A(n_0_161), .B1(n_0_348), .B2(n_0_248), .C1(n_0_371), 
      .C2(n_0_249), .ZN(n_222));
   AOI22_X1 i_0_343 (.A1(n_19), .A2(n_0_245), .B1(A_imm_2s_complement[3]), 
      .B2(n_0_218), .ZN(n_0_161));
   OAI221_X1 i_0_344 (.A(n_0_162), .B1(n_0_349), .B2(n_0_248), .C1(n_0_372), 
      .C2(n_0_249), .ZN(n_223));
   AOI22_X1 i_0_345 (.A1(n_18), .A2(n_0_245), .B1(A_imm_2s_complement[4]), 
      .B2(n_0_218), .ZN(n_0_162));
   OAI221_X1 i_0_346 (.A(n_0_163), .B1(n_0_350), .B2(n_0_248), .C1(n_0_373), 
      .C2(n_0_249), .ZN(n_224));
   AOI22_X1 i_0_347 (.A1(n_17), .A2(n_0_245), .B1(A_imm_2s_complement[5]), 
      .B2(n_0_218), .ZN(n_0_163));
   OAI221_X1 i_0_348 (.A(n_0_164), .B1(n_0_351), .B2(n_0_248), .C1(n_0_374), 
      .C2(n_0_249), .ZN(n_225));
   AOI22_X1 i_0_349 (.A1(n_16), .A2(n_0_245), .B1(A_imm_2s_complement[6]), 
      .B2(n_0_218), .ZN(n_0_164));
   OAI221_X1 i_0_350 (.A(n_0_165), .B1(n_0_352), .B2(n_0_248), .C1(n_0_375), 
      .C2(n_0_249), .ZN(n_226));
   AOI22_X1 i_0_351 (.A1(n_15), .A2(n_0_245), .B1(A_imm_2s_complement[7]), 
      .B2(n_0_218), .ZN(n_0_165));
   OAI221_X1 i_0_352 (.A(n_0_166), .B1(n_0_353), .B2(n_0_248), .C1(n_0_376), 
      .C2(n_0_249), .ZN(n_227));
   AOI22_X1 i_0_353 (.A1(n_14), .A2(n_0_245), .B1(A_imm_2s_complement[8]), 
      .B2(n_0_218), .ZN(n_0_166));
   OAI221_X1 i_0_354 (.A(n_0_167), .B1(n_0_354), .B2(n_0_248), .C1(n_0_377), 
      .C2(n_0_249), .ZN(n_228));
   AOI22_X1 i_0_355 (.A1(n_13), .A2(n_0_245), .B1(A_imm_2s_complement[9]), 
      .B2(n_0_218), .ZN(n_0_167));
   OAI221_X1 i_0_356 (.A(n_0_168), .B1(n_0_355), .B2(n_0_248), .C1(n_0_378), 
      .C2(n_0_249), .ZN(n_229));
   AOI22_X1 i_0_357 (.A1(n_12), .A2(n_0_245), .B1(A_imm_2s_complement[10]), 
      .B2(n_0_218), .ZN(n_0_168));
   OAI221_X1 i_0_358 (.A(n_0_169), .B1(n_0_356), .B2(n_0_248), .C1(n_0_379), 
      .C2(n_0_249), .ZN(n_230));
   AOI22_X1 i_0_359 (.A1(n_11), .A2(n_0_245), .B1(A_imm_2s_complement[11]), 
      .B2(n_0_218), .ZN(n_0_169));
   OAI221_X1 i_0_360 (.A(n_0_170), .B1(n_0_357), .B2(n_0_248), .C1(n_0_380), 
      .C2(n_0_249), .ZN(n_231));
   AOI22_X1 i_0_361 (.A1(n_10), .A2(n_0_245), .B1(A_imm_2s_complement[12]), 
      .B2(n_0_218), .ZN(n_0_170));
   OAI221_X1 i_0_362 (.A(n_0_171), .B1(n_0_306), .B2(n_0_248), .C1(n_0_305), 
      .C2(n_0_249), .ZN(n_232));
   AOI22_X1 i_0_363 (.A1(n_9), .A2(n_0_245), .B1(A_imm_2s_complement[13]), 
      .B2(n_0_218), .ZN(n_0_171));
   OAI221_X1 i_0_364 (.A(n_0_172), .B1(n_0_359), .B2(n_0_248), .C1(n_0_382), 
      .C2(n_0_249), .ZN(n_233));
   AOI22_X1 i_0_365 (.A1(n_8), .A2(n_0_245), .B1(A_imm_2s_complement[14]), 
      .B2(n_0_218), .ZN(n_0_172));
   OAI221_X1 i_0_366 (.A(n_0_173), .B1(n_0_360), .B2(n_0_248), .C1(n_0_383), 
      .C2(n_0_249), .ZN(n_234));
   AOI22_X1 i_0_367 (.A1(n_7), .A2(n_0_245), .B1(A_imm_2s_complement[15]), 
      .B2(n_0_218), .ZN(n_0_173));
   OAI221_X1 i_0_368 (.A(n_0_174), .B1(n_0_361), .B2(n_0_248), .C1(n_0_384), 
      .C2(n_0_249), .ZN(n_235));
   AOI22_X1 i_0_369 (.A1(n_6), .A2(n_0_245), .B1(A_imm_2s_complement[16]), 
      .B2(n_0_218), .ZN(n_0_174));
   OAI221_X1 i_0_370 (.A(n_0_175), .B1(n_0_310), .B2(n_0_248), .C1(n_0_385), 
      .C2(n_0_249), .ZN(n_236));
   AOI22_X1 i_0_371 (.A1(n_5), .A2(n_0_245), .B1(A_imm_2s_complement[17]), 
      .B2(n_0_218), .ZN(n_0_175));
   OAI221_X1 i_0_372 (.A(n_0_176), .B1(n_0_363), .B2(n_0_248), .C1(n_0_386), 
      .C2(n_0_249), .ZN(n_237));
   AOI22_X1 i_0_373 (.A1(n_4), .A2(n_0_245), .B1(A_imm_2s_complement[18]), 
      .B2(n_0_218), .ZN(n_0_176));
   OAI221_X1 i_0_374 (.A(n_0_177), .B1(n_0_404), .B2(n_0_248), .C1(n_0_403), 
      .C2(n_0_249), .ZN(n_238));
   AOI22_X1 i_0_375 (.A1(n_3), .A2(n_0_245), .B1(A_imm_2s_complement[19]), 
      .B2(n_0_218), .ZN(n_0_177));
   OAI221_X1 i_0_376 (.A(n_0_178), .B1(n_0_365), .B2(n_0_248), .C1(n_0_388), 
      .C2(n_0_249), .ZN(n_239));
   AOI22_X1 i_0_377 (.A1(n_2), .A2(n_0_245), .B1(A_imm_2s_complement[20]), 
      .B2(n_0_218), .ZN(n_0_178));
   OAI221_X1 i_0_378 (.A(n_0_179), .B1(n_0_31), .B2(n_0_248), .C1(n_0_27), 
      .C2(n_0_249), .ZN(n_240));
   AOI22_X1 i_0_379 (.A1(n_1), .A2(n_0_245), .B1(A_imm_2s_complement[21]), 
      .B2(n_0_218), .ZN(n_0_179));
   OAI221_X1 i_0_380 (.A(n_0_180), .B1(n_0_28), .B2(n_0_248), .C1(n_0_60), 
      .C2(n_0_249), .ZN(n_241));
   AOI22_X1 i_0_381 (.A1(n_0), .A2(n_0_245), .B1(A_imm_2s_complement[22]), 
      .B2(n_0_218), .ZN(n_0_180));
   OAI222_X1 i_0_383 (.A1(n_0_60), .A2(n_0_184), .B1(n_0_28), .B2(n_0_244), 
      .C1(n_0_391), .C2(n_0_249), .ZN(n_242));
   INV_X1 i_0_386 (.A(n_0_218), .ZN(n_0_184));
   NOR3_X1 i_0_390 (.A1(n_0_188), .A2(n_0_391), .A3(n_0_243), .ZN(n_243));
   NOR2_X1 i_0_392 (.A1(n_0_344), .A2(n_0_279), .ZN(n_244));
   OAI221_X1 i_0_395 (.A(n_0_190), .B1(n_0_346), .B2(n_0_282), .C1(n_0_369), 
      .C2(n_0_281), .ZN(n_245));
   AOI22_X1 i_0_396 (.A1(n_21), .A2(n_0_278), .B1(A_imm_2s_complement[1]), 
      .B2(n_0_251), .ZN(n_0_190));
   OAI221_X1 i_0_397 (.A(n_0_191), .B1(n_0_347), .B2(n_0_282), .C1(n_0_370), 
      .C2(n_0_281), .ZN(n_246));
   AOI22_X1 i_0_398 (.A1(n_20), .A2(n_0_278), .B1(A_imm_2s_complement[2]), 
      .B2(n_0_251), .ZN(n_0_191));
   OAI221_X1 i_0_399 (.A(n_0_192), .B1(n_0_348), .B2(n_0_282), .C1(n_0_371), 
      .C2(n_0_281), .ZN(n_247));
   AOI22_X1 i_0_400 (.A1(n_19), .A2(n_0_278), .B1(A_imm_2s_complement[3]), 
      .B2(n_0_251), .ZN(n_0_192));
   OAI221_X1 i_0_401 (.A(n_0_193), .B1(n_0_349), .B2(n_0_282), .C1(n_0_372), 
      .C2(n_0_281), .ZN(n_248));
   AOI22_X1 i_0_402 (.A1(n_18), .A2(n_0_278), .B1(A_imm_2s_complement[4]), 
      .B2(n_0_251), .ZN(n_0_193));
   OAI221_X1 i_0_403 (.A(n_0_194), .B1(n_0_350), .B2(n_0_282), .C1(n_0_373), 
      .C2(n_0_281), .ZN(n_249));
   AOI22_X1 i_0_404 (.A1(n_17), .A2(n_0_278), .B1(A_imm_2s_complement[5]), 
      .B2(n_0_251), .ZN(n_0_194));
   OAI221_X1 i_0_405 (.A(n_0_195), .B1(n_0_351), .B2(n_0_282), .C1(n_0_374), 
      .C2(n_0_281), .ZN(n_250));
   AOI22_X1 i_0_406 (.A1(n_16), .A2(n_0_278), .B1(A_imm_2s_complement[6]), 
      .B2(n_0_251), .ZN(n_0_195));
   OAI221_X1 i_0_407 (.A(n_0_196), .B1(n_0_352), .B2(n_0_282), .C1(n_0_375), 
      .C2(n_0_281), .ZN(n_251));
   AOI22_X1 i_0_408 (.A1(n_15), .A2(n_0_278), .B1(A_imm_2s_complement[7]), 
      .B2(n_0_251), .ZN(n_0_196));
   OAI221_X1 i_0_409 (.A(n_0_197), .B1(n_0_353), .B2(n_0_282), .C1(n_0_376), 
      .C2(n_0_281), .ZN(n_252));
   AOI22_X1 i_0_410 (.A1(n_14), .A2(n_0_278), .B1(A_imm_2s_complement[8]), 
      .B2(n_0_251), .ZN(n_0_197));
   OAI221_X1 i_0_411 (.A(n_0_198), .B1(n_0_354), .B2(n_0_282), .C1(n_0_377), 
      .C2(n_0_281), .ZN(n_253));
   AOI22_X1 i_0_412 (.A1(n_13), .A2(n_0_278), .B1(A_imm_2s_complement[9]), 
      .B2(n_0_251), .ZN(n_0_198));
   OAI221_X1 i_0_413 (.A(n_0_199), .B1(n_0_355), .B2(n_0_282), .C1(n_0_378), 
      .C2(n_0_281), .ZN(n_254));
   AOI22_X1 i_0_414 (.A1(n_12), .A2(n_0_278), .B1(A_imm_2s_complement[10]), 
      .B2(n_0_251), .ZN(n_0_199));
   OAI221_X1 i_0_415 (.A(n_0_200), .B1(n_0_356), .B2(n_0_282), .C1(n_0_379), 
      .C2(n_0_281), .ZN(n_255));
   AOI22_X1 i_0_416 (.A1(n_11), .A2(n_0_278), .B1(A_imm_2s_complement[11]), 
      .B2(n_0_251), .ZN(n_0_200));
   OAI221_X1 i_0_417 (.A(n_0_201), .B1(n_0_357), .B2(n_0_282), .C1(n_0_380), 
      .C2(n_0_281), .ZN(n_256));
   AOI22_X1 i_0_418 (.A1(n_10), .A2(n_0_278), .B1(A_imm_2s_complement[12]), 
      .B2(n_0_251), .ZN(n_0_201));
   OAI221_X1 i_0_421 (.A(n_0_203), .B1(n_0_359), .B2(n_0_282), .C1(n_0_382), 
      .C2(n_0_281), .ZN(n_257));
   AOI22_X1 i_0_422 (.A1(n_8), .A2(n_0_278), .B1(A_imm_2s_complement[14]), 
      .B2(n_0_251), .ZN(n_0_203));
   OAI221_X1 i_0_423 (.A(n_0_204), .B1(n_0_360), .B2(n_0_282), .C1(n_0_383), 
      .C2(n_0_281), .ZN(n_258));
   AOI22_X1 i_0_424 (.A1(n_7), .A2(n_0_278), .B1(A_imm_2s_complement[15]), 
      .B2(n_0_251), .ZN(n_0_204));
   OAI221_X1 i_0_425 (.A(n_0_205), .B1(n_0_361), .B2(n_0_282), .C1(n_0_384), 
      .C2(n_0_281), .ZN(n_259));
   AOI22_X1 i_0_426 (.A1(n_6), .A2(n_0_278), .B1(A_imm_2s_complement[16]), 
      .B2(n_0_251), .ZN(n_0_205));
   OAI221_X1 i_0_429 (.A(n_0_207), .B1(n_0_363), .B2(n_0_282), .C1(n_0_386), 
      .C2(n_0_281), .ZN(n_260));
   AOI22_X1 i_0_430 (.A1(n_4), .A2(n_0_278), .B1(A_imm_2s_complement[18]), 
      .B2(n_0_251), .ZN(n_0_207));
   OAI221_X1 i_0_431 (.A(n_0_208), .B1(n_0_404), .B2(n_0_282), .C1(n_0_403), 
      .C2(n_0_281), .ZN(n_261));
   AOI22_X1 i_0_432 (.A1(n_3), .A2(n_0_278), .B1(A_imm_2s_complement[19]), 
      .B2(n_0_251), .ZN(n_0_208));
   OAI221_X1 i_0_433 (.A(n_0_209), .B1(n_0_365), .B2(n_0_282), .C1(n_0_388), 
      .C2(n_0_281), .ZN(n_262));
   AOI22_X1 i_0_434 (.A1(n_2), .A2(n_0_278), .B1(A_imm_2s_complement[20]), 
      .B2(n_0_251), .ZN(n_0_209));
   OAI221_X1 i_0_435 (.A(n_0_210), .B1(n_0_31), .B2(n_0_282), .C1(n_0_27), 
      .C2(n_0_281), .ZN(n_263));
   AOI22_X1 i_0_436 (.A1(n_1), .A2(n_0_278), .B1(A_imm_2s_complement[21]), 
      .B2(n_0_251), .ZN(n_0_210));
   OAI221_X1 i_0_437 (.A(n_0_211), .B1(n_0_28), .B2(n_0_282), .C1(n_0_60), 
      .C2(n_0_281), .ZN(n_264));
   AOI22_X1 i_0_438 (.A1(n_0), .A2(n_0_278), .B1(A_imm_2s_complement[22]), 
      .B2(n_0_251), .ZN(n_0_211));
   OAI222_X1 i_0_440 (.A1(n_0_60), .A2(n_0_215), .B1(n_0_28), .B2(n_0_276), 
      .C1(n_0_391), .C2(n_0_281), .ZN(n_265));
   INV_X1 i_0_443 (.A(n_0_251), .ZN(n_0_215));
   NOR3_X1 i_0_447 (.A1(n_0_219), .A2(n_0_391), .A3(n_0_275), .ZN(n_266));
   NOR2_X1 i_0_449 (.A1(n_0_344), .A2(n_0_337), .ZN(n_267));
   OAI221_X1 i_0_452 (.A(n_0_221), .B1(n_0_346), .B2(n_0_338), .C1(n_0_369), 
      .C2(n_0_340), .ZN(n_268));
   AOI22_X1 i_0_453 (.A1(n_21), .A2(n_0_336), .B1(A_imm_2s_complement[1]), 
      .B2(n_0_311), .ZN(n_0_221));
   OAI221_X1 i_0_454 (.A(n_0_222), .B1(n_0_347), .B2(n_0_338), .C1(n_0_370), 
      .C2(n_0_340), .ZN(n_269));
   AOI22_X1 i_0_455 (.A1(n_20), .A2(n_0_336), .B1(A_imm_2s_complement[2]), 
      .B2(n_0_311), .ZN(n_0_222));
   OAI221_X1 i_0_456 (.A(n_0_223), .B1(n_0_348), .B2(n_0_338), .C1(n_0_371), 
      .C2(n_0_340), .ZN(n_270));
   AOI22_X1 i_0_457 (.A1(n_19), .A2(n_0_336), .B1(A_imm_2s_complement[3]), 
      .B2(n_0_311), .ZN(n_0_223));
   OAI221_X1 i_0_458 (.A(n_0_224), .B1(n_0_349), .B2(n_0_338), .C1(n_0_372), 
      .C2(n_0_340), .ZN(n_271));
   AOI22_X1 i_0_459 (.A1(n_18), .A2(n_0_336), .B1(A_imm_2s_complement[4]), 
      .B2(n_0_311), .ZN(n_0_224));
   OAI221_X1 i_0_460 (.A(n_0_225), .B1(n_0_350), .B2(n_0_338), .C1(n_0_373), 
      .C2(n_0_340), .ZN(n_272));
   AOI22_X1 i_0_461 (.A1(n_17), .A2(n_0_336), .B1(A_imm_2s_complement[5]), 
      .B2(n_0_311), .ZN(n_0_225));
   OAI221_X1 i_0_462 (.A(n_0_226), .B1(n_0_351), .B2(n_0_338), .C1(n_0_374), 
      .C2(n_0_340), .ZN(n_273));
   AOI22_X1 i_0_463 (.A1(n_16), .A2(n_0_336), .B1(A_imm_2s_complement[6]), 
      .B2(n_0_311), .ZN(n_0_226));
   OAI221_X1 i_0_464 (.A(n_0_227), .B1(n_0_352), .B2(n_0_338), .C1(n_0_375), 
      .C2(n_0_340), .ZN(n_274));
   AOI22_X1 i_0_465 (.A1(n_15), .A2(n_0_336), .B1(A_imm_2s_complement[7]), 
      .B2(n_0_311), .ZN(n_0_227));
   OAI221_X1 i_0_466 (.A(n_0_228), .B1(n_0_353), .B2(n_0_338), .C1(n_0_376), 
      .C2(n_0_340), .ZN(n_275));
   AOI22_X1 i_0_467 (.A1(n_14), .A2(n_0_336), .B1(A_imm_2s_complement[8]), 
      .B2(n_0_311), .ZN(n_0_228));
   OAI221_X1 i_0_468 (.A(n_0_229), .B1(n_0_354), .B2(n_0_338), .C1(n_0_377), 
      .C2(n_0_340), .ZN(n_276));
   AOI22_X1 i_0_469 (.A1(n_13), .A2(n_0_336), .B1(A_imm_2s_complement[9]), 
      .B2(n_0_311), .ZN(n_0_229));
   OAI221_X1 i_0_470 (.A(n_0_230), .B1(n_0_355), .B2(n_0_338), .C1(n_0_378), 
      .C2(n_0_340), .ZN(n_277));
   AOI22_X1 i_0_471 (.A1(n_12), .A2(n_0_336), .B1(A_imm_2s_complement[10]), 
      .B2(n_0_311), .ZN(n_0_230));
   OAI221_X1 i_0_472 (.A(n_0_231), .B1(n_0_356), .B2(n_0_338), .C1(n_0_379), 
      .C2(n_0_340), .ZN(n_278));
   AOI22_X1 i_0_473 (.A1(n_11), .A2(n_0_336), .B1(A_imm_2s_complement[11]), 
      .B2(n_0_311), .ZN(n_0_231));
   OAI221_X1 i_0_474 (.A(n_0_232), .B1(n_0_357), .B2(n_0_338), .C1(n_0_380), 
      .C2(n_0_340), .ZN(n_279));
   AOI22_X1 i_0_475 (.A1(n_10), .A2(n_0_336), .B1(A_imm_2s_complement[12]), 
      .B2(n_0_311), .ZN(n_0_232));
   OAI221_X1 i_0_476 (.A(n_0_233), .B1(n_0_306), .B2(n_0_338), .C1(n_0_305), 
      .C2(n_0_340), .ZN(n_280));
   AOI22_X1 i_0_477 (.A1(n_9), .A2(n_0_336), .B1(A_imm_2s_complement[13]), 
      .B2(n_0_311), .ZN(n_0_233));
   OAI221_X1 i_0_478 (.A(n_0_234), .B1(n_0_359), .B2(n_0_338), .C1(n_0_382), 
      .C2(n_0_340), .ZN(n_281));
   AOI22_X1 i_0_479 (.A1(n_8), .A2(n_0_336), .B1(A_imm_2s_complement[14]), 
      .B2(n_0_311), .ZN(n_0_234));
   OAI221_X1 i_0_480 (.A(n_0_235), .B1(n_0_360), .B2(n_0_338), .C1(n_0_383), 
      .C2(n_0_340), .ZN(n_282));
   AOI22_X1 i_0_481 (.A1(n_7), .A2(n_0_336), .B1(A_imm_2s_complement[15]), 
      .B2(n_0_311), .ZN(n_0_235));
   OAI221_X1 i_0_482 (.A(n_0_236), .B1(n_0_361), .B2(n_0_338), .C1(n_0_384), 
      .C2(n_0_340), .ZN(n_283));
   AOI22_X1 i_0_483 (.A1(n_6), .A2(n_0_336), .B1(A_imm_2s_complement[16]), 
      .B2(n_0_311), .ZN(n_0_236));
   OAI221_X1 i_0_110 (.A(n_0_237), .B1(n_0_310), .B2(n_0_338), .C1(n_0_385), 
      .C2(n_0_340), .ZN(n_284));
   AOI22_X1 i_0_111 (.A1(n_5), .A2(n_0_336), .B1(A_imm_2s_complement[17]), 
      .B2(n_0_311), .ZN(n_0_237));
   OAI221_X1 i_0_486 (.A(n_0_238), .B1(n_0_363), .B2(n_0_338), .C1(n_0_386), 
      .C2(n_0_340), .ZN(n_285));
   AOI22_X1 i_0_487 (.A1(n_4), .A2(n_0_336), .B1(A_imm_2s_complement[18]), 
      .B2(n_0_311), .ZN(n_0_238));
   OAI221_X1 i_0_488 (.A(n_0_239), .B1(n_0_404), .B2(n_0_338), .C1(n_0_403), 
      .C2(n_0_340), .ZN(n_286));
   AOI22_X1 i_0_489 (.A1(n_3), .A2(n_0_336), .B1(A_imm_2s_complement[19]), 
      .B2(n_0_311), .ZN(n_0_239));
   OAI221_X1 i_0_490 (.A(n_0_240), .B1(n_0_365), .B2(n_0_338), .C1(n_0_388), 
      .C2(n_0_340), .ZN(n_287));
   AOI22_X1 i_0_491 (.A1(n_2), .A2(n_0_336), .B1(A_imm_2s_complement[20]), 
      .B2(n_0_311), .ZN(n_0_240));
   OAI221_X1 i_0_492 (.A(n_0_241), .B1(n_0_31), .B2(n_0_338), .C1(n_0_27), 
      .C2(n_0_340), .ZN(n_288));
   AOI22_X1 i_0_493 (.A1(n_1), .A2(n_0_336), .B1(A_imm_2s_complement[21]), 
      .B2(n_0_311), .ZN(n_0_241));
   OAI221_X1 i_0_494 (.A(n_0_242), .B1(n_0_28), .B2(n_0_338), .C1(n_0_60), 
      .C2(n_0_340), .ZN(n_289));
   AOI22_X1 i_0_495 (.A1(n_0), .A2(n_0_336), .B1(A_imm_2s_complement[22]), 
      .B2(n_0_311), .ZN(n_0_242));
   OAI222_X1 i_0_497 (.A1(n_0_60), .A2(n_0_246), .B1(n_0_28), .B2(n_0_334), 
      .C1(n_0_391), .C2(n_0_340), .ZN(n_290));
   INV_X1 i_0_500 (.A(n_0_311), .ZN(n_0_246));
   NOR3_X1 i_0_504 (.A1(n_0_268), .A2(n_0_391), .A3(n_0_330), .ZN(n_291));
   NOR2_X1 i_0_506 (.A1(n_0_344), .A2(n_0_366), .ZN(n_292));
   OAI221_X1 i_0_509 (.A(n_0_252), .B1(n_0_346), .B2(n_0_381), .C1(n_0_369), 
      .C2(n_0_368), .ZN(n_293));
   AOI22_X1 i_0_510 (.A1(n_21), .A2(n_0_364), .B1(A_imm_2s_complement[1]), 
      .B2(n_0_342), .ZN(n_0_252));
   OAI221_X1 i_0_511 (.A(n_0_253), .B1(n_0_347), .B2(n_0_381), .C1(n_0_370), 
      .C2(n_0_368), .ZN(n_294));
   AOI22_X1 i_0_512 (.A1(n_20), .A2(n_0_364), .B1(A_imm_2s_complement[2]), 
      .B2(n_0_342), .ZN(n_0_253));
   OAI221_X1 i_0_513 (.A(n_0_254), .B1(n_0_348), .B2(n_0_381), .C1(n_0_371), 
      .C2(n_0_368), .ZN(n_295));
   AOI22_X1 i_0_514 (.A1(n_19), .A2(n_0_364), .B1(A_imm_2s_complement[3]), 
      .B2(n_0_342), .ZN(n_0_254));
   OAI221_X1 i_0_515 (.A(n_0_255), .B1(n_0_349), .B2(n_0_381), .C1(n_0_372), 
      .C2(n_0_368), .ZN(n_296));
   AOI22_X1 i_0_516 (.A1(n_18), .A2(n_0_364), .B1(A_imm_2s_complement[4]), 
      .B2(n_0_342), .ZN(n_0_255));
   OAI221_X1 i_0_517 (.A(n_0_256), .B1(n_0_350), .B2(n_0_381), .C1(n_0_373), 
      .C2(n_0_368), .ZN(n_297));
   AOI22_X1 i_0_518 (.A1(n_17), .A2(n_0_364), .B1(A_imm_2s_complement[5]), 
      .B2(n_0_342), .ZN(n_0_256));
   OAI221_X1 i_0_519 (.A(n_0_257), .B1(n_0_351), .B2(n_0_381), .C1(n_0_374), 
      .C2(n_0_368), .ZN(n_298));
   AOI22_X1 i_0_520 (.A1(n_16), .A2(n_0_364), .B1(A_imm_2s_complement[6]), 
      .B2(n_0_342), .ZN(n_0_257));
   OAI221_X1 i_0_521 (.A(n_0_258), .B1(n_0_352), .B2(n_0_381), .C1(n_0_375), 
      .C2(n_0_368), .ZN(n_299));
   AOI22_X1 i_0_522 (.A1(n_15), .A2(n_0_364), .B1(A_imm_2s_complement[7]), 
      .B2(n_0_342), .ZN(n_0_258));
   OAI221_X1 i_0_523 (.A(n_0_259), .B1(n_0_353), .B2(n_0_381), .C1(n_0_376), 
      .C2(n_0_368), .ZN(n_300));
   AOI22_X1 i_0_524 (.A1(n_14), .A2(n_0_364), .B1(A_imm_2s_complement[8]), 
      .B2(n_0_342), .ZN(n_0_259));
   OAI221_X1 i_0_525 (.A(n_0_260), .B1(n_0_354), .B2(n_0_381), .C1(n_0_377), 
      .C2(n_0_368), .ZN(n_301));
   AOI22_X1 i_0_526 (.A1(n_13), .A2(n_0_364), .B1(A_imm_2s_complement[9]), 
      .B2(n_0_342), .ZN(n_0_260));
   OAI221_X1 i_0_527 (.A(n_0_261), .B1(n_0_355), .B2(n_0_381), .C1(n_0_378), 
      .C2(n_0_368), .ZN(n_302));
   AOI22_X1 i_0_528 (.A1(n_12), .A2(n_0_364), .B1(A_imm_2s_complement[10]), 
      .B2(n_0_342), .ZN(n_0_261));
   OAI221_X1 i_0_529 (.A(n_0_262), .B1(n_0_356), .B2(n_0_381), .C1(n_0_379), 
      .C2(n_0_368), .ZN(n_303));
   AOI22_X1 i_0_530 (.A1(n_11), .A2(n_0_364), .B1(A_imm_2s_complement[11]), 
      .B2(n_0_342), .ZN(n_0_262));
   OAI221_X1 i_0_531 (.A(n_0_263), .B1(n_0_357), .B2(n_0_381), .C1(n_0_380), 
      .C2(n_0_368), .ZN(n_304));
   AOI22_X1 i_0_532 (.A1(n_10), .A2(n_0_364), .B1(A_imm_2s_complement[12]), 
      .B2(n_0_342), .ZN(n_0_263));
   OAI221_X1 i_0_533 (.A(n_0_264), .B1(n_0_306), .B2(n_0_381), .C1(n_0_305), 
      .C2(n_0_368), .ZN(n_305));
   AOI22_X1 i_0_534 (.A1(n_9), .A2(n_0_364), .B1(A_imm_2s_complement[13]), 
      .B2(n_0_342), .ZN(n_0_264));
   OAI221_X1 i_0_535 (.A(n_0_265), .B1(n_0_359), .B2(n_0_381), .C1(n_0_382), 
      .C2(n_0_368), .ZN(n_306));
   AOI22_X1 i_0_536 (.A1(n_8), .A2(n_0_364), .B1(A_imm_2s_complement[14]), 
      .B2(n_0_342), .ZN(n_0_265));
   OAI221_X1 i_0_537 (.A(n_0_266), .B1(n_0_360), .B2(n_0_381), .C1(n_0_383), 
      .C2(n_0_368), .ZN(n_307));
   AOI22_X1 i_0_538 (.A1(n_7), .A2(n_0_364), .B1(A_imm_2s_complement[15]), 
      .B2(n_0_342), .ZN(n_0_266));
   OAI221_X1 i_0_539 (.A(n_0_267), .B1(n_0_361), .B2(n_0_381), .C1(n_0_384), 
      .C2(n_0_368), .ZN(n_308));
   AOI22_X1 i_0_540 (.A1(n_6), .A2(n_0_364), .B1(A_imm_2s_complement[16]), 
      .B2(n_0_342), .ZN(n_0_267));
   OAI221_X1 i_0_543 (.A(n_0_269), .B1(n_0_363), .B2(n_0_381), .C1(n_0_386), 
      .C2(n_0_368), .ZN(n_309));
   AOI22_X1 i_0_544 (.A1(n_4), .A2(n_0_364), .B1(A_imm_2s_complement[18]), 
      .B2(n_0_342), .ZN(n_0_269));
   OAI221_X1 i_0_545 (.A(n_0_270), .B1(n_0_404), .B2(n_0_381), .C1(n_0_403), 
      .C2(n_0_368), .ZN(n_310));
   AOI22_X1 i_0_546 (.A1(n_3), .A2(n_0_364), .B1(A_imm_2s_complement[19]), 
      .B2(n_0_342), .ZN(n_0_270));
   OAI221_X1 i_0_547 (.A(n_0_271), .B1(n_0_365), .B2(n_0_381), .C1(n_0_388), 
      .C2(n_0_368), .ZN(n_311));
   AOI22_X1 i_0_548 (.A1(n_2), .A2(n_0_364), .B1(A_imm_2s_complement[20]), 
      .B2(n_0_342), .ZN(n_0_271));
   OAI221_X1 i_0_549 (.A(n_0_272), .B1(n_0_31), .B2(n_0_381), .C1(n_0_27), 
      .C2(n_0_368), .ZN(n_312));
   AOI22_X1 i_0_550 (.A1(n_1), .A2(n_0_364), .B1(A_imm_2s_complement[21]), 
      .B2(n_0_342), .ZN(n_0_272));
   OAI221_X1 i_0_551 (.A(n_0_273), .B1(n_0_28), .B2(n_0_381), .C1(n_0_60), 
      .C2(n_0_368), .ZN(n_313));
   AOI22_X1 i_0_552 (.A1(n_0), .A2(n_0_364), .B1(A_imm_2s_complement[22]), 
      .B2(n_0_342), .ZN(n_0_273));
   OAI222_X1 i_0_554 (.A1(n_0_60), .A2(n_0_277), .B1(n_0_28), .B2(n_0_362), 
      .C1(n_0_391), .C2(n_0_368), .ZN(n_314));
   INV_X1 i_0_557 (.A(n_0_342), .ZN(n_0_277));
   NOR3_X1 i_0_561 (.A1(n_0_312), .A2(n_0_391), .A3(n_0_358), .ZN(n_315));
   NOR2_X1 i_0_563 (.A1(n_0_344), .A2(n_0_397), .ZN(n_316));
   OAI221_X1 i_0_566 (.A(n_0_283), .B1(n_0_346), .B2(n_0_400), .C1(n_0_369), 
      .C2(n_0_399), .ZN(n_317));
   AOI22_X1 i_0_567 (.A1(n_21), .A2(n_0_396), .B1(A_imm_2s_complement[1]), 
      .B2(n_0_390), .ZN(n_0_283));
   OAI221_X1 i_0_568 (.A(n_0_284), .B1(n_0_347), .B2(n_0_400), .C1(n_0_370), 
      .C2(n_0_399), .ZN(n_318));
   AOI22_X1 i_0_569 (.A1(n_20), .A2(n_0_396), .B1(A_imm_2s_complement[2]), 
      .B2(n_0_390), .ZN(n_0_284));
   OAI221_X1 i_0_570 (.A(n_0_285), .B1(n_0_348), .B2(n_0_400), .C1(n_0_371), 
      .C2(n_0_399), .ZN(n_319));
   AOI22_X1 i_0_571 (.A1(n_19), .A2(n_0_396), .B1(A_imm_2s_complement[3]), 
      .B2(n_0_390), .ZN(n_0_285));
   OAI221_X1 i_0_572 (.A(n_0_286), .B1(n_0_349), .B2(n_0_400), .C1(n_0_372), 
      .C2(n_0_399), .ZN(n_320));
   AOI22_X1 i_0_573 (.A1(n_18), .A2(n_0_396), .B1(A_imm_2s_complement[4]), 
      .B2(n_0_390), .ZN(n_0_286));
   OAI221_X1 i_0_574 (.A(n_0_287), .B1(n_0_350), .B2(n_0_400), .C1(n_0_373), 
      .C2(n_0_399), .ZN(n_321));
   AOI22_X1 i_0_575 (.A1(n_17), .A2(n_0_396), .B1(A_imm_2s_complement[5]), 
      .B2(n_0_390), .ZN(n_0_287));
   OAI221_X1 i_0_576 (.A(n_0_288), .B1(n_0_351), .B2(n_0_400), .C1(n_0_374), 
      .C2(n_0_399), .ZN(n_322));
   AOI22_X1 i_0_577 (.A1(n_16), .A2(n_0_396), .B1(A_imm_2s_complement[6]), 
      .B2(n_0_390), .ZN(n_0_288));
   OAI221_X1 i_0_578 (.A(n_0_289), .B1(n_0_352), .B2(n_0_400), .C1(n_0_375), 
      .C2(n_0_399), .ZN(n_323));
   AOI22_X1 i_0_579 (.A1(n_15), .A2(n_0_396), .B1(A_imm_2s_complement[7]), 
      .B2(n_0_390), .ZN(n_0_289));
   OAI221_X1 i_0_580 (.A(n_0_290), .B1(n_0_353), .B2(n_0_400), .C1(n_0_376), 
      .C2(n_0_399), .ZN(n_324));
   AOI22_X1 i_0_581 (.A1(n_14), .A2(n_0_396), .B1(A_imm_2s_complement[8]), 
      .B2(n_0_390), .ZN(n_0_290));
   OAI221_X1 i_0_582 (.A(n_0_291), .B1(n_0_354), .B2(n_0_400), .C1(n_0_377), 
      .C2(n_0_399), .ZN(n_325));
   AOI22_X1 i_0_583 (.A1(n_13), .A2(n_0_396), .B1(A_imm_2s_complement[9]), 
      .B2(n_0_390), .ZN(n_0_291));
   OAI221_X1 i_0_584 (.A(n_0_292), .B1(n_0_355), .B2(n_0_400), .C1(n_0_378), 
      .C2(n_0_399), .ZN(n_326));
   AOI22_X1 i_0_585 (.A1(n_12), .A2(n_0_396), .B1(A_imm_2s_complement[10]), 
      .B2(n_0_390), .ZN(n_0_292));
   OAI221_X1 i_0_586 (.A(n_0_293), .B1(n_0_356), .B2(n_0_400), .C1(n_0_379), 
      .C2(n_0_399), .ZN(n_327));
   AOI22_X1 i_0_587 (.A1(n_11), .A2(n_0_396), .B1(A_imm_2s_complement[11]), 
      .B2(n_0_390), .ZN(n_0_293));
   OAI221_X1 i_0_588 (.A(n_0_294), .B1(n_0_357), .B2(n_0_400), .C1(n_0_380), 
      .C2(n_0_399), .ZN(n_328));
   AOI22_X1 i_0_589 (.A1(n_10), .A2(n_0_396), .B1(A_imm_2s_complement[12]), 
      .B2(n_0_390), .ZN(n_0_294));
   OAI221_X1 i_0_590 (.A(n_0_295), .B1(n_0_306), .B2(n_0_400), .C1(n_0_305), 
      .C2(n_0_399), .ZN(n_329));
   AOI22_X1 i_0_591 (.A1(n_9), .A2(n_0_396), .B1(A_imm_2s_complement[13]), 
      .B2(n_0_390), .ZN(n_0_295));
   OAI221_X1 i_0_592 (.A(n_0_296), .B1(n_0_359), .B2(n_0_400), .C1(n_0_382), 
      .C2(n_0_399), .ZN(n_330));
   AOI22_X1 i_0_593 (.A1(n_8), .A2(n_0_396), .B1(A_imm_2s_complement[14]), 
      .B2(n_0_390), .ZN(n_0_296));
   OAI221_X1 i_0_594 (.A(n_0_297), .B1(n_0_360), .B2(n_0_400), .C1(n_0_383), 
      .C2(n_0_399), .ZN(n_331));
   AOI22_X1 i_0_595 (.A1(n_7), .A2(n_0_396), .B1(A_imm_2s_complement[15]), 
      .B2(n_0_390), .ZN(n_0_297));
   OAI221_X1 i_0_596 (.A(n_0_298), .B1(n_0_361), .B2(n_0_400), .C1(n_0_384), 
      .C2(n_0_399), .ZN(n_332));
   AOI22_X1 i_0_597 (.A1(n_6), .A2(n_0_396), .B1(A_imm_2s_complement[16]), 
      .B2(n_0_390), .ZN(n_0_298));
   OAI221_X1 i_0_598 (.A(n_0_299), .B1(n_0_310), .B2(n_0_400), .C1(n_0_385), 
      .C2(n_0_399), .ZN(n_333));
   AOI22_X1 i_0_599 (.A1(n_5), .A2(n_0_396), .B1(A_imm_2s_complement[17]), 
      .B2(n_0_390), .ZN(n_0_299));
   OAI221_X1 i_0_600 (.A(n_0_300), .B1(n_0_363), .B2(n_0_400), .C1(n_0_386), 
      .C2(n_0_399), .ZN(n_334));
   AOI22_X1 i_0_601 (.A1(n_4), .A2(n_0_396), .B1(A_imm_2s_complement[18]), 
      .B2(n_0_390), .ZN(n_0_300));
   OAI221_X1 i_0_604 (.A(n_0_302), .B1(n_0_365), .B2(n_0_400), .C1(n_0_388), 
      .C2(n_0_399), .ZN(n_335));
   AOI22_X1 i_0_605 (.A1(n_2), .A2(n_0_396), .B1(A_imm_2s_complement[20]), 
      .B2(n_0_390), .ZN(n_0_302));
   OAI221_X1 i_0_606 (.A(n_0_303), .B1(n_0_31), .B2(n_0_400), .C1(n_0_27), 
      .C2(n_0_399), .ZN(n_336));
   AOI22_X1 i_0_607 (.A1(n_1), .A2(n_0_396), .B1(A_imm_2s_complement[21]), 
      .B2(n_0_390), .ZN(n_0_303));
   OAI222_X1 i_0_611 (.A1(n_0_60), .A2(n_0_308), .B1(n_0_28), .B2(n_0_395), 
      .C1(n_0_391), .C2(n_0_399), .ZN(n_337));
   INV_X1 i_0_614 (.A(n_0_390), .ZN(n_0_308));
   NOR3_X1 i_0_618 (.A1(n_0_343), .A2(n_0_391), .A3(n_0_394), .ZN(n_338));
   NOR2_X1 i_0_620 (.A1(n_0_344), .A2(n_0_412), .ZN(n_339));
   OAI221_X1 i_0_623 (.A(n_0_314), .B1(n_0_346), .B2(n_0_415), .C1(n_0_369), 
      .C2(n_0_414), .ZN(n_340));
   AOI22_X1 i_0_624 (.A1(n_21), .A2(n_0_411), .B1(A_imm_2s_complement[1]), 
      .B2(n_0_406), .ZN(n_0_314));
   OAI221_X1 i_0_625 (.A(n_0_315), .B1(n_0_347), .B2(n_0_415), .C1(n_0_370), 
      .C2(n_0_414), .ZN(n_341));
   AOI22_X1 i_0_626 (.A1(n_20), .A2(n_0_411), .B1(A_imm_2s_complement[2]), 
      .B2(n_0_406), .ZN(n_0_315));
   OAI221_X1 i_0_627 (.A(n_0_316), .B1(n_0_348), .B2(n_0_415), .C1(n_0_371), 
      .C2(n_0_414), .ZN(n_342));
   AOI22_X1 i_0_628 (.A1(n_19), .A2(n_0_411), .B1(A_imm_2s_complement[3]), 
      .B2(n_0_406), .ZN(n_0_316));
   OAI221_X1 i_0_629 (.A(n_0_317), .B1(n_0_349), .B2(n_0_415), .C1(n_0_372), 
      .C2(n_0_414), .ZN(n_343));
   AOI22_X1 i_0_630 (.A1(n_18), .A2(n_0_411), .B1(A_imm_2s_complement[4]), 
      .B2(n_0_406), .ZN(n_0_317));
   OAI221_X1 i_0_631 (.A(n_0_318), .B1(n_0_350), .B2(n_0_415), .C1(n_0_373), 
      .C2(n_0_414), .ZN(n_344));
   AOI22_X1 i_0_632 (.A1(n_17), .A2(n_0_411), .B1(A_imm_2s_complement[5]), 
      .B2(n_0_406), .ZN(n_0_318));
   OAI221_X1 i_0_633 (.A(n_0_319), .B1(n_0_351), .B2(n_0_415), .C1(n_0_374), 
      .C2(n_0_414), .ZN(n_345));
   AOI22_X1 i_0_634 (.A1(n_16), .A2(n_0_411), .B1(A_imm_2s_complement[6]), 
      .B2(n_0_406), .ZN(n_0_319));
   OAI221_X1 i_0_635 (.A(n_0_320), .B1(n_0_352), .B2(n_0_415), .C1(n_0_375), 
      .C2(n_0_414), .ZN(n_346));
   AOI22_X1 i_0_636 (.A1(n_15), .A2(n_0_411), .B1(A_imm_2s_complement[7]), 
      .B2(n_0_406), .ZN(n_0_320));
   OAI221_X1 i_0_637 (.A(n_0_321), .B1(n_0_353), .B2(n_0_415), .C1(n_0_376), 
      .C2(n_0_414), .ZN(n_347));
   AOI22_X1 i_0_638 (.A1(n_14), .A2(n_0_411), .B1(A_imm_2s_complement[8]), 
      .B2(n_0_406), .ZN(n_0_321));
   OAI221_X1 i_0_639 (.A(n_0_322), .B1(n_0_354), .B2(n_0_415), .C1(n_0_377), 
      .C2(n_0_414), .ZN(n_348));
   AOI22_X1 i_0_640 (.A1(n_13), .A2(n_0_411), .B1(A_imm_2s_complement[9]), 
      .B2(n_0_406), .ZN(n_0_322));
   OAI221_X1 i_0_641 (.A(n_0_323), .B1(n_0_355), .B2(n_0_415), .C1(n_0_378), 
      .C2(n_0_414), .ZN(n_349));
   AOI22_X1 i_0_642 (.A1(n_12), .A2(n_0_411), .B1(A_imm_2s_complement[10]), 
      .B2(n_0_406), .ZN(n_0_323));
   OAI221_X1 i_0_643 (.A(n_0_324), .B1(n_0_356), .B2(n_0_415), .C1(n_0_379), 
      .C2(n_0_414), .ZN(n_350));
   AOI22_X1 i_0_644 (.A1(n_11), .A2(n_0_411), .B1(A_imm_2s_complement[11]), 
      .B2(n_0_406), .ZN(n_0_324));
   OAI221_X1 i_0_645 (.A(n_0_325), .B1(n_0_357), .B2(n_0_415), .C1(n_0_380), 
      .C2(n_0_414), .ZN(n_351));
   AOI22_X1 i_0_646 (.A1(n_10), .A2(n_0_411), .B1(A_imm_2s_complement[12]), 
      .B2(n_0_406), .ZN(n_0_325));
   OAI221_X1 i_0_647 (.A(n_0_326), .B1(n_0_306), .B2(n_0_415), .C1(n_0_305), 
      .C2(n_0_414), .ZN(n_352));
   AOI22_X1 i_0_648 (.A1(n_9), .A2(n_0_411), .B1(A_imm_2s_complement[13]), 
      .B2(n_0_406), .ZN(n_0_326));
   OAI221_X1 i_0_649 (.A(n_0_327), .B1(n_0_359), .B2(n_0_415), .C1(n_0_382), 
      .C2(n_0_414), .ZN(n_353));
   AOI22_X1 i_0_650 (.A1(n_8), .A2(n_0_411), .B1(A_imm_2s_complement[14]), 
      .B2(n_0_406), .ZN(n_0_327));
   OAI221_X1 i_0_651 (.A(n_0_328), .B1(n_0_360), .B2(n_0_415), .C1(n_0_383), 
      .C2(n_0_414), .ZN(n_354));
   AOI22_X1 i_0_652 (.A1(n_7), .A2(n_0_411), .B1(A_imm_2s_complement[15]), 
      .B2(n_0_406), .ZN(n_0_328));
   OAI221_X1 i_0_653 (.A(n_0_329), .B1(n_0_361), .B2(n_0_415), .C1(n_0_384), 
      .C2(n_0_414), .ZN(n_355));
   AOI22_X1 i_0_654 (.A1(n_6), .A2(n_0_411), .B1(A_imm_2s_complement[16]), 
      .B2(n_0_406), .ZN(n_0_329));
   OAI221_X1 i_0_657 (.A(n_0_331), .B1(n_0_363), .B2(n_0_415), .C1(n_0_386), 
      .C2(n_0_414), .ZN(n_356));
   AOI22_X1 i_0_658 (.A1(n_4), .A2(n_0_411), .B1(A_imm_2s_complement[18]), 
      .B2(n_0_406), .ZN(n_0_331));
   OAI221_X1 i_0_659 (.A(n_0_332), .B1(n_0_404), .B2(n_0_415), .C1(n_0_403), 
      .C2(n_0_414), .ZN(n_357));
   AOI22_X1 i_0_660 (.A1(n_3), .A2(n_0_411), .B1(A_imm_2s_complement[19]), 
      .B2(n_0_406), .ZN(n_0_332));
   OAI221_X1 i_0_661 (.A(n_0_333), .B1(n_0_365), .B2(n_0_415), .C1(n_0_388), 
      .C2(n_0_414), .ZN(n_358));
   AOI22_X1 i_0_662 (.A1(n_2), .A2(n_0_411), .B1(A_imm_2s_complement[20]), 
      .B2(n_0_406), .ZN(n_0_333));
   OAI221_X1 i_0_665 (.A(n_0_335), .B1(n_0_28), .B2(n_0_415), .C1(n_0_60), 
      .C2(n_0_414), .ZN(n_359));
   AOI22_X1 i_0_666 (.A1(n_0), .A2(n_0_411), .B1(A_imm_2s_complement[22]), 
      .B2(n_0_406), .ZN(n_0_335));
   OAI222_X1 i_0_668 (.A1(n_0_60), .A2(n_0_339), .B1(n_0_28), .B2(n_0_410), 
      .C1(n_0_391), .C2(n_0_414), .ZN(n_360));
   INV_X1 i_0_671 (.A(n_0_406), .ZN(n_0_339));
   NOR3_X1 i_0_675 (.A1(n_0_392), .A2(n_0_391), .A3(n_0_409), .ZN(n_361));
   INV_X1 i_0_150 (.A(n_22), .ZN(n_0_344));
   INV_X1 i_0_151 (.A(n_20), .ZN(n_0_346));
   INV_X1 i_0_680 (.A(n_19), .ZN(n_0_347));
   INV_X1 i_0_681 (.A(n_18), .ZN(n_0_348));
   INV_X1 i_0_682 (.A(n_17), .ZN(n_0_349));
   INV_X1 i_0_683 (.A(n_16), .ZN(n_0_350));
   INV_X1 i_0_684 (.A(n_15), .ZN(n_0_351));
   INV_X1 i_0_685 (.A(n_14), .ZN(n_0_352));
   INV_X1 i_0_686 (.A(n_13), .ZN(n_0_353));
   INV_X1 i_0_687 (.A(n_12), .ZN(n_0_354));
   INV_X1 i_0_688 (.A(n_11), .ZN(n_0_355));
   INV_X1 i_0_689 (.A(n_10), .ZN(n_0_356));
   INV_X1 i_0_690 (.A(n_9), .ZN(n_0_357));
   INV_X1 i_0_692 (.A(n_7), .ZN(n_0_359));
   INV_X1 i_0_693 (.A(n_6), .ZN(n_0_360));
   INV_X1 i_0_694 (.A(n_5), .ZN(n_0_361));
   INV_X1 i_0_696 (.A(n_3), .ZN(n_0_363));
   INV_X1 i_0_698 (.A(n_1), .ZN(n_0_365));
   INV_X1 i_0_154 (.A(A_imm_2s_complement[2]), .ZN(n_0_369));
   INV_X1 i_0_703 (.A(A_imm_2s_complement[3]), .ZN(n_0_370));
   INV_X1 i_0_704 (.A(A_imm_2s_complement[4]), .ZN(n_0_371));
   INV_X1 i_0_705 (.A(A_imm_2s_complement[5]), .ZN(n_0_372));
   INV_X1 i_0_706 (.A(A_imm_2s_complement[6]), .ZN(n_0_373));
   INV_X1 i_0_707 (.A(A_imm_2s_complement[7]), .ZN(n_0_374));
   INV_X1 i_0_708 (.A(A_imm_2s_complement[8]), .ZN(n_0_375));
   INV_X1 i_0_709 (.A(A_imm_2s_complement[9]), .ZN(n_0_376));
   INV_X1 i_0_710 (.A(A_imm_2s_complement[10]), .ZN(n_0_377));
   INV_X1 i_0_711 (.A(A_imm_2s_complement[11]), .ZN(n_0_378));
   INV_X1 i_0_712 (.A(A_imm_2s_complement[12]), .ZN(n_0_379));
   INV_X1 i_0_713 (.A(A_imm_2s_complement[13]), .ZN(n_0_380));
   INV_X1 i_0_715 (.A(A_imm_2s_complement[15]), .ZN(n_0_382));
   INV_X1 i_0_716 (.A(A_imm_2s_complement[16]), .ZN(n_0_383));
   INV_X1 i_0_717 (.A(A_imm_2s_complement[17]), .ZN(n_0_384));
   INV_X1 i_0_719 (.A(A_imm_2s_complement[19]), .ZN(n_0_386));
   INV_X1 i_0_721 (.A(A_imm_2s_complement[21]), .ZN(n_0_388));
   INV_X1 i_0_155 (.A(A_imm_2s_complement[27]), .ZN(n_0_391));
   INV_X1 i_0_156 (.A(A_imm_2s_complement[18]), .ZN(n_0_385));
   INV_X1 i_0_157 (.A(A_imm_2s_complement[22]), .ZN(n_0_27));
   INV_X1 i_0_158 (.A(n_46), .ZN(n_0_28));
   NOR3_X1 i_0_159 (.A1(n_0_28), .A2(n_23), .A3(n_24), .ZN(n_0_29));
   INV_X1 i_0_160 (.A(n_0_29), .ZN(n_0_30));
   INV_X1 i_0_161 (.A(n_0), .ZN(n_0_31));
   INV_X1 i_0_162 (.A(n_24), .ZN(n_0_33));
   NAND2_X1 i_0_163 (.A1(n_23), .A2(n_24), .ZN(n_0_34));
   INV_X1 i_0_165 (.A(n_0_34), .ZN(n_0_57));
   NAND2_X1 i_0_166 (.A1(n_0_57), .A2(n_0_28), .ZN(n_0_59));
   INV_X1 i_0_211 (.A(A_imm_2s_complement[23]), .ZN(n_0_60));
   OAI21_X1 i_0_214 (.A(n_0_34), .B1(n_23), .B2(n_24), .ZN(n_0_61));
   OR2_X1 i_0_215 (.A1(n_0_61), .A2(n_0_28), .ZN(n_0_62));
   OAI222_X1 i_0_216 (.A1(n_0_62), .A2(n_0_60), .B1(n_0_30), .B2(n_0_27), 
      .C1(n_0_59), .C2(n_0_31), .ZN(n_362));
   INV_X1 i_0_217 (.A(n_26), .ZN(n_0_63));
   NAND2_X1 i_0_218 (.A1(n_25), .A2(n_26), .ZN(n_0_64));
   INV_X1 i_0_220 (.A(n_0_64), .ZN(n_0_65));
   NAND2_X1 i_0_222 (.A1(n_0_65), .A2(n_0_33), .ZN(n_0_88));
   INV_X1 i_0_223 (.A(n_0_88), .ZN(n_0_90));
   NOR3_X1 i_0_268 (.A1(n_25), .A2(n_26), .A3(n_0_33), .ZN(n_0_91));
   INV_X1 i_0_269 (.A(A_imm_2s_complement[1]), .ZN(n_0_92));
   OAI21_X1 i_0_270 (.A(n_0_64), .B1(n_25), .B2(n_26), .ZN(n_0_93));
   OR2_X1 i_0_271 (.A1(n_0_93), .A2(n_0_33), .ZN(n_0_94));
   INV_X1 i_0_272 (.A(n_21), .ZN(n_0_95));
   OR2_X1 i_0_273 (.A1(n_0_93), .A2(n_24), .ZN(n_0_96));
   OAI21_X1 i_0_274 (.A(n_22), .B1(n_0_90), .B2(n_0_91), .ZN(n_0_119));
   OAI221_X1 i_0_275 (.A(n_0_119), .B1(n_0_96), .B2(n_0_95), .C1(n_0_94), 
      .C2(n_0_92), .ZN(n_363));
   INV_X1 i_0_277 (.A(n_28), .ZN(n_0_120));
   NAND2_X1 i_0_279 (.A1(n_27), .A2(n_28), .ZN(n_0_121));
   INV_X1 i_0_280 (.A(n_0_121), .ZN(n_0_123));
   NAND2_X1 i_0_325 (.A1(n_0_123), .A2(n_0_63), .ZN(n_0_124));
   INV_X1 i_0_327 (.A(n_0_124), .ZN(n_0_125));
   NOR3_X1 i_0_328 (.A1(n_27), .A2(n_28), .A3(n_0_63), .ZN(n_0_126));
   OAI21_X1 i_0_330 (.A(n_0_121), .B1(n_27), .B2(n_28), .ZN(n_0_127));
   OR2_X1 i_0_331 (.A1(n_0_127), .A2(n_0_63), .ZN(n_0_150));
   OR2_X1 i_0_332 (.A1(n_0_127), .A2(n_26), .ZN(n_0_151));
   OAI21_X1 i_0_334 (.A(n_22), .B1(n_0_125), .B2(n_0_126), .ZN(n_0_152));
   OAI221_X1 i_0_336 (.A(n_0_152), .B1(n_0_151), .B2(n_0_95), .C1(n_0_150), 
      .C2(n_0_92), .ZN(n_364));
   NOR3_X1 i_0_337 (.A1(n_29), .A2(n_30), .A3(n_0_120), .ZN(n_0_154));
   INV_X1 i_0_382 (.A(n_30), .ZN(n_0_155));
   NAND2_X1 i_0_384 (.A1(n_29), .A2(n_30), .ZN(n_0_156));
   INV_X1 i_0_385 (.A(n_0_156), .ZN(n_0_157));
   NAND2_X1 i_0_387 (.A1(n_0_157), .A2(n_0_120), .ZN(n_0_158));
   INV_X1 i_0_388 (.A(n_0_158), .ZN(n_0_181));
   OAI21_X1 i_0_389 (.A(n_0_156), .B1(n_29), .B2(n_30), .ZN(n_0_182));
   OR2_X1 i_0_391 (.A1(n_0_182), .A2(n_28), .ZN(n_0_183));
   OR2_X1 i_0_393 (.A1(n_0_182), .A2(n_0_120), .ZN(n_0_185));
   OAI21_X1 i_0_394 (.A(n_22), .B1(n_0_181), .B2(n_0_154), .ZN(n_0_186));
   OAI221_X1 i_0_419 (.A(n_0_186), .B1(n_0_183), .B2(n_0_95), .C1(n_0_185), 
      .C2(n_0_92), .ZN(n_365));
   NOR3_X1 i_0_420 (.A1(n_31), .A2(n_32), .A3(n_0_155), .ZN(n_0_187));
   INV_X1 i_0_427 (.A(n_32), .ZN(n_0_188));
   NAND2_X1 i_0_428 (.A1(n_31), .A2(n_32), .ZN(n_0_189));
   INV_X1 i_0_439 (.A(n_0_189), .ZN(n_0_202));
   NAND2_X1 i_0_441 (.A1(n_0_202), .A2(n_0_155), .ZN(n_0_206));
   INV_X1 i_0_442 (.A(n_0_206), .ZN(n_0_212));
   OAI21_X1 i_0_444 (.A(n_0_189), .B1(n_31), .B2(n_32), .ZN(n_0_213));
   OR2_X1 i_0_445 (.A1(n_0_213), .A2(n_30), .ZN(n_0_214));
   OR2_X1 i_0_446 (.A1(n_0_213), .A2(n_0_155), .ZN(n_0_216));
   OAI21_X1 i_0_448 (.A(n_22), .B1(n_0_212), .B2(n_0_187), .ZN(n_0_217));
   OAI221_X1 i_0_450 (.A(n_0_217), .B1(n_0_214), .B2(n_0_95), .C1(n_0_216), 
      .C2(n_0_92), .ZN(n_366));
   NOR3_X1 i_0_451 (.A1(n_33), .A2(n_34), .A3(n_0_188), .ZN(n_0_218));
   INV_X1 i_0_484 (.A(n_34), .ZN(n_0_219));
   NAND2_X1 i_0_485 (.A1(n_33), .A2(n_34), .ZN(n_0_220));
   INV_X1 i_0_496 (.A(n_0_220), .ZN(n_0_243));
   NAND2_X1 i_0_498 (.A1(n_0_243), .A2(n_0_188), .ZN(n_0_244));
   INV_X1 i_0_499 (.A(n_0_244), .ZN(n_0_245));
   OAI21_X1 i_0_501 (.A(n_0_220), .B1(n_33), .B2(n_34), .ZN(n_0_247));
   OR2_X1 i_0_502 (.A1(n_0_247), .A2(n_32), .ZN(n_0_248));
   OR2_X1 i_0_503 (.A1(n_0_247), .A2(n_0_188), .ZN(n_0_249));
   OAI21_X1 i_0_505 (.A(n_22), .B1(n_0_245), .B2(n_0_218), .ZN(n_0_250));
   OAI221_X1 i_0_507 (.A(n_0_250), .B1(n_0_248), .B2(n_0_95), .C1(n_0_249), 
      .C2(n_0_92), .ZN(n_367));
   NOR3_X1 i_0_508 (.A1(n_35), .A2(n_36), .A3(n_0_219), .ZN(n_0_251));
   INV_X1 i_0_541 (.A(n_36), .ZN(n_0_268));
   NAND2_X1 i_0_542 (.A1(n_35), .A2(n_36), .ZN(n_0_274));
   INV_X1 i_0_553 (.A(n_0_274), .ZN(n_0_275));
   NAND2_X1 i_0_555 (.A1(n_0_275), .A2(n_0_219), .ZN(n_0_276));
   INV_X1 i_0_556 (.A(n_0_276), .ZN(n_0_278));
   OAI21_X1 i_0_558 (.A(n_0_274), .B1(n_35), .B2(n_36), .ZN(n_0_279));
   NOR2_X1 i_0_559 (.A1(n_0_279), .A2(n_0_219), .ZN(n_0_280));
   INV_X1 i_0_560 (.A(n_0_280), .ZN(n_0_281));
   OR2_X1 i_0_562 (.A1(n_0_279), .A2(n_34), .ZN(n_0_282));
   OAI21_X1 i_0_564 (.A(n_22), .B1(n_0_278), .B2(n_0_251), .ZN(n_0_301));
   OAI221_X1 i_0_565 (.A(n_0_301), .B1(n_0_282), .B2(n_0_95), .C1(n_0_281), 
      .C2(n_0_92), .ZN(n_368));
   OAI221_X1 i_0_602 (.A(n_0_304), .B1(n_0_305), .B2(n_0_281), .C1(n_0_306), 
      .C2(n_0_282), .ZN(n_369));
   AOI22_X1 i_0_603 (.A1(A_imm_2s_complement[13]), .A2(n_0_251), .B1(n_0_278), 
      .B2(n_9), .ZN(n_0_304));
   INV_X1 i_0_608 (.A(A_imm_2s_complement[14]), .ZN(n_0_305));
   INV_X1 i_0_609 (.A(n_8), .ZN(n_0_306));
   OAI221_X1 i_0_610 (.A(n_0_307), .B1(n_0_310), .B2(n_0_282), .C1(n_0_309), 
      .C2(n_0_276), .ZN(n_370));
   AOI22_X1 i_0_612 (.A1(A_imm_2s_complement[18]), .A2(n_0_280), .B1(
      A_imm_2s_complement[17]), .B2(n_0_251), .ZN(n_0_307));
   INV_X1 i_0_613 (.A(n_5), .ZN(n_0_309));
   INV_X1 i_0_615 (.A(n_4), .ZN(n_0_310));
   NOR3_X1 i_0_616 (.A1(n_37), .A2(n_38), .A3(n_0_268), .ZN(n_0_311));
   INV_X1 i_0_617 (.A(n_38), .ZN(n_0_312));
   NAND2_X1 i_0_619 (.A1(n_37), .A2(n_38), .ZN(n_0_313));
   INV_X1 i_0_621 (.A(n_0_313), .ZN(n_0_330));
   NAND2_X1 i_0_622 (.A1(n_0_330), .A2(n_0_268), .ZN(n_0_334));
   INV_X1 i_0_655 (.A(n_0_334), .ZN(n_0_336));
   OAI21_X1 i_0_656 (.A(n_0_313), .B1(n_37), .B2(n_38), .ZN(n_0_337));
   OR2_X1 i_0_663 (.A1(n_0_337), .A2(n_36), .ZN(n_0_338));
   OR2_X1 i_0_664 (.A1(n_0_337), .A2(n_0_268), .ZN(n_0_340));
   OAI21_X1 i_0_667 (.A(n_22), .B1(n_0_336), .B2(n_0_311), .ZN(n_0_341));
   OAI221_X1 i_0_669 (.A(n_0_341), .B1(n_0_338), .B2(n_0_95), .C1(n_0_340), 
      .C2(n_0_92), .ZN(n_371));
   NOR3_X1 i_0_670 (.A1(n_39), .A2(n_40), .A3(n_0_312), .ZN(n_0_342));
   INV_X1 i_0_672 (.A(n_40), .ZN(n_0_343));
   NAND2_X1 i_0_673 (.A1(n_39), .A2(n_40), .ZN(n_0_345));
   INV_X1 i_0_674 (.A(n_0_345), .ZN(n_0_358));
   NAND2_X1 i_0_676 (.A1(n_0_358), .A2(n_0_312), .ZN(n_0_362));
   INV_X1 i_0_677 (.A(n_0_362), .ZN(n_0_364));
   OAI21_X1 i_0_678 (.A(n_0_345), .B1(n_39), .B2(n_40), .ZN(n_0_366));
   NOR2_X1 i_0_679 (.A1(n_0_366), .A2(n_0_312), .ZN(n_0_367));
   INV_X1 i_0_691 (.A(n_0_367), .ZN(n_0_368));
   OR2_X1 i_0_695 (.A1(n_0_366), .A2(n_38), .ZN(n_0_381));
   OAI21_X1 i_0_697 (.A(n_22), .B1(n_0_364), .B2(n_0_342), .ZN(n_0_387));
   OAI221_X1 i_0_699 (.A(n_0_387), .B1(n_0_381), .B2(n_0_95), .C1(n_0_368), 
      .C2(n_0_92), .ZN(n_372));
   OAI221_X1 i_0_700 (.A(n_0_389), .B1(n_0_381), .B2(n_0_310), .C1(n_0_362), 
      .C2(n_0_309), .ZN(n_373));
   AOI22_X1 i_0_701 (.A1(A_imm_2s_complement[18]), .A2(n_0_367), .B1(
      A_imm_2s_complement[17]), .B2(n_0_342), .ZN(n_0_389));
   NOR3_X1 i_0_702 (.A1(n_41), .A2(n_42), .A3(n_0_343), .ZN(n_0_390));
   INV_X1 i_0_714 (.A(n_42), .ZN(n_0_392));
   NAND2_X1 i_0_718 (.A1(n_41), .A2(n_42), .ZN(n_0_393));
   INV_X1 i_0_720 (.A(n_0_393), .ZN(n_0_394));
   NAND2_X1 i_0_722 (.A1(n_0_394), .A2(n_0_343), .ZN(n_0_395));
   INV_X1 i_0_723 (.A(n_0_395), .ZN(n_0_396));
   OAI21_X1 i_0_724 (.A(n_0_393), .B1(n_41), .B2(n_42), .ZN(n_0_397));
   NOR2_X1 i_0_725 (.A1(n_0_397), .A2(n_0_343), .ZN(n_0_398));
   INV_X1 i_0_726 (.A(n_0_398), .ZN(n_0_399));
   OR2_X1 i_0_727 (.A1(n_0_397), .A2(n_40), .ZN(n_0_400));
   OAI21_X1 i_0_728 (.A(n_22), .B1(n_0_396), .B2(n_0_390), .ZN(n_0_401));
   OAI221_X1 i_0_729 (.A(n_0_401), .B1(n_0_400), .B2(n_0_95), .C1(n_0_399), 
      .C2(n_0_92), .ZN(n_374));
   OAI221_X1 i_0_730 (.A(n_0_402), .B1(n_0_403), .B2(n_0_399), .C1(n_0_404), 
      .C2(n_0_400), .ZN(n_375));
   AOI22_X1 i_0_731 (.A1(A_imm_2s_complement[19]), .A2(n_0_390), .B1(n_0_396), 
      .B2(n_3), .ZN(n_0_402));
   INV_X1 i_0_732 (.A(A_imm_2s_complement[20]), .ZN(n_0_403));
   INV_X1 i_0_733 (.A(n_2), .ZN(n_0_404));
   OAI221_X1 i_0_734 (.A(n_0_405), .B1(n_0_400), .B2(n_0_28), .C1(n_0_395), 
      .C2(n_0_31), .ZN(n_376));
   AOI22_X1 i_0_735 (.A1(A_imm_2s_complement[23]), .A2(n_0_398), .B1(
      A_imm_2s_complement[22]), .B2(n_0_390), .ZN(n_0_405));
   NOR3_X1 i_0_736 (.A1(n_43), .A2(n_44), .A3(n_0_392), .ZN(n_0_406));
   INV_X1 i_0_737 (.A(n_44), .ZN(n_0_407));
   NAND2_X1 i_0_738 (.A1(n_43), .A2(n_44), .ZN(n_0_408));
   INV_X1 i_0_739 (.A(n_0_408), .ZN(n_0_409));
   NAND2_X1 i_0_740 (.A1(n_0_409), .A2(n_0_392), .ZN(n_0_410));
   INV_X1 i_0_741 (.A(n_0_410), .ZN(n_0_411));
   OAI21_X1 i_0_742 (.A(n_0_408), .B1(n_43), .B2(n_44), .ZN(n_0_412));
   NOR2_X1 i_0_743 (.A1(n_0_412), .A2(n_0_392), .ZN(n_0_413));
   INV_X1 i_0_744 (.A(n_0_413), .ZN(n_0_414));
   OR2_X1 i_0_745 (.A1(n_0_412), .A2(n_42), .ZN(n_0_415));
   OAI21_X1 i_0_746 (.A(n_22), .B1(n_0_411), .B2(n_0_406), .ZN(n_0_416));
   OAI221_X1 i_0_747 (.A(n_0_416), .B1(n_0_415), .B2(n_0_95), .C1(n_0_414), 
      .C2(n_0_92), .ZN(n_377));
   OAI221_X1 i_0_748 (.A(n_0_417), .B1(n_0_415), .B2(n_0_310), .C1(n_0_410), 
      .C2(n_0_309), .ZN(n_378));
   AOI22_X1 i_0_749 (.A1(A_imm_2s_complement[18]), .A2(n_0_413), .B1(
      A_imm_2s_complement[17]), .B2(n_0_406), .ZN(n_0_417));
   OAI221_X1 i_0_750 (.A(n_0_418), .B1(n_0_27), .B2(n_0_414), .C1(n_0_415), 
      .C2(n_0_31), .ZN(n_379));
   AOI22_X1 i_0_751 (.A1(A_imm_2s_complement[21]), .A2(n_0_406), .B1(n_0_411), 
      .B2(n_1), .ZN(n_0_418));
   AND2_X1 i_1_0 (.A1(n_1_0__1), .A2(\aggregated_res[14] [23]), .ZN(n_380));
   AND2_X1 i_1_1 (.A1(n_1_0__1), .A2(\aggregated_res[14] [24]), .ZN(n_381));
   AND2_X1 i_1_2 (.A1(n_1_0__1), .A2(\aggregated_res[14] [25]), .ZN(n_382));
   AND2_X1 i_1_3 (.A1(n_1_0__1), .A2(\aggregated_res[14] [26]), .ZN(n_383));
   AND2_X1 i_1_4 (.A1(n_1_0__1), .A2(\aggregated_res[14] [27]), .ZN(n_384));
   AND2_X1 i_1_5 (.A1(n_1_0__1), .A2(\aggregated_res[14] [28]), .ZN(n_385));
   AND2_X1 i_1_6 (.A1(n_1_0__1), .A2(\aggregated_res[14] [29]), .ZN(n_386));
   AND2_X1 i_1_7 (.A1(n_1_0__1), .A2(\aggregated_res[14] [30]), .ZN(n_387));
   AND2_X1 i_1_8 (.A1(n_1_0__1), .A2(\aggregated_res[14] [31]), .ZN(n_388));
   AND2_X1 i_1_9 (.A1(n_1_0__1), .A2(\aggregated_res[14] [32]), .ZN(n_389));
   AND2_X1 i_1_10 (.A1(n_1_0__1), .A2(\aggregated_res[14] [33]), .ZN(n_390));
   AND2_X1 i_1_11 (.A1(n_1_0__1), .A2(\aggregated_res[14] [34]), .ZN(n_391));
   AND2_X1 i_1_12 (.A1(n_1_0__1), .A2(\aggregated_res[14] [35]), .ZN(n_392));
   AND2_X1 i_1_13 (.A1(n_1_0__1), .A2(\aggregated_res[14] [36]), .ZN(n_393));
   AND2_X1 i_1_14 (.A1(n_1_0__1), .A2(\aggregated_res[14] [37]), .ZN(n_394));
   AND2_X1 i_1_15 (.A1(n_1_0__1), .A2(\aggregated_res[14] [38]), .ZN(n_395));
   AND2_X1 i_1_16 (.A1(n_1_0__1), .A2(\aggregated_res[14] [39]), .ZN(n_396));
   AND2_X1 i_1_17 (.A1(n_1_0__1), .A2(\aggregated_res[14] [40]), .ZN(n_397));
   AND2_X1 i_1_18 (.A1(n_1_0__1), .A2(\aggregated_res[14] [41]), .ZN(n_398));
   AND2_X1 i_1_19 (.A1(n_1_0__1), .A2(\aggregated_res[14] [42]), .ZN(n_399));
   AND2_X1 i_1_20 (.A1(n_1_0__1), .A2(\aggregated_res[14] [43]), .ZN(n_400));
   AND2_X1 i_1_21 (.A1(n_1_0__1), .A2(\aggregated_res[14] [44]), .ZN(n_401));
   AND2_X1 i_1_22 (.A1(n_1_0__1), .A2(\aggregated_res[14] [45]), .ZN(n_402));
   AND2_X1 i_1_23 (.A1(n_1_0__1), .A2(\aggregated_res[14] [46]), .ZN(n_403));
   AND2_X1 i_1_24 (.A1(n_1_0__1), .A2(\aggregated_res[14] [47]), .ZN(n_404));
   AND2_X1 i_1_25 (.A1(n_1_0__1), .A2(B[0]), .ZN(n_405));
   AND2_X1 i_1_26 (.A1(n_1_0__1), .A2(B[1]), .ZN(n_406));
   AND2_X1 i_1_27 (.A1(n_1_0__1), .A2(B[2]), .ZN(n_407));
   AND2_X1 i_1_28 (.A1(n_1_0__1), .A2(B[3]), .ZN(n_408));
   AND2_X1 i_1_29 (.A1(n_1_0__1), .A2(B[4]), .ZN(n_409));
   AND2_X1 i_1_30 (.A1(n_1_0__1), .A2(B[5]), .ZN(n_410));
   AND2_X1 i_1_31 (.A1(n_1_0__1), .A2(B[6]), .ZN(n_411));
   AND2_X1 i_1_32 (.A1(n_1_0__1), .A2(B[7]), .ZN(n_412));
   AND2_X1 i_1_33 (.A1(n_1_0__1), .A2(B[8]), .ZN(n_413));
   AND2_X1 i_1_34 (.A1(n_1_0__1), .A2(B[9]), .ZN(n_414));
   AND2_X1 i_1_35 (.A1(n_1_0__1), .A2(B[10]), .ZN(n_415));
   AND2_X1 i_1_36 (.A1(n_1_0__1), .A2(B[11]), .ZN(n_416));
   AND2_X1 i_1_37 (.A1(n_1_0__1), .A2(B[12]), .ZN(n_417));
   AND2_X1 i_1_38 (.A1(n_1_0__1), .A2(B[13]), .ZN(n_418));
   AND2_X1 i_1_39 (.A1(n_1_0__1), .A2(B[14]), .ZN(n_419));
   AND2_X1 i_1_40 (.A1(n_1_0__1), .A2(B[15]), .ZN(n_420));
   AND2_X1 i_1_41 (.A1(n_1_0__1), .A2(B[16]), .ZN(n_421));
   AND2_X1 i_1_42 (.A1(n_1_0__1), .A2(B[17]), .ZN(n_422));
   AND2_X1 i_1_43 (.A1(n_1_0__1), .A2(B[18]), .ZN(n_423));
   AND2_X1 i_1_44 (.A1(n_1_0__1), .A2(B[19]), .ZN(n_424));
   AND2_X1 i_1_45 (.A1(n_1_0__1), .A2(B[20]), .ZN(n_425));
   AND2_X1 i_1_46 (.A1(n_1_0__1), .A2(B[21]), .ZN(n_426));
   AND2_X1 i_1_47 (.A1(n_1_0__1), .A2(B[22]), .ZN(n_427));
   INV_X1 i_1_48 (.A(n_1_0__0), .ZN(n_428));
   AOI21_X1 i_1_49 (.A(reset), .B1(clk), .B2(enable), .ZN(n_1_0__0));
   AND2_X1 i_1_50 (.A1(n_1_0__1), .A2(A[0]), .ZN(n_429));
   AND2_X1 i_1_51 (.A1(n_1_0__1), .A2(A[1]), .ZN(n_430));
   AND2_X1 i_1_52 (.A1(n_1_0__1), .A2(A[2]), .ZN(n_431));
   AND2_X1 i_1_53 (.A1(n_1_0__1), .A2(A[3]), .ZN(n_432));
   AND2_X1 i_1_54 (.A1(n_1_0__1), .A2(A[4]), .ZN(n_433));
   AND2_X1 i_1_55 (.A1(n_1_0__1), .A2(A[5]), .ZN(n_434));
   AND2_X1 i_1_56 (.A1(n_1_0__1), .A2(A[6]), .ZN(n_435));
   AND2_X1 i_1_57 (.A1(n_1_0__1), .A2(A[7]), .ZN(n_436));
   AND2_X1 i_1_58 (.A1(n_1_0__1), .A2(A[8]), .ZN(n_437));
   AND2_X1 i_1_59 (.A1(n_1_0__1), .A2(A[9]), .ZN(n_438));
   AND2_X1 i_1_60 (.A1(n_1_0__1), .A2(A[10]), .ZN(n_439));
   AND2_X1 i_1_61 (.A1(n_1_0__1), .A2(A[11]), .ZN(n_440));
   AND2_X1 i_1_62 (.A1(n_1_0__1), .A2(A[12]), .ZN(n_441));
   AND2_X1 i_1_63 (.A1(n_1_0__1), .A2(A[13]), .ZN(n_442));
   AND2_X1 i_1_64 (.A1(n_1_0__1), .A2(A[14]), .ZN(n_443));
   AND2_X1 i_1_65 (.A1(n_1_0__1), .A2(A[15]), .ZN(n_444));
   AND2_X1 i_1_66 (.A1(n_1_0__1), .A2(A[16]), .ZN(n_445));
   AND2_X1 i_1_67 (.A1(n_1_0__1), .A2(A[17]), .ZN(n_446));
   AND2_X1 i_1_68 (.A1(n_1_0__1), .A2(A[18]), .ZN(n_447));
   AND2_X1 i_1_69 (.A1(n_1_0__1), .A2(A[19]), .ZN(n_448));
   AND2_X1 i_1_70 (.A1(n_1_0__1), .A2(A[20]), .ZN(n_449));
   AND2_X1 i_1_71 (.A1(n_1_0__1), .A2(A[21]), .ZN(n_450));
   AND2_X1 i_1_72 (.A1(n_1_0__1), .A2(A[22]), .ZN(n_451));
   NAND2_X1 i_1_73 (.A1(n_1_0__1), .A2(clk), .ZN(n_452));
   INV_X1 i_1_74 (.A(reset), .ZN(n_1_0__1));
endmodule

module datapath__0_78(M_multiplied, p_0, M_resultTruncated);
   input M_multiplied;
   input [22:0]p_0;
   output [22:0]M_resultTruncated;

   HA_X1 i_0 (.A(M_multiplied), .B(p_0[0]), .CO(n_0), .S(M_resultTruncated[0]));
   HA_X1 i_1 (.A(p_0[1]), .B(n_0), .CO(n_1), .S(M_resultTruncated[1]));
   HA_X1 i_2 (.A(p_0[2]), .B(n_1), .CO(n_2), .S(M_resultTruncated[2]));
   HA_X1 i_3 (.A(p_0[3]), .B(n_2), .CO(n_3), .S(M_resultTruncated[3]));
   HA_X1 i_4 (.A(p_0[4]), .B(n_3), .CO(n_4), .S(M_resultTruncated[4]));
   HA_X1 i_5 (.A(p_0[5]), .B(n_4), .CO(n_5), .S(M_resultTruncated[5]));
   HA_X1 i_6 (.A(p_0[6]), .B(n_5), .CO(n_6), .S(M_resultTruncated[6]));
   HA_X1 i_7 (.A(p_0[7]), .B(n_6), .CO(n_7), .S(M_resultTruncated[7]));
   HA_X1 i_8 (.A(p_0[8]), .B(n_7), .CO(n_8), .S(M_resultTruncated[8]));
   HA_X1 i_9 (.A(p_0[9]), .B(n_8), .CO(n_9), .S(M_resultTruncated[9]));
   HA_X1 i_10 (.A(p_0[10]), .B(n_9), .CO(n_10), .S(M_resultTruncated[10]));
   HA_X1 i_11 (.A(p_0[11]), .B(n_10), .CO(n_11), .S(M_resultTruncated[11]));
   HA_X1 i_12 (.A(p_0[12]), .B(n_11), .CO(n_12), .S(M_resultTruncated[12]));
   HA_X1 i_13 (.A(p_0[13]), .B(n_12), .CO(n_13), .S(M_resultTruncated[13]));
   HA_X1 i_14 (.A(p_0[14]), .B(n_13), .CO(n_14), .S(M_resultTruncated[14]));
   HA_X1 i_15 (.A(p_0[15]), .B(n_14), .CO(n_15), .S(M_resultTruncated[15]));
   HA_X1 i_16 (.A(p_0[16]), .B(n_15), .CO(n_16), .S(M_resultTruncated[16]));
   HA_X1 i_17 (.A(p_0[17]), .B(n_16), .CO(n_17), .S(M_resultTruncated[17]));
   HA_X1 i_18 (.A(p_0[18]), .B(n_17), .CO(n_18), .S(M_resultTruncated[18]));
   HA_X1 i_19 (.A(p_0[19]), .B(n_18), .CO(n_19), .S(M_resultTruncated[19]));
   HA_X1 i_20 (.A(p_0[20]), .B(n_19), .CO(n_20), .S(M_resultTruncated[20]));
   HA_X1 i_21 (.A(p_0[21]), .B(n_20), .CO(n_21), .S(M_resultTruncated[21]));
   XOR2_X1 i_22 (.A(p_0[22]), .B(n_21), .Z(M_resultTruncated[22]));
endmodule

module FPU_boothAlgoR4(Res, A, B, clk, reset, enable);
   output [31:0]Res;
   input [31:0]A;
   input [31:0]B;
   input clk;
   input reset;
   input enable;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire [22:0]M_resultTruncated;
   wire [7:0]EA;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire [7:0]EB;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire A_reg;
   wire B_reg;
   wire n_0_1_2;
   wire n_0_1_3;
   wire n_0_1_4;
   wire n_0_1_5;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_1_8;
   wire n_0_1_9;
   wire n_0_1_10;
   wire n_0_1_11;
   wire n_0_1_12;
   wire n_0_1_13;
   wire n_0_1_14;
   wire n_0_1_15;
   wire n_0_1_22;
   wire n_0_1_16;
   wire n_0_1_23;
   wire n_0_1_17;
   wire n_0_1_24;
   wire n_0_1_18;
   wire n_0_1_25;
   wire n_0_1_19;
   wire n_0_1_26;
   wire n_0_1_20;
   wire n_0_1_27;
   wire n_0_1_21;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_72;
   wire n_0_1_32;
   wire n_0_73;
   wire n_0_1_33;
   wire n_0_74;
   wire n_0_1_34;
   wire n_0_75;
   wire n_0_1_35;
   wire n_0_76;
   wire n_0_1_36;
   wire n_0_77;
   wire n_0_1_37;
   wire n_0_78;
   wire n_0_1_38;
   wire n_0_79;
   wire n_0_1_39;
   wire n_0_80;
   wire n_0_1_40;
   wire n_0_81;
   wire n_0_1_41;
   wire n_0_82;
   wire n_0_1_42;
   wire n_0_83;
   wire n_0_1_43;
   wire n_0_84;
   wire n_0_1_44;
   wire n_0_85;
   wire n_0_1_45;
   wire n_0_86;
   wire n_0_1_46;
   wire n_0_87;
   wire n_0_1_47;
   wire n_0_88;
   wire n_0_1_48;
   wire n_0_89;
   wire n_0_1_49;
   wire n_0_90;
   wire n_0_1_50;
   wire n_0_91;
   wire n_0_1_51;
   wire n_0_92;
   wire n_0_1_52;
   wire n_0_93;
   wire n_0_1_53;
   wire n_0_1_54;
   wire n_0_1_55;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_1_56;
   wire n_0_1_57;
   wire n_0_1_58;
   wire n_0_1_59;
   wire n_0_1_60;
   wire n_0_1_62;
   wire n_0_1_64;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_1_105;
   wire n_0_1_106;
   wire n_0_1_107;
   wire n_0_1_108;
   wire n_0_1_109;
   wire n_0_1_110;
   wire n_0_1_111;
   wire n_0_1_112;
   wire n_0_1_28;
   wire n_0_1_29;
   wire n_0_71;
   wire n_0_1_30;
   wire n_0_1_31;
   wire n_0_1_61;
   wire n_0_1_63;
   wire n_0_1_65;
   wire n_0_1_66;
   wire n_0_1_67;
   wire n_0_1_68;
   wire n_0_1_69;
   wire n_0_1_70;
   wire n_0_1_71;
   wire n_0_1_72;
   wire n_0_1_73;
   wire n_0_1_74;
   wire n_0_1_75;
   wire n_0_1_76;
   wire n_0_1_77;
   wire n_0_1_78;
   wire n_0_1_79;
   wire n_0_1_80;
   wire n_0_1_81;
   wire n_0_1_82;
   wire n_0_1_83;
   wire n_0_1_84;
   wire n_0_1_85;
   wire n_0_1_86;
   wire n_0_1_87;
   wire n_0_1_88;
   wire n_0_1_89;
   wire n_0_1_90;
   wire n_0_1_91;
   wire n_0_1_92;
   wire n_0_1_93;
   wire n_0_1_94;
   wire n_0_1_95;
   wire n_0_1_96;
   wire n_0_1_97;
   wire n_0_1_98;
   wire n_0_1_99;
   wire n_0_1_100;
   wire n_0_1_101;
   wire n_0_1_102;
   wire n_0_1_103;
   wire n_0_102;
   wire n_0_1_104;

   boothAlgoR4 multiplier (.Res({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, 
      uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, n_0_24, n_0_23, 
      n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, 
      n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, 
      n_0_3, n_0_2, n_0_1, n_0_0, uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, 
      uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, 
      uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, uc_38}), .OVF(), .A({uc_39, 
      uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, n_0_25, n_0_26, 
      n_0_27, n_0_28, n_0_29, n_0_30, n_0_31, n_0_32, n_0_33, n_0_34, n_0_35, 
      n_0_36, n_0_37, n_0_38, n_0_39, n_0_40, n_0_41, n_0_42, n_0_43, n_0_44, 
      n_0_45, n_0_46, n_0_47}), .B({uc_48, uc_49, uc_50, uc_51, uc_52, uc_53, 
      uc_54, uc_55, uc_56, n_0_48, n_0_49, n_0_50, n_0_51, n_0_52, n_0_53, 
      n_0_54, n_0_55, n_0_56, n_0_57, n_0_58, n_0_59, n_0_60, n_0_61, n_0_62, 
      n_0_63, n_0_64, n_0_65, n_0_66, n_0_67, n_0_68, n_0_69, n_0_70}), .clk(clk), 
      .reset(reset), .enable(enable));
   datapath__0_78 i_0_0 (.M_multiplied(n_0_0), .p_0({n_0_23, n_0_22, n_0_21, 
      n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, 
      n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, 
      n_0_1}), .M_resultTruncated(M_resultTruncated));
   DLH_X1 \Res_reg[31]  (.D(n_0_102), .G(n_0_168), .Q(Res[31]));
   DLH_X1 \Res_reg[30]  (.D(n_0_101), .G(n_0_168), .Q(Res[30]));
   DLH_X1 \Res_reg[29]  (.D(n_0_100), .G(n_0_168), .Q(Res[29]));
   DLH_X1 \Res_reg[28]  (.D(n_0_99), .G(n_0_168), .Q(Res[28]));
   DLH_X1 \Res_reg[27]  (.D(n_0_98), .G(n_0_168), .Q(Res[27]));
   DLH_X1 \Res_reg[26]  (.D(n_0_97), .G(n_0_168), .Q(Res[26]));
   DLH_X1 \Res_reg[25]  (.D(n_0_96), .G(n_0_168), .Q(Res[25]));
   DLH_X1 \Res_reg[24]  (.D(n_0_95), .G(n_0_168), .Q(Res[24]));
   DLH_X1 \Res_reg[23]  (.D(n_0_94), .G(n_0_168), .Q(Res[23]));
   DLH_X1 \Res_reg[22]  (.D(n_0_93), .G(n_0_168), .Q(Res[22]));
   DLH_X1 \Res_reg[21]  (.D(n_0_92), .G(n_0_168), .Q(Res[21]));
   DLH_X1 \Res_reg[20]  (.D(n_0_91), .G(n_0_168), .Q(Res[20]));
   DLH_X1 \Res_reg[19]  (.D(n_0_90), .G(n_0_168), .Q(Res[19]));
   DLH_X1 \Res_reg[18]  (.D(n_0_89), .G(n_0_168), .Q(Res[18]));
   DLH_X1 \Res_reg[17]  (.D(n_0_88), .G(n_0_168), .Q(Res[17]));
   DLH_X1 \Res_reg[16]  (.D(n_0_87), .G(n_0_168), .Q(Res[16]));
   DLH_X1 \Res_reg[15]  (.D(n_0_86), .G(n_0_168), .Q(Res[15]));
   DLH_X1 \Res_reg[14]  (.D(n_0_85), .G(n_0_168), .Q(Res[14]));
   DLH_X1 \Res_reg[13]  (.D(n_0_84), .G(n_0_168), .Q(Res[13]));
   DLH_X1 \Res_reg[12]  (.D(n_0_83), .G(n_0_168), .Q(Res[12]));
   DLH_X1 \Res_reg[11]  (.D(n_0_82), .G(n_0_168), .Q(Res[11]));
   DLH_X1 \Res_reg[10]  (.D(n_0_81), .G(n_0_168), .Q(Res[10]));
   DLH_X1 \Res_reg[9]  (.D(n_0_80), .G(n_0_168), .Q(Res[9]));
   DLH_X1 \Res_reg[8]  (.D(n_0_79), .G(n_0_168), .Q(Res[8]));
   DLH_X1 \Res_reg[7]  (.D(n_0_78), .G(n_0_168), .Q(Res[7]));
   DLH_X1 \Res_reg[6]  (.D(n_0_77), .G(n_0_168), .Q(Res[6]));
   DLH_X1 \Res_reg[5]  (.D(n_0_76), .G(n_0_168), .Q(Res[5]));
   DLH_X1 \Res_reg[4]  (.D(n_0_75), .G(n_0_168), .Q(Res[4]));
   DLH_X1 \Res_reg[3]  (.D(n_0_74), .G(n_0_168), .Q(Res[3]));
   DLH_X1 \Res_reg[2]  (.D(n_0_73), .G(n_0_168), .Q(Res[2]));
   DLH_X1 \Res_reg[1]  (.D(n_0_72), .G(n_0_168), .Q(Res[1]));
   DLH_X1 \Res_reg[0]  (.D(n_0_71), .G(n_0_168), .Q(Res[0]));
   DLH_X1 \A_reg_reg[30]  (.D(n_0_136), .G(n_0_104), .Q(EA[7]));
   DLH_X1 \A_reg_reg[29]  (.D(n_0_135), .G(n_0_104), .Q(EA[6]));
   DLH_X1 \A_reg_reg[28]  (.D(n_0_134), .G(n_0_104), .Q(EA[5]));
   DLH_X1 \A_reg_reg[27]  (.D(n_0_133), .G(n_0_104), .Q(EA[4]));
   DLH_X1 \A_reg_reg[26]  (.D(n_0_132), .G(n_0_104), .Q(EA[3]));
   DLH_X1 \A_reg_reg[25]  (.D(n_0_131), .G(n_0_104), .Q(EA[2]));
   DLH_X1 \A_reg_reg[24]  (.D(n_0_130), .G(n_0_104), .Q(EA[1]));
   DLH_X1 \A_reg_reg[23]  (.D(n_0_129), .G(n_0_104), .Q(EA[0]));
   DLH_X1 \A_reg_reg[22]  (.D(n_0_128), .G(n_0_104), .Q(n_0_25));
   DLH_X1 \A_reg_reg[21]  (.D(n_0_127), .G(n_0_104), .Q(n_0_26));
   DLH_X1 \A_reg_reg[20]  (.D(n_0_126), .G(n_0_104), .Q(n_0_27));
   DLH_X1 \A_reg_reg[19]  (.D(n_0_125), .G(n_0_104), .Q(n_0_28));
   DLH_X1 \A_reg_reg[18]  (.D(n_0_124), .G(n_0_104), .Q(n_0_29));
   DLH_X1 \A_reg_reg[17]  (.D(n_0_123), .G(n_0_104), .Q(n_0_30));
   DLH_X1 \A_reg_reg[16]  (.D(n_0_122), .G(n_0_104), .Q(n_0_31));
   DLH_X1 \A_reg_reg[15]  (.D(n_0_121), .G(n_0_104), .Q(n_0_32));
   DLH_X1 \A_reg_reg[14]  (.D(n_0_120), .G(n_0_104), .Q(n_0_33));
   DLH_X1 \A_reg_reg[13]  (.D(n_0_119), .G(n_0_104), .Q(n_0_34));
   DLH_X1 \A_reg_reg[12]  (.D(n_0_118), .G(n_0_104), .Q(n_0_35));
   DLH_X1 \A_reg_reg[11]  (.D(n_0_117), .G(n_0_104), .Q(n_0_36));
   DLH_X1 \A_reg_reg[10]  (.D(n_0_116), .G(n_0_104), .Q(n_0_37));
   DLH_X1 \A_reg_reg[9]  (.D(n_0_115), .G(n_0_104), .Q(n_0_38));
   DLH_X1 \A_reg_reg[8]  (.D(n_0_114), .G(n_0_104), .Q(n_0_39));
   DLH_X1 \A_reg_reg[7]  (.D(n_0_113), .G(n_0_104), .Q(n_0_40));
   DLH_X1 \A_reg_reg[6]  (.D(n_0_112), .G(n_0_104), .Q(n_0_41));
   DLH_X1 \A_reg_reg[5]  (.D(n_0_111), .G(n_0_104), .Q(n_0_42));
   DLH_X1 \A_reg_reg[4]  (.D(n_0_110), .G(n_0_104), .Q(n_0_43));
   DLH_X1 \A_reg_reg[3]  (.D(n_0_109), .G(n_0_104), .Q(n_0_44));
   DLH_X1 \A_reg_reg[2]  (.D(n_0_108), .G(n_0_104), .Q(n_0_45));
   DLH_X1 \A_reg_reg[1]  (.D(n_0_107), .G(n_0_104), .Q(n_0_46));
   DLH_X1 \A_reg_reg[0]  (.D(n_0_106), .G(n_0_104), .Q(n_0_47));
   DLH_X1 \B_reg_reg[30]  (.D(n_0_167), .G(n_0_104), .Q(EB[7]));
   DLH_X1 \B_reg_reg[29]  (.D(n_0_166), .G(n_0_104), .Q(EB[6]));
   DLH_X1 \B_reg_reg[28]  (.D(n_0_165), .G(n_0_104), .Q(EB[5]));
   DLH_X1 \B_reg_reg[27]  (.D(n_0_164), .G(n_0_104), .Q(EB[4]));
   DLH_X1 \B_reg_reg[26]  (.D(n_0_163), .G(n_0_104), .Q(EB[3]));
   DLH_X1 \B_reg_reg[25]  (.D(n_0_162), .G(n_0_104), .Q(EB[2]));
   DLH_X1 \B_reg_reg[24]  (.D(n_0_161), .G(n_0_104), .Q(EB[1]));
   DLH_X1 \B_reg_reg[23]  (.D(n_0_160), .G(n_0_104), .Q(EB[0]));
   DLH_X1 \B_reg_reg[22]  (.D(n_0_159), .G(n_0_104), .Q(n_0_48));
   DLH_X1 \B_reg_reg[21]  (.D(n_0_158), .G(n_0_104), .Q(n_0_49));
   DLH_X1 \B_reg_reg[20]  (.D(n_0_157), .G(n_0_104), .Q(n_0_50));
   DLH_X1 \B_reg_reg[19]  (.D(n_0_156), .G(n_0_104), .Q(n_0_51));
   DLH_X1 \B_reg_reg[18]  (.D(n_0_155), .G(n_0_104), .Q(n_0_52));
   DLH_X1 \B_reg_reg[17]  (.D(n_0_154), .G(n_0_104), .Q(n_0_53));
   DLH_X1 \B_reg_reg[16]  (.D(n_0_153), .G(n_0_104), .Q(n_0_54));
   DLH_X1 \B_reg_reg[15]  (.D(n_0_152), .G(n_0_104), .Q(n_0_55));
   DLH_X1 \B_reg_reg[14]  (.D(n_0_151), .G(n_0_104), .Q(n_0_56));
   DLH_X1 \B_reg_reg[13]  (.D(n_0_150), .G(n_0_104), .Q(n_0_57));
   DLH_X1 \B_reg_reg[12]  (.D(n_0_149), .G(n_0_104), .Q(n_0_58));
   DLH_X1 \B_reg_reg[11]  (.D(n_0_148), .G(n_0_104), .Q(n_0_59));
   DLH_X1 \B_reg_reg[10]  (.D(n_0_147), .G(n_0_104), .Q(n_0_60));
   DLH_X1 \B_reg_reg[9]  (.D(n_0_146), .G(n_0_104), .Q(n_0_61));
   DLH_X1 \B_reg_reg[8]  (.D(n_0_145), .G(n_0_104), .Q(n_0_62));
   DLH_X1 \B_reg_reg[7]  (.D(n_0_144), .G(n_0_104), .Q(n_0_63));
   DLH_X1 \B_reg_reg[6]  (.D(n_0_143), .G(n_0_104), .Q(n_0_64));
   DLH_X1 \B_reg_reg[5]  (.D(n_0_142), .G(n_0_104), .Q(n_0_65));
   DLH_X1 \B_reg_reg[4]  (.D(n_0_141), .G(n_0_104), .Q(n_0_66));
   DLH_X1 \B_reg_reg[3]  (.D(n_0_140), .G(n_0_104), .Q(n_0_67));
   DLH_X1 \B_reg_reg[2]  (.D(n_0_139), .G(n_0_104), .Q(n_0_68));
   DLH_X1 \B_reg_reg[1]  (.D(n_0_138), .G(n_0_104), .Q(n_0_69));
   DLH_X1 \B_reg_reg[0]  (.D(n_0_137), .G(n_0_104), .Q(n_0_70));
   DLH_X1 \A_reg_reg[31]  (.D(n_0_103), .G(n_0_104), .Q(A_reg));
   DLH_X1 \B_reg_reg[31]  (.D(n_0_105), .G(n_0_104), .Q(B_reg));
   HA_X1 i_0_1_0 (.A(EB[1]), .B(EA[1]), .CO(n_0_1_3), .S(n_0_1_2));
   HA_X1 i_0_1_1 (.A(EB[2]), .B(EA[2]), .CO(n_0_1_5), .S(n_0_1_4));
   HA_X1 i_0_1_2 (.A(EB[3]), .B(EA[3]), .CO(n_0_1_7), .S(n_0_1_6));
   HA_X1 i_0_1_3 (.A(EB[4]), .B(EA[4]), .CO(n_0_1_9), .S(n_0_1_8));
   HA_X1 i_0_1_4 (.A(EB[5]), .B(EA[5]), .CO(n_0_1_11), .S(n_0_1_10));
   HA_X1 i_0_1_5 (.A(EB[6]), .B(EA[6]), .CO(n_0_1_13), .S(n_0_1_12));
   HA_X1 i_0_1_6 (.A(EA[0]), .B(n_0_1_0), .CO(n_0_1_15), .S(n_0_1_14));
   FA_X1 i_0_1_7 (.A(n_0_1_1), .B(n_0_1_2), .CI(n_0_1_15), .CO(n_0_1_16), 
      .S(n_0_1_22));
   FA_X1 i_0_1_8 (.A(n_0_1_3), .B(n_0_1_4), .CI(n_0_1_16), .CO(n_0_1_17), 
      .S(n_0_1_23));
   FA_X1 i_0_1_9 (.A(n_0_1_5), .B(n_0_1_6), .CI(n_0_1_17), .CO(n_0_1_18), 
      .S(n_0_1_24));
   FA_X1 i_0_1_10 (.A(n_0_1_7), .B(n_0_1_8), .CI(n_0_1_18), .CO(n_0_1_19), 
      .S(n_0_1_25));
   FA_X1 i_0_1_11 (.A(n_0_1_9), .B(n_0_1_10), .CI(n_0_1_19), .CO(n_0_1_20), 
      .S(n_0_1_26));
   FA_X1 i_0_1_12 (.A(n_0_1_11), .B(n_0_1_12), .CI(n_0_1_20), .CO(n_0_1_21), 
      .S(n_0_1_27));
   XNOR2_X1 i_0_1_13 (.A(EB[0]), .B(n_0_24), .ZN(n_0_1_0));
   OR2_X1 i_0_1_14 (.A1(EB[0]), .A2(n_0_24), .ZN(n_0_1_1));
   INV_X1 i_0_1_15 (.A(n_0_1_32), .ZN(n_0_72));
   AOI22_X1 i_0_1_16 (.A1(M_resultTruncated[1]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_1), .ZN(n_0_1_32));
   INV_X1 i_0_1_22 (.A(n_0_1_33), .ZN(n_0_73));
   AOI22_X1 i_0_1_23 (.A1(M_resultTruncated[2]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_2), .ZN(n_0_1_33));
   INV_X1 i_0_1_24 (.A(n_0_1_34), .ZN(n_0_74));
   AOI22_X1 i_0_1_25 (.A1(M_resultTruncated[3]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_3), .ZN(n_0_1_34));
   INV_X1 i_0_1_26 (.A(n_0_1_35), .ZN(n_0_75));
   AOI22_X1 i_0_1_27 (.A1(M_resultTruncated[4]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_4), .ZN(n_0_1_35));
   INV_X1 i_0_1_28 (.A(n_0_1_36), .ZN(n_0_76));
   AOI22_X1 i_0_1_29 (.A1(M_resultTruncated[5]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_5), .ZN(n_0_1_36));
   INV_X1 i_0_1_30 (.A(n_0_1_37), .ZN(n_0_77));
   AOI22_X1 i_0_1_31 (.A1(M_resultTruncated[6]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_6), .ZN(n_0_1_37));
   INV_X1 i_0_1_32 (.A(n_0_1_38), .ZN(n_0_78));
   AOI22_X1 i_0_1_33 (.A1(M_resultTruncated[7]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_7), .ZN(n_0_1_38));
   INV_X1 i_0_1_34 (.A(n_0_1_39), .ZN(n_0_79));
   AOI22_X1 i_0_1_35 (.A1(M_resultTruncated[8]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_8), .ZN(n_0_1_39));
   INV_X1 i_0_1_36 (.A(n_0_1_40), .ZN(n_0_80));
   AOI22_X1 i_0_1_37 (.A1(M_resultTruncated[9]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_9), .ZN(n_0_1_40));
   INV_X1 i_0_1_38 (.A(n_0_1_41), .ZN(n_0_81));
   AOI22_X1 i_0_1_39 (.A1(M_resultTruncated[10]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_10), .ZN(n_0_1_41));
   INV_X1 i_0_1_40 (.A(n_0_1_42), .ZN(n_0_82));
   AOI22_X1 i_0_1_41 (.A1(M_resultTruncated[11]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_11), .ZN(n_0_1_42));
   INV_X1 i_0_1_42 (.A(n_0_1_43), .ZN(n_0_83));
   AOI22_X1 i_0_1_43 (.A1(M_resultTruncated[12]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_12), .ZN(n_0_1_43));
   INV_X1 i_0_1_44 (.A(n_0_1_44), .ZN(n_0_84));
   AOI22_X1 i_0_1_45 (.A1(M_resultTruncated[13]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_13), .ZN(n_0_1_44));
   INV_X1 i_0_1_46 (.A(n_0_1_45), .ZN(n_0_85));
   AOI22_X1 i_0_1_47 (.A1(M_resultTruncated[14]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_14), .ZN(n_0_1_45));
   INV_X1 i_0_1_48 (.A(n_0_1_46), .ZN(n_0_86));
   AOI22_X1 i_0_1_49 (.A1(M_resultTruncated[15]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_15), .ZN(n_0_1_46));
   INV_X1 i_0_1_50 (.A(n_0_1_47), .ZN(n_0_87));
   AOI22_X1 i_0_1_51 (.A1(M_resultTruncated[16]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_16), .ZN(n_0_1_47));
   INV_X1 i_0_1_52 (.A(n_0_1_48), .ZN(n_0_88));
   AOI22_X1 i_0_1_53 (.A1(M_resultTruncated[17]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_17), .ZN(n_0_1_48));
   INV_X1 i_0_1_54 (.A(n_0_1_49), .ZN(n_0_89));
   AOI22_X1 i_0_1_55 (.A1(M_resultTruncated[18]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_18), .ZN(n_0_1_49));
   INV_X1 i_0_1_56 (.A(n_0_1_50), .ZN(n_0_90));
   AOI22_X1 i_0_1_57 (.A1(M_resultTruncated[19]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_19), .ZN(n_0_1_50));
   INV_X1 i_0_1_58 (.A(n_0_1_51), .ZN(n_0_91));
   AOI22_X1 i_0_1_59 (.A1(M_resultTruncated[20]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_20), .ZN(n_0_1_51));
   INV_X1 i_0_1_60 (.A(n_0_1_52), .ZN(n_0_92));
   AOI22_X1 i_0_1_61 (.A1(M_resultTruncated[21]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_21), .ZN(n_0_1_52));
   INV_X1 i_0_1_62 (.A(n_0_1_53), .ZN(n_0_93));
   AOI22_X1 i_0_1_63 (.A1(M_resultTruncated[22]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_22), .ZN(n_0_1_53));
   NOR3_X1 i_0_1_17 (.A1(n_0_1_60), .A2(n_0_24), .A3(n_0_1_64), .ZN(n_0_1_54));
   NOR3_X1 i_0_1_18 (.A1(n_0_1_29), .A2(n_0_1_64), .A3(n_0_1_60), .ZN(n_0_1_55));
   OAI21_X1 i_0_1_19 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_111), .ZN(n_0_94));
   OAI21_X1 i_0_1_67 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_110), .ZN(n_0_95));
   OAI21_X1 i_0_1_68 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_109), .ZN(n_0_96));
   OAI21_X1 i_0_1_69 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_108), .ZN(n_0_97));
   OAI21_X1 i_0_1_70 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_107), .ZN(n_0_98));
   OAI21_X1 i_0_1_71 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_106), .ZN(n_0_99));
   OAI21_X1 i_0_1_72 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_105), .ZN(n_0_100));
   OAI21_X1 i_0_1_73 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_56), .ZN(n_0_101));
   XNOR2_X1 i_0_1_74 (.A(n_0_1_58), .B(n_0_1_57), .ZN(n_0_1_56));
   XNOR2_X1 i_0_1_75 (.A(n_0_1_13), .B(n_0_1_21), .ZN(n_0_1_57));
   NOR2_X1 i_0_1_76 (.A1(n_0_1_68), .A2(n_0_1_59), .ZN(n_0_1_58));
   NOR2_X1 i_0_1_77 (.A1(EB[7]), .A2(EA[7]), .ZN(n_0_1_59));
   NAND2_X1 i_0_1_20 (.A1(n_0_1_69), .A2(n_0_1_66), .ZN(n_0_1_60));
   AOI21_X1 i_0_1_21 (.A(n_0_1_72), .B1(n_0_1_69), .B2(n_0_1_64), .ZN(n_0_1_62));
   NAND3_X1 i_0_1_64 (.A1(n_0_1_100), .A2(n_0_1_97), .A3(n_0_1_67), .ZN(n_0_1_64));
   AND2_X1 i_0_1_65 (.A1(n_0_1_112), .A2(A[31]), .ZN(n_0_103));
   OAI21_X1 i_0_1_125 (.A(n_0_1_112), .B1(n_0_1_28), .B2(clk), .ZN(n_0_104));
   AND2_X1 i_0_1_126 (.A1(n_0_1_112), .A2(B[31]), .ZN(n_0_105));
   AND2_X1 i_0_1_127 (.A1(n_0_1_112), .A2(A[0]), .ZN(n_0_106));
   AND2_X1 i_0_1_128 (.A1(n_0_1_112), .A2(A[1]), .ZN(n_0_107));
   AND2_X1 i_0_1_129 (.A1(n_0_1_112), .A2(A[2]), .ZN(n_0_108));
   AND2_X1 i_0_1_130 (.A1(n_0_1_112), .A2(A[3]), .ZN(n_0_109));
   AND2_X1 i_0_1_131 (.A1(n_0_1_112), .A2(A[4]), .ZN(n_0_110));
   AND2_X1 i_0_1_132 (.A1(n_0_1_112), .A2(A[5]), .ZN(n_0_111));
   AND2_X1 i_0_1_133 (.A1(n_0_1_112), .A2(A[6]), .ZN(n_0_112));
   AND2_X1 i_0_1_134 (.A1(n_0_1_112), .A2(A[7]), .ZN(n_0_113));
   AND2_X1 i_0_1_135 (.A1(n_0_1_112), .A2(A[8]), .ZN(n_0_114));
   AND2_X1 i_0_1_136 (.A1(n_0_1_112), .A2(A[9]), .ZN(n_0_115));
   AND2_X1 i_0_1_137 (.A1(n_0_1_112), .A2(A[10]), .ZN(n_0_116));
   AND2_X1 i_0_1_138 (.A1(n_0_1_112), .A2(A[11]), .ZN(n_0_117));
   AND2_X1 i_0_1_139 (.A1(n_0_1_112), .A2(A[12]), .ZN(n_0_118));
   AND2_X1 i_0_1_140 (.A1(n_0_1_112), .A2(A[13]), .ZN(n_0_119));
   AND2_X1 i_0_1_141 (.A1(n_0_1_112), .A2(A[14]), .ZN(n_0_120));
   AND2_X1 i_0_1_142 (.A1(n_0_1_112), .A2(A[15]), .ZN(n_0_121));
   AND2_X1 i_0_1_143 (.A1(n_0_1_112), .A2(A[16]), .ZN(n_0_122));
   AND2_X1 i_0_1_144 (.A1(n_0_1_112), .A2(A[17]), .ZN(n_0_123));
   AND2_X1 i_0_1_145 (.A1(n_0_1_112), .A2(A[18]), .ZN(n_0_124));
   AND2_X1 i_0_1_146 (.A1(n_0_1_112), .A2(A[19]), .ZN(n_0_125));
   AND2_X1 i_0_1_147 (.A1(n_0_1_112), .A2(A[20]), .ZN(n_0_126));
   AND2_X1 i_0_1_148 (.A1(n_0_1_112), .A2(A[21]), .ZN(n_0_127));
   AND2_X1 i_0_1_149 (.A1(n_0_1_112), .A2(A[22]), .ZN(n_0_128));
   AND2_X1 i_0_1_150 (.A1(n_0_1_112), .A2(A[23]), .ZN(n_0_129));
   AND2_X1 i_0_1_151 (.A1(n_0_1_112), .A2(A[24]), .ZN(n_0_130));
   AND2_X1 i_0_1_152 (.A1(n_0_1_112), .A2(A[25]), .ZN(n_0_131));
   AND2_X1 i_0_1_153 (.A1(n_0_1_112), .A2(A[26]), .ZN(n_0_132));
   AND2_X1 i_0_1_154 (.A1(n_0_1_112), .A2(A[27]), .ZN(n_0_133));
   AND2_X1 i_0_1_155 (.A1(n_0_1_112), .A2(A[28]), .ZN(n_0_134));
   AND2_X1 i_0_1_156 (.A1(n_0_1_112), .A2(A[29]), .ZN(n_0_135));
   AND2_X1 i_0_1_157 (.A1(n_0_1_112), .A2(A[30]), .ZN(n_0_136));
   AND2_X1 i_0_1_158 (.A1(n_0_1_112), .A2(B[0]), .ZN(n_0_137));
   AND2_X1 i_0_1_159 (.A1(n_0_1_112), .A2(B[1]), .ZN(n_0_138));
   AND2_X1 i_0_1_160 (.A1(n_0_1_112), .A2(B[2]), .ZN(n_0_139));
   AND2_X1 i_0_1_161 (.A1(n_0_1_112), .A2(B[3]), .ZN(n_0_140));
   AND2_X1 i_0_1_162 (.A1(n_0_1_112), .A2(B[4]), .ZN(n_0_141));
   AND2_X1 i_0_1_163 (.A1(n_0_1_112), .A2(B[5]), .ZN(n_0_142));
   AND2_X1 i_0_1_164 (.A1(n_0_1_112), .A2(B[6]), .ZN(n_0_143));
   AND2_X1 i_0_1_165 (.A1(n_0_1_112), .A2(B[7]), .ZN(n_0_144));
   AND2_X1 i_0_1_166 (.A1(n_0_1_112), .A2(B[8]), .ZN(n_0_145));
   AND2_X1 i_0_1_167 (.A1(n_0_1_112), .A2(B[9]), .ZN(n_0_146));
   AND2_X1 i_0_1_168 (.A1(n_0_1_112), .A2(B[10]), .ZN(n_0_147));
   AND2_X1 i_0_1_169 (.A1(n_0_1_112), .A2(B[11]), .ZN(n_0_148));
   AND2_X1 i_0_1_170 (.A1(n_0_1_112), .A2(B[12]), .ZN(n_0_149));
   AND2_X1 i_0_1_171 (.A1(n_0_1_112), .A2(B[13]), .ZN(n_0_150));
   AND2_X1 i_0_1_172 (.A1(n_0_1_112), .A2(B[14]), .ZN(n_0_151));
   AND2_X1 i_0_1_173 (.A1(n_0_1_112), .A2(B[15]), .ZN(n_0_152));
   AND2_X1 i_0_1_174 (.A1(n_0_1_112), .A2(B[16]), .ZN(n_0_153));
   AND2_X1 i_0_1_175 (.A1(n_0_1_112), .A2(B[17]), .ZN(n_0_154));
   AND2_X1 i_0_1_176 (.A1(n_0_1_112), .A2(B[18]), .ZN(n_0_155));
   AND2_X1 i_0_1_177 (.A1(n_0_1_112), .A2(B[19]), .ZN(n_0_156));
   AND2_X1 i_0_1_178 (.A1(n_0_1_112), .A2(B[20]), .ZN(n_0_157));
   AND2_X1 i_0_1_179 (.A1(n_0_1_112), .A2(B[21]), .ZN(n_0_158));
   AND2_X1 i_0_1_180 (.A1(n_0_1_112), .A2(B[22]), .ZN(n_0_159));
   AND2_X1 i_0_1_181 (.A1(n_0_1_112), .A2(B[23]), .ZN(n_0_160));
   AND2_X1 i_0_1_182 (.A1(n_0_1_112), .A2(B[24]), .ZN(n_0_161));
   AND2_X1 i_0_1_183 (.A1(n_0_1_112), .A2(B[25]), .ZN(n_0_162));
   AND2_X1 i_0_1_184 (.A1(n_0_1_112), .A2(B[26]), .ZN(n_0_163));
   AND2_X1 i_0_1_185 (.A1(n_0_1_112), .A2(B[27]), .ZN(n_0_164));
   AND2_X1 i_0_1_186 (.A1(n_0_1_112), .A2(B[28]), .ZN(n_0_165));
   AND2_X1 i_0_1_187 (.A1(n_0_1_112), .A2(B[29]), .ZN(n_0_166));
   AND2_X1 i_0_1_188 (.A1(n_0_1_112), .A2(B[30]), .ZN(n_0_167));
   OR2_X1 i_0_1_189 (.A1(clk), .A2(reset), .ZN(n_0_168));
   INV_X1 i_0_1_190 (.A(n_0_1_27), .ZN(n_0_1_105));
   INV_X1 i_0_1_191 (.A(n_0_1_26), .ZN(n_0_1_106));
   INV_X1 i_0_1_192 (.A(n_0_1_25), .ZN(n_0_1_107));
   INV_X1 i_0_1_193 (.A(n_0_1_24), .ZN(n_0_1_108));
   INV_X1 i_0_1_194 (.A(n_0_1_23), .ZN(n_0_1_109));
   INV_X1 i_0_1_195 (.A(n_0_1_22), .ZN(n_0_1_110));
   INV_X1 i_0_1_66 (.A(n_0_1_14), .ZN(n_0_1_111));
   INV_X1 i_0_1_78 (.A(reset), .ZN(n_0_1_112));
   INV_X1 i_0_1_198 (.A(enable), .ZN(n_0_1_28));
   INV_X1 i_0_1_79 (.A(n_0_24), .ZN(n_0_1_29));
   OAI21_X1 i_0_1_80 (.A(n_0_1_71), .B1(n_0_1_31), .B2(n_0_1_30), .ZN(n_0_71));
   OAI221_X1 i_0_1_81 (.A(n_0_1_69), .B1(n_0_1_100), .B2(n_0_1_81), .C1(n_0_1_97), 
      .C2(n_0_1_73), .ZN(n_0_1_30));
   INV_X1 i_0_1_82 (.A(n_0_1_61), .ZN(n_0_1_31));
   OAI211_X1 i_0_1_83 (.A(n_0_1_100), .B(n_0_1_97), .C1(n_0_1_65), .C2(n_0_1_63), 
      .ZN(n_0_1_61));
   NAND2_X1 i_0_1_84 (.A1(n_0_1_67), .A2(n_0_1_66), .ZN(n_0_1_63));
   AOI22_X1 i_0_1_85 (.A1(n_0_1_103), .A2(n_0_0), .B1(n_0_24), .B2(
      M_resultTruncated[0]), .ZN(n_0_1_65));
   OR4_X1 i_0_1_86 (.A1(n_0_1_101), .A2(n_0_1_98), .A3(n_0_1_92), .A4(n_0_1_95), 
      .ZN(n_0_1_66));
   OAI221_X1 i_0_1_87 (.A(n_0_1_68), .B1(EA[6]), .B2(n_0_1_98), .C1(EB[6]), 
      .C2(n_0_1_101), .ZN(n_0_1_67));
   AND2_X1 i_0_1_88 (.A1(EA[7]), .A2(EB[7]), .ZN(n_0_1_68));
   NOR2_X1 i_0_1_89 (.A1(reset), .A2(n_0_1_70), .ZN(n_0_1_69));
   OAI22_X1 i_0_1_90 (.A1(n_0_1_91), .A2(n_0_1_81), .B1(n_0_1_94), .B2(n_0_1_73), 
      .ZN(n_0_1_70));
   INV_X1 i_0_1_91 (.A(n_0_1_72), .ZN(n_0_1_71));
   NOR4_X1 i_0_1_92 (.A1(reset), .A2(n_0_1_73), .A3(n_0_1_81), .A4(n_0_1_89), 
      .ZN(n_0_1_72));
   NAND3_X1 i_0_1_93 (.A1(n_0_1_78), .A2(n_0_1_77), .A3(n_0_1_74), .ZN(n_0_1_73));
   AND4_X1 i_0_1_94 (.A1(n_0_1_80), .A2(n_0_1_79), .A3(n_0_1_76), .A4(n_0_1_75), 
      .ZN(n_0_1_74));
   NOR4_X1 i_0_1_95 (.A1(n_0_45), .A2(n_0_47), .A3(n_0_41), .A4(n_0_44), 
      .ZN(n_0_1_75));
   NOR4_X1 i_0_1_96 (.A1(n_0_37), .A2(n_0_40), .A3(n_0_34), .A4(n_0_35), 
      .ZN(n_0_1_76));
   NOR3_X1 i_0_1_97 (.A1(n_0_42), .A2(n_0_43), .A3(n_0_46), .ZN(n_0_1_77));
   NOR4_X1 i_0_1_98 (.A1(n_0_38), .A2(n_0_39), .A3(n_0_33), .A4(n_0_36), 
      .ZN(n_0_1_78));
   NOR4_X1 i_0_1_99 (.A1(n_0_25), .A2(n_0_26), .A3(n_0_27), .A4(n_0_28), 
      .ZN(n_0_1_79));
   NOR4_X1 i_0_1_100 (.A1(n_0_29), .A2(n_0_30), .A3(n_0_31), .A4(n_0_32), 
      .ZN(n_0_1_80));
   NAND3_X1 i_0_1_101 (.A1(n_0_1_86), .A2(n_0_1_85), .A3(n_0_1_82), .ZN(n_0_1_81));
   AND4_X1 i_0_1_102 (.A1(n_0_1_88), .A2(n_0_1_87), .A3(n_0_1_84), .A4(n_0_1_83), 
      .ZN(n_0_1_82));
   NOR4_X1 i_0_1_103 (.A1(n_0_68), .A2(n_0_70), .A3(n_0_64), .A4(n_0_67), 
      .ZN(n_0_1_83));
   NOR4_X1 i_0_1_104 (.A1(n_0_60), .A2(n_0_63), .A3(n_0_57), .A4(n_0_58), 
      .ZN(n_0_1_84));
   NOR3_X1 i_0_1_105 (.A1(n_0_65), .A2(n_0_66), .A3(n_0_69), .ZN(n_0_1_85));
   NOR4_X1 i_0_1_106 (.A1(n_0_61), .A2(n_0_62), .A3(n_0_56), .A4(n_0_59), 
      .ZN(n_0_1_86));
   NOR4_X1 i_0_1_107 (.A1(n_0_48), .A2(n_0_49), .A3(n_0_50), .A4(n_0_51), 
      .ZN(n_0_1_87));
   NOR4_X1 i_0_1_108 (.A1(n_0_52), .A2(n_0_53), .A3(n_0_54), .A4(n_0_55), 
      .ZN(n_0_1_88));
   INV_X1 i_0_1_109 (.A(n_0_1_90), .ZN(n_0_1_89));
   OAI22_X1 i_0_1_110 (.A1(n_0_1_100), .A2(n_0_1_94), .B1(n_0_1_97), .B2(
      n_0_1_91), .ZN(n_0_1_90));
   OR4_X1 i_0_1_111 (.A1(n_0_1_93), .A2(n_0_1_92), .A3(EB[5]), .A4(EB[4]), 
      .ZN(n_0_1_91));
   OR2_X1 i_0_1_112 (.A1(EB[7]), .A2(EB[6]), .ZN(n_0_1_92));
   OR4_X1 i_0_1_113 (.A1(EB[3]), .A2(EB[2]), .A3(EB[1]), .A4(EB[0]), .ZN(
      n_0_1_93));
   OR4_X1 i_0_1_114 (.A1(n_0_1_96), .A2(n_0_1_95), .A3(EA[5]), .A4(EA[4]), 
      .ZN(n_0_1_94));
   OR2_X1 i_0_1_115 (.A1(EA[7]), .A2(EA[6]), .ZN(n_0_1_95));
   OR4_X1 i_0_1_116 (.A1(EA[3]), .A2(EA[2]), .A3(EA[1]), .A4(EA[0]), .ZN(
      n_0_1_96));
   NAND3_X1 i_0_1_117 (.A1(EA[7]), .A2(n_0_1_98), .A3(EA[6]), .ZN(n_0_1_97));
   AND3_X1 i_0_1_118 (.A1(EA[2]), .A2(EA[1]), .A3(n_0_1_99), .ZN(n_0_1_98));
   AND4_X1 i_0_1_119 (.A1(EA[5]), .A2(EA[4]), .A3(EA[3]), .A4(EA[0]), .ZN(
      n_0_1_99));
   NAND3_X1 i_0_1_120 (.A1(EB[7]), .A2(n_0_1_101), .A3(EB[6]), .ZN(n_0_1_100));
   AND3_X1 i_0_1_121 (.A1(EB[2]), .A2(EB[1]), .A3(n_0_1_102), .ZN(n_0_1_101));
   AND4_X1 i_0_1_122 (.A1(EB[5]), .A2(EB[4]), .A3(EB[3]), .A4(EB[0]), .ZN(
      n_0_1_102));
   INV_X1 i_0_1_123 (.A(n_0_24), .ZN(n_0_1_103));
   AOI211_X1 i_0_1_124 (.A(reset), .B(n_0_1_104), .C1(B_reg), .C2(A_reg), 
      .ZN(n_0_102));
   NOR2_X1 i_0_1_196 (.A1(B_reg), .A2(A_reg), .ZN(n_0_1_104));
endmodule
