/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 16 23:26:02 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1899911067 */

module datapath__0_2(B_imm, A_imm, Res_imm);
   input [31:0]B_imm;
   input [31:0]A_imm;
   output [63:0]Res_imm;

   HA_X1 i_0 (.A(n_1538), .B(n_1723), .CO(n_1), .S(n_0));
   FA_X1 i_1 (.A(n_1514), .B(n_1537), .CI(n_1560), .CO(n_3), .S(n_2));
   HA_X1 i_2 (.A(n_1581), .B(n_1), .CO(n_5), .S(n_4));
   FA_X1 i_3 (.A(n_1559), .B(n_1580), .CI(n_5), .CO(n_8), .S(n_6));
   FA_X1 i_4 (.A(n_1466), .B(n_1489), .CI(n_1512), .CO(n_13), .S(n_9));
   FA_X1 i_5 (.A(n_1535), .B(n_1558), .CI(n_1579), .CO(n_15), .S(n_10));
   FA_X1 i_6 (.A(n_1442), .B(n_1465), .CI(n_1488), .CO(n_21), .S(n_12));
   FA_X1 i_7 (.A(n_1511), .B(n_1534), .CI(n_1557), .CO(n_23), .S(n_14));
   FA_X1 i_8 (.A(n_1578), .B(n_15), .CI(n_13), .CO(n_25), .S(n_20));
   FA_X1 i_9 (.A(n_1418), .B(n_1441), .CI(n_1464), .CO(n_31), .S(n_22));
   FA_X1 i_10 (.A(n_1487), .B(n_1510), .CI(n_1533), .CO(n_33), .S(n_24));
   FA_X1 i_11 (.A(n_1556), .B(n_1577), .CI(n_23), .CO(n_35), .S(n_34));
   FA_X1 i_12 (.A(n_21), .B(n_25), .CI(n_34), .CO(n_32), .S(n_30));
   FA_X1 i_13 (.A(n_1394), .B(n_1417), .CI(n_1440), .CO(n_43), .S(n_42));
   FA_X1 i_14 (.A(n_1463), .B(n_1486), .CI(n_1509), .CO(n_45), .S(n_44));
   FA_X1 i_15 (.A(n_1532), .B(n_1555), .CI(n_1576), .CO(n_47), .S(n_46));
   FA_X1 i_16 (.A(n_33), .B(n_31), .CI(n_35), .CO(n_49), .S(n_36));
   FA_X1 i_17 (.A(n_46), .B(n_44), .CI(n_42), .CO(n_48), .S(n_37));
   FA_X1 i_18 (.A(n_1370), .B(n_1393), .CI(n_1416), .CO(n_57), .S(n_56));
   FA_X1 i_19 (.A(n_1439), .B(n_1462), .CI(n_1485), .CO(n_59), .S(n_58));
   FA_X1 i_20 (.A(n_1508), .B(n_1531), .CI(n_1554), .CO(n_61), .S(n_60));
   FA_X1 i_21 (.A(n_1575), .B(n_47), .CI(n_45), .CO(n_63), .S(n_62));
   FA_X1 i_22 (.A(n_43), .B(n_60), .CI(n_58), .CO(n_65), .S(n_50));
   FA_X1 i_23 (.A(n_56), .B(n_49), .CI(n_62), .CO(n_64), .S(n_51));
   FA_X1 i_24 (.A(n_1346), .B(n_1369), .CI(n_1392), .CO(n_73), .S(n_72));
   FA_X1 i_25 (.A(n_1415), .B(n_1438), .CI(n_1461), .CO(n_75), .S(n_74));
   FA_X1 i_26 (.A(n_1484), .B(n_1507), .CI(n_1530), .CO(n_77), .S(n_76));
   FA_X1 i_27 (.A(n_1553), .B(n_1574), .CI(n_61), .CO(n_66), .S(n_78));
   FA_X1 i_28 (.A(n_59), .B(n_57), .CI(n_63), .CO(n_67), .S(n_80));
   FA_X1 i_29 (.A(n_78), .B(n_76), .CI(n_74), .CO(n_81), .S(n_79));
   FA_X1 i_30 (.A(n_72), .B(n_80), .CI(n_65), .CO(n_83), .S(n_82));
   FA_X1 i_45 (.A(n_1322), .B(n_1345), .CI(n_1368), .CO(n_85), .S(n_84));
   FA_X1 i_46 (.A(n_1391), .B(n_1414), .CI(n_1437), .CO(n_91), .S(n_90));
   FA_X1 i_47 (.A(n_1460), .B(n_1483), .CI(n_1506), .CO(n_95), .S(n_92));
   FA_X1 i_48 (.A(n_1529), .B(n_1552), .CI(n_1573), .CO(n_97), .S(n_93));
   FA_X1 i_31 (.A(n_77), .B(n_75), .CI(n_73), .CO(n_96), .S(n_94));
   FA_X1 i_32 (.A(n_1298), .B(n_1321), .CI(n_1344), .CO(n_99), .S(n_98));
   FA_X1 i_56 (.A(n_1367), .B(n_1390), .CI(n_1413), .CO(n_111), .S(n_110));
   FA_X1 i_57 (.A(n_1436), .B(n_1459), .CI(n_1482), .CO(n_113), .S(n_112));
   FA_X1 i_33 (.A(n_1505), .B(n_1528), .CI(n_1551), .CO(n_117), .S(n_114));
   FA_X1 i_34 (.A(n_1572), .B(n_97), .CI(n_95), .CO(n_116), .S(n_115));
   FA_X1 i_35 (.A(n_1274), .B(n_1297), .CI(n_1320), .CO(n_133), .S(n_118));
   FA_X1 i_36 (.A(n_1343), .B(n_1366), .CI(n_1389), .CO(n_135), .S(n_119));
   FA_X1 i_37 (.A(n_1412), .B(n_1435), .CI(n_1458), .CO(n_137), .S(n_132));
   FA_X1 i_38 (.A(n_1481), .B(n_1504), .CI(n_1527), .CO(n_139), .S(n_134));
   FA_X1 i_39 (.A(n_1550), .B(n_1571), .CI(n_117), .CO(n_141), .S(n_136));
   FA_X1 i_40 (.A(n_1250), .B(n_1273), .CI(n_1296), .CO(n_140), .S(n_138));
   FA_X1 i_41 (.A(n_1319), .B(n_1342), .CI(n_1365), .CO(n_156), .S(n_143));
   FA_X1 i_42 (.A(n_1388), .B(n_1411), .CI(n_1434), .CO(n_158), .S(n_157));
   FA_X1 i_43 (.A(n_1457), .B(n_1480), .CI(n_1503), .CO(n_160), .S(n_159));
   FA_X1 i_44 (.A(n_1526), .B(n_1549), .CI(n_1570), .CO(n_162), .S(n_161));
   FA_X1 i_49 (.A(n_139), .B(n_137), .CI(n_135), .CO(n_164), .S(n_163));
   FA_X1 i_50 (.A(n_133), .B(n_939), .CI(n_141), .CO(n_166), .S(n_165));
   FA_X1 i_51 (.A(n_1032), .B(n_1055), .CI(n_1078), .CO(n_551), .S(n_550));
   FA_X1 i_52 (.A(n_1101), .B(n_1124), .CI(n_1147), .CO(n_553), .S(n_552));
   FA_X1 i_53 (.A(n_1170), .B(n_1193), .CI(n_1216), .CO(n_555), .S(n_554));
   FA_X1 i_54 (.A(n_1239), .B(n_1262), .CI(n_1285), .CO(n_557), .S(n_556));
   FA_X1 i_55 (.A(n_1308), .B(n_1331), .CI(n_1354), .CO(n_559), .S(n_558));
   FA_X1 i_58 (.A(n_1377), .B(n_1400), .CI(n_1423), .CO(n_561), .S(n_560));
   FA_X1 i_59 (.A(n_1446), .B(n_1469), .CI(n_1492), .CO(n_563), .S(n_562));
   FA_X1 i_60 (.A(n_1515), .B(n_800), .CI(n_801), .CO(n_565), .S(n_564));
   FA_X1 i_61 (.A(n_788), .B(n_789), .CI(n_790), .CO(n_567), .S(n_566));
   FA_X1 i_62 (.A(n_785), .B(n_786), .CI(n_776), .CO(n_569), .S(n_568));
   FA_X1 i_63 (.A(n_778), .B(n_793), .CI(n_562), .CO(n_571), .S(n_570));
   FA_X1 i_64 (.A(n_560), .B(n_558), .CI(n_556), .CO(n_573), .S(n_572));
   FA_X1 i_65 (.A(n_554), .B(n_552), .CI(n_550), .CO(n_575), .S(n_574));
   FA_X1 i_66 (.A(n_829), .B(n_568), .CI(n_566), .CO(n_577), .S(n_576));
   FA_X1 i_67 (.A(n_564), .B(n_791), .CI(n_828), .CO(n_579), .S(n_578));
   FA_X1 i_68 (.A(n_787), .B(n_570), .CI(n_780), .CO(n_581), .S(n_580));
   FA_X1 i_69 (.A(n_574), .B(n_572), .CI(n_854), .CO(n_583), .S(n_582));
   FA_X1 i_70 (.A(n_578), .B(n_576), .CI(n_792), .CO(n_585), .S(n_584));
   FA_X1 i_71 (.A(n_580), .B(n_855), .CI(n_783), .CO(n_587), .S(n_586));
   FA_X1 i_72 (.A(n_582), .B(n_584), .CI(n_878), .CO(n_589), .S(n_588));
   FA_X1 i_73 (.A(n_586), .B(n_588), .CI(n_879), .CO(n_591), .S(n_590));
   FA_X1 i_74 (.A(n_1031), .B(n_1054), .CI(n_1077), .CO(n_593), .S(n_592));
   FA_X1 i_75 (.A(n_1100), .B(n_1123), .CI(n_1146), .CO(n_595), .S(n_594));
   FA_X1 i_76 (.A(n_1169), .B(n_1192), .CI(n_1215), .CO(n_597), .S(n_596));
   FA_X1 i_77 (.A(n_1238), .B(n_1261), .CI(n_1284), .CO(n_599), .S(n_598));
   FA_X1 i_78 (.A(n_1307), .B(n_1330), .CI(n_1353), .CO(n_601), .S(n_600));
   FA_X1 i_79 (.A(n_1376), .B(n_1399), .CI(n_1422), .CO(n_603), .S(n_602));
   FA_X1 i_80 (.A(n_1445), .B(n_1468), .CI(n_1491), .CO(n_605), .S(n_604));
   FA_X1 i_81 (.A(n_563), .B(n_561), .CI(n_559), .CO(n_607), .S(n_606));
   FA_X1 i_82 (.A(n_557), .B(n_555), .CI(n_553), .CO(n_609), .S(n_608));
   FA_X1 i_83 (.A(n_551), .B(n_567), .CI(n_565), .CO(n_611), .S(n_610));
   FA_X1 i_84 (.A(n_604), .B(n_602), .CI(n_600), .CO(n_613), .S(n_612));
   FA_X1 i_85 (.A(n_598), .B(n_596), .CI(n_594), .CO(n_615), .S(n_614));
   FA_X1 i_86 (.A(n_592), .B(n_569), .CI(n_608), .CO(n_617), .S(n_616));
   FA_X1 i_87 (.A(n_606), .B(n_575), .CI(n_573), .CO(n_619), .S(n_618));
   FA_X1 i_88 (.A(n_571), .B(n_610), .CI(n_579), .CO(n_621), .S(n_620));
   FA_X1 i_89 (.A(n_577), .B(n_614), .CI(n_612), .CO(n_623), .S(n_622));
   FA_X1 i_90 (.A(n_616), .B(n_581), .CI(n_618), .CO(n_625), .S(n_624));
   FA_X1 i_91 (.A(n_583), .B(n_620), .CI(n_585), .CO(n_627), .S(n_626));
   FA_X1 i_92 (.A(n_622), .B(n_624), .CI(n_587), .CO(n_167), .S(n_628));
   FA_X1 i_93 (.A(n_626), .B(n_589), .CI(n_628), .CO(n_168), .S(n_630));
   FA_X1 i_94 (.A(n_1030), .B(n_1053), .CI(n_1076), .CO(n_633), .S(n_632));
   FA_X1 i_95 (.A(n_1099), .B(n_1122), .CI(n_1145), .CO(n_635), .S(n_634));
   FA_X1 i_96 (.A(n_1168), .B(n_1191), .CI(n_1214), .CO(n_637), .S(n_636));
   FA_X1 i_97 (.A(n_1237), .B(n_1260), .CI(n_1283), .CO(n_639), .S(n_638));
   FA_X1 i_98 (.A(n_1306), .B(n_1329), .CI(n_1352), .CO(n_641), .S(n_640));
   FA_X1 i_99 (.A(n_1375), .B(n_1398), .CI(n_1421), .CO(n_643), .S(n_642));
   FA_X1 i_100 (.A(n_1444), .B(n_1467), .CI(n_605), .CO(n_645), .S(n_644));
   FA_X1 i_101 (.A(n_603), .B(n_601), .CI(n_599), .CO(n_647), .S(n_646));
   FA_X1 i_102 (.A(n_597), .B(n_595), .CI(n_593), .CO(n_649), .S(n_648));
   FA_X1 i_103 (.A(n_609), .B(n_607), .CI(n_644), .CO(n_651), .S(n_650));
   FA_X1 i_104 (.A(n_642), .B(n_640), .CI(n_638), .CO(n_653), .S(n_652));
   FA_X1 i_105 (.A(n_636), .B(n_634), .CI(n_632), .CO(n_655), .S(n_654));
   FA_X1 i_106 (.A(n_611), .B(n_648), .CI(n_646), .CO(n_657), .S(n_656));
   FA_X1 i_107 (.A(n_615), .B(n_613), .CI(n_650), .CO(n_659), .S(n_658));
   FA_X1 i_108 (.A(n_619), .B(n_617), .CI(n_654), .CO(n_661), .S(n_660));
   FA_X1 i_109 (.A(n_652), .B(n_621), .CI(n_658), .CO(n_663), .S(n_662));
   FA_X1 i_110 (.A(n_656), .B(n_623), .CI(n_660), .CO(n_665), .S(n_169));
   FA_X1 i_111 (.A(n_625), .B(n_662), .CI(n_627), .CO(n_504), .S(n_461));
   FA_X1 i_112 (.A(n_1029), .B(n_1052), .CI(n_1075), .CO(n_671), .S(n_670));
   FA_X1 i_113 (.A(n_1098), .B(n_1121), .CI(n_1144), .CO(n_673), .S(n_672));
   FA_X1 i_114 (.A(n_1167), .B(n_1190), .CI(n_1213), .CO(n_675), .S(n_674));
   FA_X1 i_115 (.A(n_1236), .B(n_1259), .CI(n_1282), .CO(n_677), .S(n_676));
   FA_X1 i_116 (.A(n_1305), .B(n_1328), .CI(n_1351), .CO(n_679), .S(n_678));
   FA_X1 i_117 (.A(n_1374), .B(n_1397), .CI(n_1420), .CO(n_681), .S(n_680));
   FA_X1 i_118 (.A(n_1443), .B(n_643), .CI(n_641), .CO(n_683), .S(n_682));
   FA_X1 i_119 (.A(n_639), .B(n_637), .CI(n_635), .CO(n_685), .S(n_684));
   FA_X1 i_120 (.A(n_633), .B(n_649), .CI(n_647), .CO(n_687), .S(n_686));
   FA_X1 i_121 (.A(n_645), .B(n_680), .CI(n_678), .CO(n_689), .S(n_688));
   FA_X1 i_122 (.A(n_676), .B(n_674), .CI(n_672), .CO(n_691), .S(n_690));
   FA_X1 i_123 (.A(n_670), .B(n_684), .CI(n_682), .CO(n_693), .S(n_692));
   FA_X1 i_124 (.A(n_655), .B(n_653), .CI(n_651), .CO(n_695), .S(n_694));
   FA_X1 i_125 (.A(n_686), .B(n_657), .CI(n_690), .CO(n_697), .S(n_696));
   FA_X1 i_126 (.A(n_688), .B(n_659), .CI(n_694), .CO(n_699), .S(n_698));
   FA_X1 i_127 (.A(n_692), .B(n_661), .CI(n_696), .CO(n_701), .S(n_505));
   FA_X1 i_128 (.A(n_663), .B(n_698), .CI(n_665), .CO(n_509), .S(n_507));
   FA_X1 i_129 (.A(n_1028), .B(n_1051), .CI(n_1074), .CO(n_707), .S(n_706));
   FA_X1 i_130 (.A(n_1097), .B(n_1120), .CI(n_1143), .CO(n_709), .S(n_708));
   FA_X1 i_131 (.A(n_1166), .B(n_1189), .CI(n_1212), .CO(n_711), .S(n_710));
   FA_X1 i_132 (.A(n_1235), .B(n_1258), .CI(n_1281), .CO(n_713), .S(n_712));
   FA_X1 i_133 (.A(n_1304), .B(n_1327), .CI(n_1350), .CO(n_715), .S(n_714));
   FA_X1 i_134 (.A(n_1373), .B(n_1396), .CI(n_1419), .CO(n_717), .S(n_716));
   FA_X1 i_135 (.A(n_681), .B(n_679), .CI(n_677), .CO(n_719), .S(n_718));
   FA_X1 i_136 (.A(n_675), .B(n_673), .CI(n_671), .CO(n_721), .S(n_720));
   FA_X1 i_137 (.A(n_685), .B(n_683), .CI(n_716), .CO(n_723), .S(n_722));
   FA_X1 i_138 (.A(n_714), .B(n_712), .CI(n_710), .CO(n_725), .S(n_724));
   FA_X1 i_139 (.A(n_708), .B(n_706), .CI(n_687), .CO(n_727), .S(n_726));
   FA_X1 i_140 (.A(n_720), .B(n_718), .CI(n_691), .CO(n_511), .S(n_728));
   FA_X1 i_141 (.A(n_689), .B(n_722), .CI(n_695), .CO(n_513), .S(n_730));
   FA_X1 i_142 (.A(n_693), .B(n_726), .CI(n_724), .CO(n_733), .S(n_732));
   FA_X1 i_143 (.A(n_728), .B(n_697), .CI(n_730), .CO(n_735), .S(n_515));
   FA_X1 i_144 (.A(n_699), .B(n_732), .CI(n_701), .CO(n_519), .S(n_517));
   FA_X1 i_145 (.A(n_1027), .B(n_1050), .CI(n_1073), .CO(n_741), .S(n_740));
   FA_X1 i_146 (.A(n_1096), .B(n_1119), .CI(n_1142), .CO(n_743), .S(n_742));
   FA_X1 i_147 (.A(n_1165), .B(n_1188), .CI(n_1211), .CO(n_745), .S(n_744));
   FA_X1 i_148 (.A(n_1234), .B(n_1257), .CI(n_1280), .CO(n_747), .S(n_746));
   FA_X1 i_149 (.A(n_1303), .B(n_1326), .CI(n_1349), .CO(n_749), .S(n_748));
   FA_X1 i_150 (.A(n_1372), .B(n_1395), .CI(n_717), .CO(n_751), .S(n_750));
   FA_X1 i_151 (.A(n_715), .B(n_713), .CI(n_711), .CO(n_753), .S(n_752));
   FA_X1 i_152 (.A(n_709), .B(n_707), .CI(n_721), .CO(n_755), .S(n_754));
   FA_X1 i_153 (.A(n_719), .B(n_750), .CI(n_748), .CO(n_757), .S(n_521));
   FA_X1 i_154 (.A(n_746), .B(n_744), .CI(n_742), .CO(n_759), .S(n_523));
   FA_X1 i_155 (.A(n_740), .B(n_754), .CI(n_752), .CO(n_527), .S(n_525));
   FA_X1 i_156 (.A(n_725), .B(n_723), .CI(n_727), .CO(n_531), .S(n_529));
   FA_X1 i_157 (.A(n_733), .B(n_1700), .CI(n_735), .CO(n_535), .S(n_533));
   FA_X1 i_158 (.A(n_1026), .B(n_1049), .CI(n_1072), .CO(n_537), .S(n_772));
   FA_X1 i_159 (.A(n_1095), .B(n_1118), .CI(n_1141), .CO(n_539), .S(n_774));
   FA_X1 i_160 (.A(n_1371), .B(n_749), .CI(n_747), .CO(n_541), .S(n_782));
   FA_X1 i_161 (.A(n_745), .B(n_743), .CI(n_741), .CO(n_543), .S(n_784));
   FA_X1 i_162 (.A(n_753), .B(n_751), .CI(n_1688), .CO(n_547), .S(n_545));
   FA_X1 i_163 (.A(n_1690), .B(n_1691), .CI(n_774), .CO(n_549), .S(n_548));
   FA_X1 i_164 (.A(n_772), .B(n_755), .CI(n_784), .CO(n_631), .S(n_629));
   FA_X1 i_165 (.A(n_782), .B(n_759), .CI(n_757), .CO(n_666), .S(n_664));
   NOR2_X1 i_166 (.A1(n_1654), .A2(n_1639), .ZN(n_1026));
   NOR2_X1 i_167 (.A1(n_1654), .A2(n_1634), .ZN(n_1027));
   NOR2_X1 i_168 (.A1(n_1654), .A2(n_1633), .ZN(n_1028));
   NOR2_X1 i_169 (.A1(n_1654), .A2(n_1632), .ZN(n_1029));
   NOR2_X1 i_170 (.A1(n_1654), .A2(n_1631), .ZN(n_1030));
   NOR2_X1 i_171 (.A1(n_1654), .A2(n_1630), .ZN(n_1031));
   NOR2_X1 i_172 (.A1(n_1654), .A2(n_1629), .ZN(n_1032));
   NOR2_X1 i_173 (.A1(n_1678), .A2(n_1640), .ZN(n_1049));
   NOR2_X1 i_174 (.A1(n_1678), .A2(n_1639), .ZN(n_1050));
   NOR2_X1 i_175 (.A1(n_1678), .A2(n_1634), .ZN(n_1051));
   NOR2_X1 i_176 (.A1(n_1678), .A2(n_1633), .ZN(n_1052));
   NOR2_X1 i_177 (.A1(n_1678), .A2(n_1632), .ZN(n_1053));
   NOR2_X1 i_178 (.A1(n_1678), .A2(n_1631), .ZN(n_1054));
   NOR2_X1 i_179 (.A1(n_1678), .A2(n_1630), .ZN(n_1055));
   NOR2_X1 i_180 (.A1(n_1677), .A2(n_1641), .ZN(n_1072));
   NOR2_X1 i_181 (.A1(n_1677), .A2(n_1640), .ZN(n_1073));
   NOR2_X1 i_182 (.A1(n_1677), .A2(n_1639), .ZN(n_1074));
   NOR2_X1 i_183 (.A1(n_1677), .A2(n_1634), .ZN(n_1075));
   NOR2_X1 i_184 (.A1(n_1677), .A2(n_1633), .ZN(n_1076));
   NOR2_X1 i_185 (.A1(n_1677), .A2(n_1632), .ZN(n_1077));
   NOR2_X1 i_186 (.A1(n_1677), .A2(n_1631), .ZN(n_1078));
   NOR2_X1 i_187 (.A1(n_1676), .A2(n_1642), .ZN(n_1095));
   NOR2_X1 i_188 (.A1(n_1676), .A2(n_1641), .ZN(n_1096));
   NOR2_X1 i_189 (.A1(n_1676), .A2(n_1640), .ZN(n_1097));
   NOR2_X1 i_190 (.A1(n_1676), .A2(n_1639), .ZN(n_1098));
   NOR2_X1 i_191 (.A1(n_1676), .A2(n_1634), .ZN(n_1099));
   NOR2_X1 i_192 (.A1(n_1676), .A2(n_1633), .ZN(n_1100));
   NOR2_X1 i_193 (.A1(n_1676), .A2(n_1632), .ZN(n_1101));
   NOR2_X1 i_194 (.A1(n_1675), .A2(n_1643), .ZN(n_1118));
   NOR2_X1 i_195 (.A1(n_1675), .A2(n_1642), .ZN(n_1119));
   NOR2_X1 i_196 (.A1(n_1675), .A2(n_1641), .ZN(n_1120));
   NOR2_X1 i_197 (.A1(n_1675), .A2(n_1640), .ZN(n_1121));
   NOR2_X1 i_198 (.A1(n_1675), .A2(n_1639), .ZN(n_1122));
   NOR2_X1 i_199 (.A1(n_1675), .A2(n_1634), .ZN(n_1123));
   NOR2_X1 i_200 (.A1(n_1675), .A2(n_1633), .ZN(n_1124));
   NOR2_X1 i_201 (.A1(n_1674), .A2(n_1644), .ZN(n_1141));
   NOR2_X1 i_202 (.A1(n_1674), .A2(n_1643), .ZN(n_1142));
   NOR2_X1 i_203 (.A1(n_1674), .A2(n_1642), .ZN(n_1143));
   NOR2_X1 i_204 (.A1(n_1674), .A2(n_1641), .ZN(n_1144));
   NOR2_X1 i_205 (.A1(n_1674), .A2(n_1640), .ZN(n_1145));
   NOR2_X1 i_206 (.A1(n_1674), .A2(n_1639), .ZN(n_1146));
   NOR2_X1 i_207 (.A1(n_1674), .A2(n_1634), .ZN(n_1147));
   NOR2_X1 i_208 (.A1(n_1673), .A2(n_1645), .ZN(n_667));
   NOR2_X1 i_209 (.A1(n_1673), .A2(n_1644), .ZN(n_1165));
   NOR2_X1 i_210 (.A1(n_1673), .A2(n_1643), .ZN(n_1166));
   NOR2_X1 i_211 (.A1(n_1673), .A2(n_1642), .ZN(n_1167));
   NOR2_X1 i_212 (.A1(n_1673), .A2(n_1641), .ZN(n_1168));
   NOR2_X1 i_213 (.A1(n_1673), .A2(n_1640), .ZN(n_1169));
   NOR2_X1 i_214 (.A1(n_1673), .A2(n_1639), .ZN(n_1170));
   NOR2_X1 i_215 (.A1(n_1672), .A2(n_1646), .ZN(n_668));
   NOR2_X1 i_216 (.A1(n_1672), .A2(n_1645), .ZN(n_1188));
   NOR2_X1 i_217 (.A1(n_1672), .A2(n_1644), .ZN(n_1189));
   NOR2_X1 i_218 (.A1(n_1672), .A2(n_1643), .ZN(n_1190));
   NOR2_X1 i_219 (.A1(n_1672), .A2(n_1642), .ZN(n_1191));
   NOR2_X1 i_220 (.A1(n_1672), .A2(n_1641), .ZN(n_1192));
   NOR2_X1 i_221 (.A1(n_1672), .A2(n_1640), .ZN(n_1193));
   NOR2_X1 i_222 (.A1(n_1670), .A2(n_1647), .ZN(n_669));
   NOR2_X1 i_223 (.A1(n_1670), .A2(n_1646), .ZN(n_1211));
   NOR2_X1 i_224 (.A1(n_1670), .A2(n_1645), .ZN(n_1212));
   NOR2_X1 i_225 (.A1(n_1670), .A2(n_1644), .ZN(n_1213));
   NOR2_X1 i_226 (.A1(n_1670), .A2(n_1643), .ZN(n_1214));
   NOR2_X1 i_227 (.A1(n_1670), .A2(n_1642), .ZN(n_1215));
   NOR2_X1 i_228 (.A1(n_1670), .A2(n_1641), .ZN(n_1216));
   NOR2_X1 i_229 (.A1(n_1670), .A2(n_1625), .ZN(n_700));
   NOR2_X1 i_230 (.A1(n_1669), .A2(n_1648), .ZN(n_702));
   NOR2_X1 i_231 (.A1(n_1669), .A2(n_1647), .ZN(n_1234));
   NOR2_X1 i_232 (.A1(n_1669), .A2(n_1646), .ZN(n_1235));
   NOR2_X1 i_233 (.A1(n_1669), .A2(n_1645), .ZN(n_1236));
   NOR2_X1 i_234 (.A1(n_1669), .A2(n_1644), .ZN(n_1237));
   NOR2_X1 i_235 (.A1(n_1669), .A2(n_1643), .ZN(n_1238));
   NOR2_X1 i_236 (.A1(n_1669), .A2(n_1642), .ZN(n_1239));
   NOR2_X1 i_237 (.A1(n_1669), .A2(n_1628), .ZN(n_703));
   NOR2_X1 i_744 (.A1(n_1669), .A2(n_1625), .ZN(n_1250));
   NOR2_X1 i_238 (.A1(n_1668), .A2(n_1649), .ZN(n_704));
   NOR2_X1 i_239 (.A1(n_1668), .A2(n_1648), .ZN(n_1257));
   NOR2_X1 i_240 (.A1(n_1668), .A2(n_1647), .ZN(n_1258));
   NOR2_X1 i_241 (.A1(n_1668), .A2(n_1646), .ZN(n_1259));
   NOR2_X1 i_242 (.A1(n_1668), .A2(n_1645), .ZN(n_1260));
   NOR2_X1 i_243 (.A1(n_1668), .A2(n_1644), .ZN(n_1261));
   NOR2_X1 i_244 (.A1(n_1668), .A2(n_1643), .ZN(n_1262));
   NOR2_X1 i_245 (.A1(n_1668), .A2(n_1629), .ZN(n_705));
   NOR2_X1 i_767 (.A1(n_1668), .A2(n_1628), .ZN(n_1273));
   NOR2_X1 i_246 (.A1(n_1668), .A2(n_1625), .ZN(n_1274));
   NOR2_X1 i_247 (.A1(n_1667), .A2(n_1650), .ZN(n_729));
   NOR2_X1 i_248 (.A1(n_1667), .A2(n_1649), .ZN(n_1280));
   NOR2_X1 i_249 (.A1(n_1667), .A2(n_1648), .ZN(n_1281));
   NOR2_X1 i_250 (.A1(n_1667), .A2(n_1647), .ZN(n_1282));
   NOR2_X1 i_251 (.A1(n_1667), .A2(n_1646), .ZN(n_1283));
   NOR2_X1 i_252 (.A1(n_1667), .A2(n_1645), .ZN(n_1284));
   NOR2_X1 i_253 (.A1(n_1667), .A2(n_1644), .ZN(n_1285));
   NOR2_X1 i_790 (.A1(n_1667), .A2(n_1629), .ZN(n_1296));
   NOR2_X1 i_254 (.A1(n_1667), .A2(n_1628), .ZN(n_1297));
   NOR2_X1 i_792 (.A1(n_1667), .A2(n_1625), .ZN(n_1298));
   NOR2_X1 i_255 (.A1(n_1666), .A2(n_1651), .ZN(n_731));
   NOR2_X1 i_256 (.A1(n_1666), .A2(n_1650), .ZN(n_1303));
   NOR2_X1 i_257 (.A1(n_1666), .A2(n_1649), .ZN(n_1304));
   NOR2_X1 i_258 (.A1(n_1666), .A2(n_1648), .ZN(n_1305));
   NOR2_X1 i_259 (.A1(n_1666), .A2(n_1647), .ZN(n_1306));
   NOR2_X1 i_260 (.A1(n_1666), .A2(n_1646), .ZN(n_1307));
   NOR2_X1 i_261 (.A1(n_1666), .A2(n_1645), .ZN(n_1308));
   NOR2_X1 i_813 (.A1(n_1666), .A2(n_1630), .ZN(n_1319));
   NOR2_X1 i_262 (.A1(n_1666), .A2(n_1629), .ZN(n_1320));
   NOR2_X1 i_815 (.A1(n_1666), .A2(n_1628), .ZN(n_1321));
   NOR2_X1 i_816 (.A1(n_1666), .A2(n_1625), .ZN(n_1322));
   NOR2_X1 i_263 (.A1(n_1665), .A2(n_1652), .ZN(n_734));
   NOR2_X1 i_264 (.A1(n_1665), .A2(n_1651), .ZN(n_1326));
   NOR2_X1 i_265 (.A1(n_1665), .A2(n_1650), .ZN(n_1327));
   NOR2_X1 i_266 (.A1(n_1665), .A2(n_1649), .ZN(n_1328));
   NOR2_X1 i_267 (.A1(n_1665), .A2(n_1648), .ZN(n_1329));
   NOR2_X1 i_268 (.A1(n_1665), .A2(n_1647), .ZN(n_1330));
   NOR2_X1 i_269 (.A1(n_1665), .A2(n_1646), .ZN(n_1331));
   NOR2_X1 i_836 (.A1(n_1665), .A2(n_1631), .ZN(n_1342));
   NOR2_X1 i_837 (.A1(n_1665), .A2(n_1630), .ZN(n_1343));
   NOR2_X1 i_838 (.A1(n_1665), .A2(n_1629), .ZN(n_1344));
   NOR2_X1 i_839 (.A1(n_1665), .A2(n_1628), .ZN(n_1345));
   NOR2_X1 i_270 (.A1(n_1665), .A2(n_1625), .ZN(n_1346));
   NOR2_X1 i_271 (.A1(n_1664), .A2(n_1653), .ZN(n_736));
   NOR2_X1 i_272 (.A1(n_1664), .A2(n_1652), .ZN(n_1349));
   NOR2_X1 i_273 (.A1(n_1664), .A2(n_1651), .ZN(n_1350));
   NOR2_X1 i_274 (.A1(n_1664), .A2(n_1650), .ZN(n_1351));
   NOR2_X1 i_275 (.A1(n_1664), .A2(n_1649), .ZN(n_1352));
   NOR2_X1 i_276 (.A1(n_1664), .A2(n_1648), .ZN(n_1353));
   NOR2_X1 i_277 (.A1(n_1664), .A2(n_1647), .ZN(n_1354));
   NOR2_X1 i_859 (.A1(n_1664), .A2(n_1632), .ZN(n_1365));
   NOR2_X1 i_860 (.A1(n_1664), .A2(n_1631), .ZN(n_1366));
   NOR2_X1 i_861 (.A1(n_1664), .A2(n_1630), .ZN(n_1367));
   NOR2_X1 i_862 (.A1(n_1664), .A2(n_1629), .ZN(n_1368));
   NOR2_X1 i_278 (.A1(n_1664), .A2(n_1628), .ZN(n_1369));
   NOR2_X1 i_279 (.A1(n_1664), .A2(n_1625), .ZN(n_1370));
   NOR2_X1 i_280 (.A1(n_1663), .A2(n_1654), .ZN(n_1371));
   NOR2_X1 i_281 (.A1(n_1663), .A2(n_1653), .ZN(n_1372));
   NOR2_X1 i_282 (.A1(n_1663), .A2(n_1652), .ZN(n_1373));
   NOR2_X1 i_283 (.A1(n_1663), .A2(n_1651), .ZN(n_1374));
   NOR2_X1 i_284 (.A1(n_1663), .A2(n_1650), .ZN(n_1375));
   NOR2_X1 i_285 (.A1(n_1663), .A2(n_1649), .ZN(n_1376));
   NOR2_X1 i_286 (.A1(n_1663), .A2(n_1648), .ZN(n_1377));
   NOR2_X1 i_882 (.A1(n_1663), .A2(n_1633), .ZN(n_1388));
   NOR2_X1 i_883 (.A1(n_1663), .A2(n_1632), .ZN(n_1389));
   NOR2_X1 i_884 (.A1(n_1663), .A2(n_1631), .ZN(n_1390));
   NOR2_X1 i_885 (.A1(n_1663), .A2(n_1630), .ZN(n_1391));
   NOR2_X1 i_287 (.A1(n_1663), .A2(n_1629), .ZN(n_1392));
   NOR2_X1 i_288 (.A1(n_1663), .A2(n_1628), .ZN(n_1393));
   NOR2_X1 i_289 (.A1(n_1663), .A2(n_1625), .ZN(n_1394));
   NOR2_X1 i_290 (.A1(n_1662), .A2(n_1654), .ZN(n_1395));
   NOR2_X1 i_291 (.A1(n_1662), .A2(n_1653), .ZN(n_1396));
   NOR2_X1 i_292 (.A1(n_1662), .A2(n_1652), .ZN(n_1397));
   NOR2_X1 i_293 (.A1(n_1662), .A2(n_1651), .ZN(n_1398));
   NOR2_X1 i_294 (.A1(n_1662), .A2(n_1650), .ZN(n_1399));
   NOR2_X1 i_295 (.A1(n_1662), .A2(n_1649), .ZN(n_1400));
   NOR2_X1 i_905 (.A1(n_1662), .A2(n_1634), .ZN(n_1411));
   NOR2_X1 i_906 (.A1(n_1662), .A2(n_1633), .ZN(n_1412));
   NOR2_X1 i_907 (.A1(n_1662), .A2(n_1632), .ZN(n_1413));
   NOR2_X1 i_908 (.A1(n_1662), .A2(n_1631), .ZN(n_1414));
   NOR2_X1 i_296 (.A1(n_1662), .A2(n_1630), .ZN(n_1415));
   NOR2_X1 i_297 (.A1(n_1662), .A2(n_1629), .ZN(n_1416));
   NOR2_X1 i_298 (.A1(n_1662), .A2(n_1628), .ZN(n_1417));
   NOR2_X1 i_299 (.A1(n_1662), .A2(n_1625), .ZN(n_1418));
   NOR2_X1 i_300 (.A1(n_1661), .A2(n_1654), .ZN(n_1419));
   NOR2_X1 i_301 (.A1(n_1661), .A2(n_1653), .ZN(n_1420));
   NOR2_X1 i_302 (.A1(n_1661), .A2(n_1652), .ZN(n_1421));
   NOR2_X1 i_303 (.A1(n_1661), .A2(n_1651), .ZN(n_1422));
   NOR2_X1 i_304 (.A1(n_1661), .A2(n_1650), .ZN(n_1423));
   NOR2_X1 i_928 (.A1(n_1661), .A2(n_1639), .ZN(n_1434));
   NOR2_X1 i_929 (.A1(n_1661), .A2(n_1634), .ZN(n_1435));
   NOR2_X1 i_930 (.A1(n_1661), .A2(n_1633), .ZN(n_1436));
   NOR2_X1 i_931 (.A1(n_1661), .A2(n_1632), .ZN(n_1437));
   NOR2_X1 i_305 (.A1(n_1661), .A2(n_1631), .ZN(n_1438));
   NOR2_X1 i_306 (.A1(n_1661), .A2(n_1630), .ZN(n_1439));
   NOR2_X1 i_307 (.A1(n_1661), .A2(n_1629), .ZN(n_1440));
   NOR2_X1 i_308 (.A1(n_1661), .A2(n_1628), .ZN(n_1441));
   NOR2_X1 i_309 (.A1(n_1661), .A2(n_1625), .ZN(n_1442));
   NOR2_X1 i_310 (.A1(n_1660), .A2(n_1654), .ZN(n_1443));
   NOR2_X1 i_311 (.A1(n_1660), .A2(n_1653), .ZN(n_1444));
   NOR2_X1 i_312 (.A1(n_1660), .A2(n_1652), .ZN(n_1445));
   NOR2_X1 i_313 (.A1(n_1660), .A2(n_1651), .ZN(n_1446));
   NOR2_X1 i_951 (.A1(n_1660), .A2(n_1640), .ZN(n_1457));
   NOR2_X1 i_952 (.A1(n_1660), .A2(n_1639), .ZN(n_1458));
   NOR2_X1 i_953 (.A1(n_1660), .A2(n_1634), .ZN(n_1459));
   NOR2_X1 i_954 (.A1(n_1660), .A2(n_1633), .ZN(n_1460));
   NOR2_X1 i_314 (.A1(n_1660), .A2(n_1632), .ZN(n_1461));
   NOR2_X1 i_315 (.A1(n_1660), .A2(n_1631), .ZN(n_1462));
   NOR2_X1 i_316 (.A1(n_1660), .A2(n_1630), .ZN(n_1463));
   NOR2_X1 i_317 (.A1(n_1660), .A2(n_1629), .ZN(n_1464));
   NOR2_X1 i_318 (.A1(n_1660), .A2(n_1628), .ZN(n_1465));
   NOR2_X1 i_319 (.A1(n_1660), .A2(n_1625), .ZN(n_1466));
   NOR2_X1 i_320 (.A1(n_1659), .A2(n_1654), .ZN(n_1467));
   NOR2_X1 i_321 (.A1(n_1659), .A2(n_1653), .ZN(n_1468));
   NOR2_X1 i_322 (.A1(n_1659), .A2(n_1652), .ZN(n_1469));
   NOR2_X1 i_974 (.A1(n_1659), .A2(n_1641), .ZN(n_1480));
   NOR2_X1 i_975 (.A1(n_1659), .A2(n_1640), .ZN(n_1481));
   NOR2_X1 i_976 (.A1(n_1659), .A2(n_1639), .ZN(n_1482));
   NOR2_X1 i_977 (.A1(n_1659), .A2(n_1634), .ZN(n_1483));
   NOR2_X1 i_323 (.A1(n_1659), .A2(n_1633), .ZN(n_1484));
   NOR2_X1 i_324 (.A1(n_1659), .A2(n_1632), .ZN(n_1485));
   NOR2_X1 i_325 (.A1(n_1659), .A2(n_1631), .ZN(n_1486));
   NOR2_X1 i_326 (.A1(n_1659), .A2(n_1630), .ZN(n_1487));
   NOR2_X1 i_327 (.A1(n_1659), .A2(n_1629), .ZN(n_1488));
   NOR2_X1 i_328 (.A1(n_1659), .A2(n_1628), .ZN(n_1489));
   NOR2_X1 i_329 (.A1(n_1659), .A2(n_1625), .ZN(n_737));
   NOR2_X1 i_330 (.A1(n_1658), .A2(n_1654), .ZN(n_1491));
   NOR2_X1 i_331 (.A1(n_1658), .A2(n_1653), .ZN(n_1492));
   NOR2_X1 i_997 (.A1(n_1658), .A2(n_1642), .ZN(n_1503));
   NOR2_X1 i_998 (.A1(n_1658), .A2(n_1641), .ZN(n_1504));
   NOR2_X1 i_332 (.A1(n_1658), .A2(n_1640), .ZN(n_1505));
   NOR2_X1 i_1000 (.A1(n_1658), .A2(n_1639), .ZN(n_1506));
   NOR2_X1 i_333 (.A1(n_1658), .A2(n_1634), .ZN(n_1507));
   NOR2_X1 i_334 (.A1(n_1658), .A2(n_1633), .ZN(n_1508));
   NOR2_X1 i_335 (.A1(n_1658), .A2(n_1632), .ZN(n_1509));
   NOR2_X1 i_336 (.A1(n_1658), .A2(n_1631), .ZN(n_1510));
   NOR2_X1 i_337 (.A1(n_1658), .A2(n_1630), .ZN(n_1511));
   NOR2_X1 i_338 (.A1(n_1658), .A2(n_1629), .ZN(n_1512));
   NOR2_X1 i_339 (.A1(n_1658), .A2(n_1628), .ZN(n_738));
   NOR2_X1 i_340 (.A1(n_1658), .A2(n_1625), .ZN(n_1514));
   NOR2_X1 i_341 (.A1(n_1657), .A2(n_1654), .ZN(n_1515));
   NOR2_X1 i_1020 (.A1(n_1657), .A2(n_1643), .ZN(n_1526));
   NOR2_X1 i_1021 (.A1(n_1657), .A2(n_1642), .ZN(n_1527));
   NOR2_X1 i_342 (.A1(n_1657), .A2(n_1641), .ZN(n_1528));
   NOR2_X1 i_1023 (.A1(n_1657), .A2(n_1640), .ZN(n_1529));
   NOR2_X1 i_343 (.A1(n_1657), .A2(n_1639), .ZN(n_1530));
   NOR2_X1 i_344 (.A1(n_1657), .A2(n_1634), .ZN(n_1531));
   NOR2_X1 i_345 (.A1(n_1657), .A2(n_1633), .ZN(n_1532));
   NOR2_X1 i_346 (.A1(n_1657), .A2(n_1632), .ZN(n_1533));
   NOR2_X1 i_347 (.A1(n_1657), .A2(n_1631), .ZN(n_1534));
   NOR2_X1 i_348 (.A1(n_1657), .A2(n_1630), .ZN(n_1535));
   NOR2_X1 i_349 (.A1(n_1657), .A2(n_1629), .ZN(n_739));
   NOR2_X1 i_350 (.A1(n_1657), .A2(n_1628), .ZN(n_1537));
   NOR2_X1 i_351 (.A1(n_1657), .A2(n_1625), .ZN(n_1538));
   NOR2_X1 i_1043 (.A1(n_1656), .A2(n_1644), .ZN(n_1549));
   NOR2_X1 i_352 (.A1(n_1656), .A2(n_1643), .ZN(n_1550));
   NOR2_X1 i_353 (.A1(n_1656), .A2(n_1642), .ZN(n_1551));
   NOR2_X1 i_1046 (.A1(n_1656), .A2(n_1641), .ZN(n_1552));
   NOR2_X1 i_354 (.A1(n_1656), .A2(n_1640), .ZN(n_1553));
   NOR2_X1 i_355 (.A1(n_1656), .A2(n_1639), .ZN(n_1554));
   NOR2_X1 i_356 (.A1(n_1656), .A2(n_1634), .ZN(n_1555));
   NOR2_X1 i_357 (.A1(n_1656), .A2(n_1633), .ZN(n_1556));
   NOR2_X1 i_358 (.A1(n_1656), .A2(n_1632), .ZN(n_1557));
   NOR2_X1 i_359 (.A1(n_1656), .A2(n_1631), .ZN(n_1558));
   NOR2_X1 i_360 (.A1(n_1656), .A2(n_1630), .ZN(n_1559));
   NOR2_X1 i_361 (.A1(n_1656), .A2(n_1629), .ZN(n_1560));
   NOR2_X1 i_362 (.A1(n_1655), .A2(n_1646), .ZN(n_756));
   NOR2_X1 i_1064 (.A1(n_1655), .A2(n_1645), .ZN(n_1570));
   NOR2_X1 i_363 (.A1(n_1655), .A2(n_1644), .ZN(n_1571));
   NOR2_X1 i_1066 (.A1(n_1655), .A2(n_1643), .ZN(n_1572));
   NOR2_X1 i_1067 (.A1(n_1655), .A2(n_1642), .ZN(n_1573));
   NOR2_X1 i_364 (.A1(n_1655), .A2(n_1641), .ZN(n_1574));
   NOR2_X1 i_365 (.A1(n_1655), .A2(n_1640), .ZN(n_1575));
   NOR2_X1 i_366 (.A1(n_1655), .A2(n_1639), .ZN(n_1576));
   NOR2_X1 i_367 (.A1(n_1655), .A2(n_1634), .ZN(n_1577));
   NOR2_X1 i_368 (.A1(n_1655), .A2(n_1633), .ZN(n_1578));
   NOR2_X1 i_369 (.A1(n_1655), .A2(n_1632), .ZN(n_1579));
   NOR2_X1 i_370 (.A1(n_1655), .A2(n_1631), .ZN(n_1580));
   NOR2_X1 i_371 (.A1(n_1655), .A2(n_1630), .ZN(n_1581));
   XOR2_X1 i_372 (.A(n_973), .B(n_1582), .Z(Res_imm[23]));
   NOR2_X1 i_373 (.A1(n_1763), .A2(n_1584), .ZN(n_1582));
   XOR2_X1 i_374 (.A(n_1605), .B(n_1593), .Z(Res_imm[25]));
   XOR2_X1 i_375 (.A(n_1592), .B(n_1589), .Z(Res_imm[26]));
   XOR2_X1 i_376 (.A(n_1590), .B(n_1587), .Z(Res_imm[27]));
   NOR2_X1 i_377 (.A1(n_1748), .A2(n_1751), .ZN(n_1587));
   XNOR2_X1 i_378 (.A(n_1594), .B(n_1588), .ZN(Res_imm[28]));
   OAI21_X1 i_379 (.A(n_1747), .B1(n_1751), .B2(n_1590), .ZN(n_1588));
   NOR2_X1 i_380 (.A1(n_1750), .A2(n_1689), .ZN(n_1589));
   INV_X1 i_381 (.A(n_1591), .ZN(n_1590));
   OAI21_X1 i_382 (.A(n_1749), .B1(n_1689), .B2(n_1592), .ZN(n_1591));
   AOI21_X1 i_383 (.A(n_764), .B1(n_760), .B2(n_1605), .ZN(n_1592));
   OAI21_X1 i_384 (.A(n_760), .B1(n_921), .B2(n_590), .ZN(n_1593));
   AOI21_X1 i_385 (.A(n_769), .B1(n_1713), .B2(n_1708), .ZN(n_1594));
   XNOR2_X1 i_386 (.A(n_1604), .B(n_1603), .ZN(Res_imm[29]));
   INV_X1 i_387 (.A(n_1595), .ZN(Res_imm[30]));
   AOI21_X1 i_388 (.A(n_1599), .B1(n_1601), .B2(n_1600), .ZN(n_1595));
   XOR2_X1 i_389 (.A(n_1597), .B(n_1596), .Z(Res_imm[31]));
   OAI21_X1 i_390 (.A(n_1756), .B1(n_1744), .B2(n_1601), .ZN(n_1596));
   OAI21_X1 i_391 (.A(n_1752), .B1(n_1707), .B2(n_1704), .ZN(n_1597));
   XNOR2_X1 i_392 (.A(n_1609), .B(n_1598), .ZN(Res_imm[32]));
   OAI21_X1 i_393 (.A(n_1752), .B1(n_770), .B2(n_1599), .ZN(n_1598));
   NOR2_X1 i_394 (.A1(n_1601), .A2(n_1600), .ZN(n_1599));
   OR2_X1 i_395 (.A1(n_1757), .A2(n_1744), .ZN(n_1600));
   INV_X1 i_396 (.A(n_1602), .ZN(n_1601));
   OAI22_X1 i_397 (.A1(n_1709), .A2(n_1710), .B1(n_1775), .B2(n_1604), .ZN(
      n_1602));
   OAI21_X1 i_398 (.A(n_761), .B1(n_1709), .B2(n_1710), .ZN(n_1603));
   OAI21_X1 i_399 (.A(n_1745), .B1(n_1742), .B2(n_1605), .ZN(n_1604));
   INV_X1 i_400 (.A(n_1606), .ZN(n_1605));
   OAI21_X1 i_401 (.A(n_1740), .B1(n_1738), .B2(n_1607), .ZN(n_1606));
   INV_X1 i_402 (.A(n_977), .ZN(n_1607));
   OAI22_X1 i_403 (.A1(n_1705), .A2(n_1701), .B1(n_1777), .B2(n_1778), .ZN(
      n_1609));
   XOR2_X1 i_404 (.A(n_1729), .B(n_1616), .Z(Res_imm[33]));
   XOR2_X1 i_405 (.A(n_1615), .B(n_1612), .Z(Res_imm[34]));
   XOR2_X1 i_406 (.A(n_1613), .B(n_1610), .Z(Res_imm[35]));
   NOR2_X1 i_407 (.A1(n_1759), .A2(n_1671), .ZN(n_1610));
   XNOR2_X1 i_408 (.A(n_1617), .B(n_1611), .ZN(Res_imm[36]));
   OAI22_X1 i_409 (.A1(n_1697), .A2(n_1695), .B1(n_1671), .B2(n_1613), .ZN(
      n_1611));
   AOI21_X1 i_410 (.A(n_1758), .B1(n_1699), .B2(n_1696), .ZN(n_1612));
   AOI21_X1 i_411 (.A(n_1758), .B1(n_1754), .B2(n_1614), .ZN(n_1613));
   INV_X1 i_412 (.A(n_1615), .ZN(n_1614));
   AOI21_X1 i_413 (.A(n_1753), .B1(n_1729), .B2(n_1755), .ZN(n_1615));
   OAI21_X1 i_414 (.A(n_1755), .B1(n_1703), .B2(n_1698), .ZN(n_1616));
   NOR2_X1 i_415 (.A1(n_1761), .A2(n_1762), .ZN(n_1617));
   XOR2_X1 i_416 (.A(n_1720), .B(n_1624), .Z(Res_imm[37]));
   XOR2_X1 i_417 (.A(n_1718), .B(n_1620), .Z(Res_imm[38]));
   XOR2_X1 i_418 (.A(n_1716), .B(n_1618), .Z(Res_imm[39]));
   NOR2_X1 i_419 (.A1(n_1791), .A2(n_1770), .ZN(n_1618));
   AOI21_X1 i_420 (.A(n_1769), .B1(n_1693), .B2(n_1686), .ZN(n_1620));
   OAI21_X1 i_421 (.A(n_1719), .B1(n_1694), .B2(n_1692), .ZN(n_1624));
   XOR2_X1 i_422 (.A(n_1804), .B(n_1810), .Z(Res_imm[42]));
   XNOR2_X1 i_423 (.A(n_1627), .B(n_1626), .ZN(Res_imm[43]));
   OAI22_X1 i_424 (.A1(n_1784), .A2(n_1796), .B1(n_1806), .B2(n_1804), .ZN(
      n_1626));
   NOR2_X1 i_425 (.A1(n_1800), .A2(n_1811), .ZN(n_1627));
   XNOR2_X1 i_426 (.A(n_1637), .B(n_1635), .ZN(Res_imm[46]));
   OAI21_X1 i_427 (.A(n_1765), .B1(n_1654), .B2(n_1767), .ZN(n_1635));
   OAI21_X1 i_428 (.A(n_1636), .B1(n_1654), .B2(n_1767), .ZN(Res_imm[47]));
   NAND2_X1 i_429 (.A1(n_1765), .A2(n_1637), .ZN(n_1636));
   AOI21_X1 i_430 (.A(n_1638), .B1(n_1819), .B2(n_1821), .ZN(n_1637));
   AOI21_X1 i_431 (.A(n_1815), .B1(n_1795), .B2(n_1812), .ZN(n_1638));
   INV_X1 i_432 (.A(n_1760), .ZN(n_1671));
   INV_X1 i_433 (.A(n_758), .ZN(n_1689));
   NAND2_X1 i_434 (.A1(n_591), .A2(n_630), .ZN(n_758));
   NAND2_X1 i_435 (.A1(n_921), .A2(n_590), .ZN(n_760));
   NAND2_X1 i_436 (.A1(n_1709), .A2(n_1710), .ZN(n_761));
   OAI21_X1 i_437 (.A(n_771), .B1(n_1513), .B2(n_1702), .ZN(n_762));
   INV_X1 i_438 (.A(n_1569), .ZN(n_1702));
   OAI222_X1 i_439 (.A1(n_954), .A2(n_955), .B1(n_2), .B2(n_4), .C1(n_1724), 
      .C2(n_1721), .ZN(n_763));
   AOI211_X1 i_440 (.A(n_1655), .B(n_1722), .C1(n_1629), .C2(n_1773), .ZN(n_1721));
   AOI22_X1 i_441 (.A1(A_imm[2]), .A2(n_0), .B1(A_imm[0]), .B2(n_1723), .ZN(
      n_1722));
   NOR2_X1 i_442 (.A1(n_1656), .A2(n_1628), .ZN(n_1723));
   AND2_X1 i_443 (.A1(n_2), .A2(n_4), .ZN(n_1724));
   NOR2_X1 i_444 (.A1(n_921), .A2(n_590), .ZN(n_764));
   NAND3_X1 i_445 (.A1(n_1776), .A2(n_1747), .A3(n_1749), .ZN(n_768));
   INV_X1 i_446 (.A(n_1748), .ZN(n_1747));
   NOR2_X1 i_447 (.A1(n_168), .A2(n_1712), .ZN(n_1748));
   INV_X1 i_448 (.A(n_1750), .ZN(n_1749));
   NOR2_X1 i_449 (.A1(n_591), .A2(n_630), .ZN(n_1750));
   NOR2_X1 i_450 (.A1(n_1713), .A2(n_1708), .ZN(n_769));
   OAI21_X1 i_451 (.A(n_1756), .B1(n_1707), .B2(n_1704), .ZN(n_770));
   INV_X1 i_452 (.A(n_1757), .ZN(n_1756));
   NOR2_X1 i_453 (.A1(n_1711), .A2(n_1706), .ZN(n_1757));
   NOR3_X1 i_454 (.A1(n_1763), .A2(n_1586), .A3(n_1583), .ZN(n_771));
   NOR2_X1 i_455 (.A1(n_938), .A2(n_773), .ZN(n_1763));
   NAND2_X1 i_456 (.A1(n_1654), .A2(n_1767), .ZN(n_1765));
   INV_X1 i_457 (.A(n_1813), .ZN(n_1767));
   INV_X1 i_458 (.A(n_0), .ZN(n_1773));
   FA_X1 i_459 (.A(n_1451), .B(n_1474), .CI(n_1497), .CO(n_353), .S(n_352));
   FA_X1 i_460 (.A(n_1382), .B(n_1405), .CI(n_1428), .CO(n_351), .S(n_350));
   FA_X1 i_461 (.A(n_1313), .B(n_1336), .CI(n_1359), .CO(n_349), .S(n_348));
   FA_X1 i_462 (.A(n_352), .B(n_350), .CI(n_348), .CO(n_363), .S(n_362));
   FA_X1 i_463 (.A(n_1430), .B(n_1453), .CI(n_1476), .CO(n_281), .S(n_280));
   FA_X1 i_464 (.A(n_1361), .B(n_1384), .CI(n_1407), .CO(n_279), .S(n_278));
   FA_X1 i_465 (.A(n_1292), .B(n_1315), .CI(n_1338), .CO(n_277), .S(n_276));
   FA_X1 i_466 (.A(n_281), .B(n_279), .CI(n_277), .CO(n_321), .S(n_320));
   FA_X1 i_467 (.A(n_1499), .B(n_1522), .CI(n_1545), .CO(n_283), .S(n_282));
   FA_X1 i_468 (.A(n_1544), .B(n_1565), .CI(n_283), .CO(n_319), .S(n_318));
   FA_X1 i_469 (.A(n_1520), .B(n_1543), .CI(n_1564), .CO(n_355), .S(n_354));
   FA_X1 i_470 (.A(n_321), .B(n_319), .CI(n_354), .CO(n_361), .S(n_360));
   FA_X1 i_471 (.A(n_1223), .B(n_1246), .CI(n_1269), .CO(n_275), .S(n_274));
   FA_X1 i_472 (.A(n_1154), .B(n_1177), .CI(n_1200), .CO(n_273), .S(n_272));
   FA_X1 i_473 (.A(n_1385), .B(n_1408), .CI(n_1431), .CO(n_247), .S(n_246));
   FA_X1 i_474 (.A(n_1316), .B(n_1339), .CI(n_1362), .CO(n_245), .S(n_244));
   FA_X1 i_475 (.A(n_1247), .B(n_1270), .CI(n_1293), .CO(n_243), .S(n_242));
   FA_X1 i_476 (.A(n_247), .B(n_245), .CI(n_243), .CO(n_287), .S(n_286));
   FA_X1 i_477 (.A(n_275), .B(n_273), .CI(n_287), .CO(n_323), .S(n_322));
   FA_X1 i_478 (.A(n_1268), .B(n_1291), .CI(n_1314), .CO(n_311), .S(n_310));
   FA_X1 i_479 (.A(n_1199), .B(n_1222), .CI(n_1245), .CO(n_309), .S(n_308));
   FA_X1 i_480 (.A(n_1130), .B(n_1153), .CI(n_1176), .CO(n_307), .S(n_306));
   FA_X1 i_481 (.A(n_311), .B(n_309), .CI(n_307), .CO(n_359), .S(n_358));
   FA_X1 i_482 (.A(n_1475), .B(n_1498), .CI(n_1521), .CO(n_317), .S(n_316));
   FA_X1 i_483 (.A(n_1406), .B(n_1429), .CI(n_1452), .CO(n_315), .S(n_314));
   FA_X1 i_484 (.A(n_1337), .B(n_1360), .CI(n_1383), .CO(n_313), .S(n_312));
   FA_X1 i_485 (.A(n_317), .B(n_315), .CI(n_313), .CO(n_357), .S(n_356));
   FA_X1 i_486 (.A(n_323), .B(n_358), .CI(n_356), .CO(n_367), .S(n_366));
   FA_X1 i_487 (.A(n_363), .B(n_361), .CI(n_367), .CO(n_409), .S(n_408));
   FA_X1 i_488 (.A(n_1427), .B(n_1450), .CI(n_1473), .CO(n_391), .S(n_390));
   FA_X1 i_489 (.A(n_1358), .B(n_1381), .CI(n_1404), .CO(n_389), .S(n_388));
   FA_X1 i_490 (.A(n_1289), .B(n_1312), .CI(n_1335), .CO(n_387), .S(n_386));
   FA_X1 i_491 (.A(n_391), .B(n_389), .CI(n_387), .CO(n_437), .S(n_436));
   FA_X1 i_492 (.A(n_1220), .B(n_1243), .CI(n_1266), .CO(n_385), .S(n_384));
   FA_X1 i_493 (.A(n_388), .B(n_386), .CI(n_384), .CO(n_403), .S(n_402));
   FA_X1 i_494 (.A(n_1496), .B(n_1519), .CI(n_1542), .CO(n_393), .S(n_392));
   FA_X1 i_495 (.A(n_357), .B(n_392), .CI(n_390), .CO(n_401), .S(n_400));
   FA_X1 i_496 (.A(n_436), .B(n_403), .CI(n_401), .CO(n_449), .S(n_448));
   FA_X1 i_497 (.A(n_1151), .B(n_1174), .CI(n_1197), .CO(n_383), .S(n_382));
   FA_X1 i_498 (.A(n_1082), .B(n_1105), .CI(n_1128), .CO(n_381), .S(n_380));
   FA_X1 i_499 (.A(n_1175), .B(n_1198), .CI(n_1221), .CO(n_345), .S(n_344));
   FA_X1 i_500 (.A(n_1106), .B(n_1129), .CI(n_1152), .CO(n_343), .S(n_342));
   FA_X1 i_501 (.A(n_345), .B(n_343), .CI(n_359), .CO(n_399), .S(n_398));
   FA_X1 i_502 (.A(n_382), .B(n_380), .CI(n_398), .CO(n_405), .S(n_404));
   FA_X1 i_503 (.A(n_404), .B(n_402), .CI(n_400), .CO(n_411), .S(n_410));
   FA_X1 i_504 (.A(n_409), .B(n_448), .CI(n_411), .CO(n_455), .S(n_454));
   FA_X1 i_505 (.A(n_280), .B(n_278), .CI(n_276), .CO(n_291), .S(n_290));
   FA_X1 i_506 (.A(n_1178), .B(n_1201), .CI(n_1224), .CO(n_241), .S(n_240));
   FA_X1 i_507 (.A(n_1478), .B(n_1501), .CI(n_1524), .CO(n_219), .S(n_218));
   FA_X1 i_508 (.A(n_1409), .B(n_1432), .CI(n_1455), .CO(n_217), .S(n_216));
   FA_X1 i_509 (.A(n_1340), .B(n_1363), .CI(n_1386), .CO(n_215), .S(n_214));
   FA_X1 i_510 (.A(n_219), .B(n_217), .CI(n_215), .CO(n_253), .S(n_252));
   FA_X1 i_511 (.A(n_241), .B(n_253), .CI(n_282), .CO(n_289), .S(n_288));
   FA_X1 i_512 (.A(n_320), .B(n_291), .CI(n_289), .CO(n_331), .S(n_330));
   FA_X1 i_513 (.A(n_308), .B(n_306), .CI(n_322), .CO(n_329), .S(n_328));
   FA_X1 i_514 (.A(n_1244), .B(n_1267), .CI(n_1290), .CO(n_347), .S(n_346));
   FA_X1 i_515 (.A(n_346), .B(n_344), .CI(n_342), .CO(n_365), .S(n_364));
   FA_X1 i_516 (.A(n_331), .B(n_329), .CI(n_364), .CO(n_371), .S(n_370));
   FA_X1 i_517 (.A(n_314), .B(n_312), .CI(n_310), .CO(n_327), .S(n_326));
   FA_X1 i_518 (.A(n_1523), .B(n_1546), .CI(n_1567), .CO(n_251), .S(n_250));
   FA_X1 i_519 (.A(n_1454), .B(n_1477), .CI(n_1500), .CO(n_249), .S(n_248));
   FA_X1 i_520 (.A(n_1566), .B(n_251), .CI(n_249), .CO(n_285), .S(n_284));
   FA_X1 i_521 (.A(n_285), .B(n_318), .CI(n_316), .CO(n_325), .S(n_324));
   FA_X1 i_522 (.A(n_327), .B(n_325), .CI(n_360), .CO(n_369), .S(n_368));
   FA_X1 i_523 (.A(n_362), .B(n_368), .CI(n_366), .CO(n_373), .S(n_372));
   FA_X1 i_524 (.A(n_371), .B(n_373), .CI(n_410), .CO(n_415), .S(n_414));
   FA_X1 i_525 (.A(n_351), .B(n_349), .CI(n_347), .CO(n_397), .S(n_396));
   FA_X1 i_526 (.A(n_1563), .B(n_355), .CI(n_353), .CO(n_395), .S(n_394));
   FA_X1 i_527 (.A(n_1541), .B(n_1562), .CI(n_393), .CO(n_435), .S(n_434));
   FA_X1 i_528 (.A(n_397), .B(n_395), .CI(n_434), .CO(n_441), .S(n_440));
   FA_X1 i_529 (.A(n_396), .B(n_394), .CI(n_365), .CO(n_407), .S(n_406));
   FA_X1 i_530 (.A(n_440), .B(n_407), .CI(n_405), .CO(n_451), .S(n_450));
   FA_X1 i_531 (.A(n_369), .B(n_408), .CI(n_406), .CO(n_413), .S(n_412));
   FA_X1 i_532 (.A(n_1265), .B(n_1288), .CI(n_1311), .CO(n_427), .S(n_426));
   FA_X1 i_533 (.A(n_1196), .B(n_1219), .CI(n_1242), .CO(n_425), .S(n_424));
   FA_X1 i_534 (.A(n_1127), .B(n_1150), .CI(n_1173), .CO(n_423), .S(n_422));
   FA_X1 i_535 (.A(n_426), .B(n_424), .CI(n_422), .CO(n_445), .S(n_444));
   FA_X1 i_536 (.A(n_1472), .B(n_1495), .CI(n_1518), .CO(n_433), .S(n_432));
   FA_X1 i_537 (.A(n_1403), .B(n_1426), .CI(n_1449), .CO(n_431), .S(n_430));
   FA_X1 i_538 (.A(n_1334), .B(n_1357), .CI(n_1380), .CO(n_429), .S(n_428));
   FA_X1 i_539 (.A(n_432), .B(n_430), .CI(n_428), .CO(n_443), .S(n_442));
   FA_X1 i_540 (.A(n_1058), .B(n_1081), .CI(n_1104), .CO(n_421), .S(n_420));
   FA_X1 i_541 (.A(n_385), .B(n_383), .CI(n_381), .CO(n_439), .S(n_438));
   FA_X1 i_542 (.A(n_420), .B(n_399), .CI(n_438), .CO(n_447), .S(n_446));
   FA_X1 i_543 (.A(n_444), .B(n_442), .CI(n_446), .CO(n_453), .S(n_452));
   FA_X1 i_544 (.A(n_450), .B(n_413), .CI(n_452), .CO(n_457), .S(n_456));
   FA_X1 i_545 (.A(n_454), .B(n_415), .CI(n_456), .CO(n_459), .S(n_458));
   FA_X1 i_546 (.A(n_421), .B(n_439), .CI(n_437), .CO(n_483), .S(n_482));
   FA_X1 i_547 (.A(n_443), .B(n_441), .CI(n_482), .CO(n_493), .S(n_492));
   FA_X1 i_548 (.A(n_427), .B(n_425), .CI(n_423), .CO(n_481), .S(n_480));
   FA_X1 i_549 (.A(n_433), .B(n_431), .CI(n_429), .CO(n_479), .S(n_478));
   FA_X1 i_550 (.A(n_480), .B(n_478), .CI(n_445), .CO(n_491), .S(n_490));
   FA_X1 i_551 (.A(n_492), .B(n_490), .CI(n_453), .CO(n_499), .S(n_498));
   FA_X1 i_552 (.A(n_1172), .B(n_1195), .CI(n_1218), .CO(n_467), .S(n_466));
   FA_X1 i_553 (.A(n_1103), .B(n_1126), .CI(n_1149), .CO(n_465), .S(n_464));
   FA_X1 i_554 (.A(n_1034), .B(n_1057), .CI(n_1080), .CO(n_463), .S(n_462));
   FA_X1 i_555 (.A(n_466), .B(n_464), .CI(n_462), .CO(n_489), .S(n_488));
   FA_X1 i_556 (.A(n_449), .B(n_447), .CI(n_488), .CO(n_495), .S(n_494));
   FA_X1 i_557 (.A(n_1379), .B(n_1402), .CI(n_1425), .CO(n_473), .S(n_472));
   FA_X1 i_558 (.A(n_1310), .B(n_1333), .CI(n_1356), .CO(n_471), .S(n_470));
   FA_X1 i_559 (.A(n_1241), .B(n_1264), .CI(n_1287), .CO(n_469), .S(n_468));
   FA_X1 i_560 (.A(n_472), .B(n_470), .CI(n_468), .CO(n_487), .S(n_486));
   FA_X1 i_561 (.A(n_1517), .B(n_1540), .CI(n_1561), .CO(n_477), .S(n_476));
   FA_X1 i_562 (.A(n_1448), .B(n_1471), .CI(n_1494), .CO(n_475), .S(n_474));
   FA_X1 i_563 (.A(n_435), .B(n_476), .CI(n_474), .CO(n_485), .S(n_484));
   FA_X1 i_564 (.A(n_486), .B(n_484), .CI(n_451), .CO(n_497), .S(n_496));
   FA_X1 i_565 (.A(n_494), .B(n_455), .CI(n_496), .CO(n_501), .S(n_500));
   FA_X1 i_566 (.A(n_498), .B(n_457), .CI(n_500), .CO(n_503), .S(n_502));
   HA_X1 i_567 (.A(n_459), .B(n_502), .CO(n_775), .S(n_773));
   FA_X1 i_568 (.A(n_469), .B(n_467), .CI(n_465), .CO(n_776), .S(n_524));
   FA_X1 i_569 (.A(n_475), .B(n_473), .CI(n_471), .CO(n_778), .S(n_522));
   FA_X1 i_570 (.A(n_524), .B(n_522), .CI(n_489), .CO(n_780), .S(n_534));
   FA_X1 i_571 (.A(n_534), .B(n_495), .CI(n_497), .CO(n_783), .S(n_542));
   FA_X1 i_572 (.A(n_1102), .B(n_1125), .CI(n_1148), .CO(n_785), .S(n_508));
   FA_X1 i_573 (.A(n_1033), .B(n_1056), .CI(n_1079), .CO(n_786), .S(n_506));
   FA_X1 i_574 (.A(n_508), .B(n_506), .CI(n_483), .CO(n_787), .S(n_532));
   FA_X1 i_575 (.A(n_1309), .B(n_1332), .CI(n_1355), .CO(n_788), .S(n_514));
   FA_X1 i_576 (.A(n_1240), .B(n_1263), .CI(n_1286), .CO(n_789), .S(n_512));
   FA_X1 i_577 (.A(n_1171), .B(n_1194), .CI(n_1217), .CO(n_790), .S(n_510));
   FA_X1 i_578 (.A(n_514), .B(n_512), .CI(n_510), .CO(n_791), .S(n_530));
   FA_X1 i_579 (.A(n_491), .B(n_532), .CI(n_530), .CO(n_792), .S(n_538));
   FA_X1 i_580 (.A(n_1516), .B(n_1539), .CI(n_477), .CO(n_793), .S(n_520));
   FA_X1 i_581 (.A(n_1447), .B(n_1470), .CI(n_1493), .CO(n_800), .S(n_518));
   FA_X1 i_582 (.A(n_1378), .B(n_1401), .CI(n_1424), .CO(n_801), .S(n_516));
   FA_X1 i_583 (.A(n_520), .B(n_518), .CI(n_516), .CO(n_828), .S(n_528));
   FA_X1 i_584 (.A(n_463), .B(n_481), .CI(n_479), .CO(n_829), .S(n_526));
   FA_X1 i_585 (.A(n_487), .B(n_485), .CI(n_526), .CO(n_854), .S(n_536));
   FA_X1 i_586 (.A(n_528), .B(n_493), .CI(n_536), .CO(n_855), .S(n_540));
   FA_X1 i_587 (.A(n_499), .B(n_538), .CI(n_540), .CO(n_878), .S(n_544));
   FA_X1 i_588 (.A(n_542), .B(n_501), .CI(n_544), .CO(n_879), .S(n_546));
   HA_X1 i_589 (.A(n_503), .B(n_546), .CO(n_921), .S(n_900));
   FA_X1 i_590 (.A(n_1271), .B(n_1294), .CI(n_1317), .CO(n_213), .S(n_212));
   FA_X1 i_591 (.A(n_1202), .B(n_1225), .CI(n_1248), .CO(n_211), .S(n_210));
   FA_X1 i_592 (.A(n_1433), .B(n_1456), .CI(n_1479), .CO(n_189), .S(n_188));
   FA_X1 i_593 (.A(n_1364), .B(n_1387), .CI(n_1410), .CO(n_187), .S(n_186));
   FA_X1 i_594 (.A(n_1295), .B(n_1318), .CI(n_1341), .CO(n_185), .S(n_184));
   FA_X1 i_595 (.A(n_189), .B(n_187), .CI(n_185), .CO(n_223), .S(n_222));
   FA_X1 i_596 (.A(n_213), .B(n_211), .CI(n_223), .CO(n_255), .S(n_254));
   FA_X1 i_597 (.A(n_274), .B(n_272), .CI(n_255), .CO(n_293), .S(n_292));
   FA_X1 i_598 (.A(n_246), .B(n_244), .CI(n_242), .CO(n_259), .S(n_258));
   FA_X1 i_599 (.A(n_286), .B(n_284), .CI(n_259), .CO(n_295), .S(n_294));
   FA_X1 i_600 (.A(n_293), .B(n_295), .CI(n_328), .CO(n_333), .S(n_332));
   FA_X1 i_601 (.A(n_1502), .B(n_1525), .CI(n_1548), .CO(n_191), .S(n_190));
   FA_X1 i_602 (.A(n_1547), .B(n_1568), .CI(n_191), .CO(n_221), .S(n_220));
   FA_X1 i_603 (.A(n_221), .B(n_250), .CI(n_248), .CO(n_257), .S(n_256));
   FA_X1 i_604 (.A(n_214), .B(n_212), .CI(n_210), .CO(n_229), .S(n_228));
   FA_X1 i_605 (.A(n_220), .B(n_218), .CI(n_216), .CO(n_227), .S(n_226));
   FA_X1 i_606 (.A(n_252), .B(n_229), .CI(n_227), .CO(n_263), .S(n_262));
   FA_X1 i_607 (.A(n_257), .B(n_288), .CI(n_263), .CO(n_297), .S(n_296));
   FA_X1 i_608 (.A(n_326), .B(n_324), .CI(n_297), .CO(n_335), .S(n_334));
   FA_X1 i_609 (.A(n_333), .B(n_335), .CI(n_370), .CO(n_375), .S(n_374));
   FA_X1 i_610 (.A(n_375), .B(n_412), .CI(n_414), .CO(n_417), .S(n_416));
   HA_X1 i_611 (.A(n_417), .B(n_458), .CO(n_938), .S(n_460));
   FA_X1 i_612 (.A(n_700), .B(n_703), .CI(n_705), .CO(n_183), .S(n_182));
   FA_X1 i_613 (.A(n_158), .B(n_156), .CI(n_140), .CO(n_195), .S(n_194));
   FA_X1 i_614 (.A(n_756), .B(n_162), .CI(n_160), .CO(n_193), .S(n_192));
   FA_X1 i_615 (.A(n_183), .B(n_195), .CI(n_193), .CO(n_225), .S(n_224));
   FA_X1 i_616 (.A(n_240), .B(n_225), .CI(n_254), .CO(n_261), .S(n_260));
   FA_X1 i_617 (.A(n_261), .B(n_292), .CI(n_290), .CO(n_299), .S(n_298));
   FA_X1 i_618 (.A(n_330), .B(n_299), .CI(n_332), .CO(n_337), .S(n_336));
   FA_X1 i_619 (.A(n_337), .B(n_372), .CI(n_374), .CO(n_377), .S(n_376));
   HA_X1 i_620 (.A(n_377), .B(n_416), .CO(n_419), .S(n_418));
   FA_X1 i_621 (.A(n_222), .B(n_199), .CI(n_197), .CO(n_231), .S(n_230));
   FA_X1 i_622 (.A(n_231), .B(n_258), .CI(n_256), .CO(n_265), .S(n_264));
   FA_X1 i_623 (.A(n_294), .B(n_265), .CI(n_296), .CO(n_301), .S(n_300));
   FA_X1 i_624 (.A(n_334), .B(n_301), .CI(n_336), .CO(n_339), .S(n_338));
   FA_X1 i_625 (.A(n_224), .B(n_201), .CI(n_228), .CO(n_233), .S(n_232));
   FA_X1 i_626 (.A(n_260), .B(n_262), .CI(n_233), .CO(n_267), .S(n_266));
   FA_X1 i_627 (.A(n_267), .B(n_298), .CI(n_300), .CO(n_303), .S(n_302));
   HA_X1 i_628 (.A(n_303), .B(n_338), .CO(n_341), .S(n_340));
   HA_X1 i_629 (.A(n_339), .B(n_341), .CO(n_379), .S(n_378));
   FA_X1 i_630 (.A(n_226), .B(n_230), .CI(n_203), .CO(n_235), .S(n_234));
   FA_X1 i_631 (.A(n_235), .B(n_264), .CI(n_266), .CO(n_269), .S(n_268));
   HA_X1 i_632 (.A(n_269), .B(n_302), .CO(n_305), .S(n_304));
   FA_X1 i_633 (.A(n_196), .B(n_175), .CI(n_200), .CO(n_205), .S(n_204));
   FA_X1 i_634 (.A(n_232), .B(n_205), .CI(n_234), .CO(n_237), .S(n_236));
   FA_X1 i_635 (.A(n_177), .B(n_202), .CI(n_204), .CO(n_207), .S(n_206));
   HA_X1 i_636 (.A(n_179), .B(n_181), .CO(n_209), .S(n_208));
   HA_X1 i_637 (.A(n_207), .B(n_209), .CO(n_239), .S(n_238));
   HA_X1 i_638 (.A(n_237), .B(n_239), .CO(n_271), .S(n_270));
   FA_X1 i_639 (.A(n_121), .B(n_142), .CI(n_123), .CO(n_149), .S(n_148));
   FA_X1 i_640 (.A(n_143), .B(n_138), .CI(n_163), .CO(n_173), .S(n_172));
   FA_X1 i_641 (.A(n_161), .B(n_159), .CI(n_157), .CO(n_171), .S(n_170));
   FA_X1 i_642 (.A(n_149), .B(n_172), .CI(n_170), .CO(n_177), .S(n_176));
   FA_X1 i_643 (.A(n_186), .B(n_184), .CI(n_182), .CO(n_199), .S(n_198));
   FA_X1 i_644 (.A(n_171), .B(n_173), .CI(n_198), .CO(n_203), .S(n_202));
   FA_X1 i_645 (.A(n_164), .B(n_190), .CI(n_188), .CO(n_197), .S(n_196));
   FA_X1 i_646 (.A(n_147), .B(n_145), .CI(n_165), .CO(n_175), .S(n_174));
   FA_X1 i_647 (.A(n_166), .B(n_194), .CI(n_192), .CO(n_201), .S(n_200));
   FA_X1 i_648 (.A(n_125), .B(n_146), .CI(n_144), .CO(n_151), .S(n_150));
   FA_X1 i_649 (.A(n_174), .B(n_151), .CI(n_176), .CO(n_179), .S(n_178));
   FA_X1 i_650 (.A(n_148), .B(n_127), .CI(n_129), .CO(n_153), .S(n_152));
   HA_X1 i_651 (.A(n_150), .B(n_131), .CO(n_155), .S(n_154));
   HA_X1 i_652 (.A(n_153), .B(n_155), .CO(n_181), .S(n_180));
   FA_X1 i_653 (.A(n_91), .B(n_85), .CI(n_96), .CO(n_121), .S(n_120));
   FA_X1 i_654 (.A(n_113), .B(n_111), .CI(n_99), .CO(n_939), .S(n_142));
   FA_X1 i_655 (.A(n_114), .B(n_112), .CI(n_110), .CO(n_123), .S(n_122));
   FA_X1 i_656 (.A(n_66), .B(n_93), .CI(n_92), .CO(n_101), .S(n_100));
   FA_X1 i_657 (.A(n_90), .B(n_84), .CI(n_67), .CO(n_103), .S(n_102));
   FA_X1 i_658 (.A(n_101), .B(n_103), .CI(n_122), .CO(n_127), .S(n_126));
   FA_X1 i_659 (.A(n_94), .B(n_81), .CI(n_83), .CO(n_105), .S(n_104));
   FA_X1 i_660 (.A(n_98), .B(n_120), .CI(n_115), .CO(n_125), .S(n_124));
   FA_X1 i_661 (.A(n_105), .B(n_124), .CI(n_126), .CO(n_129), .S(n_128));
   FA_X1 i_662 (.A(n_132), .B(n_119), .CI(n_118), .CO(n_147), .S(n_146));
   FA_X1 i_663 (.A(n_116), .B(n_136), .CI(n_134), .CO(n_145), .S(n_144));
   FA_X1 i_664 (.A(n_102), .B(n_100), .CI(n_104), .CO(n_107), .S(n_106));
   HA_X1 i_665 (.A(n_89), .B(n_87), .CO(n_109), .S(n_108));
   HA_X1 i_666 (.A(n_107), .B(n_109), .CO(n_131), .S(n_130));
   FA_X1 i_667 (.A(n_64), .B(n_79), .CI(n_82), .CO(n_87), .S(n_86));
   HA_X1 i_668 (.A(n_71), .B(n_69), .CO(n_89), .S(n_88));
   FA_X1 i_669 (.A(n_48), .B(n_50), .CI(n_51), .CO(n_69), .S(n_68));
   HA_X1 i_670 (.A(n_55), .B(n_53), .CO(n_71), .S(n_70));
   FA_X1 i_671 (.A(n_24), .B(n_22), .CI(n_29), .CO(n_39), .S(n_38));
   HA_X1 i_672 (.A(n_30), .B(n_27), .CO(n_41), .S(n_40));
   FA_X1 i_673 (.A(n_36), .B(n_32), .CI(n_41), .CO(n_53), .S(n_52));
   HA_X1 i_674 (.A(n_39), .B(n_37), .CO(n_55), .S(n_54));
   FA_X1 i_675 (.A(n_14), .B(n_12), .CI(n_20), .CO(n_27), .S(n_26));
   HA_X1 i_676 (.A(n_19), .B(n_17), .CO(n_29), .S(n_28));
   FA_X1 i_677 (.A(n_7), .B(n_8), .CI(n_10), .CO(n_17), .S(n_16));
   HA_X1 i_678 (.A(n_9), .B(n_11), .CO(n_19), .S(n_18));
   FA_X1 i_679 (.A(n_737), .B(n_738), .CI(n_739), .CO(n_7), .S(n_954));
   HA_X1 i_680 (.A(n_3), .B(n_6), .CO(n_11), .S(n_955));
   NOR2_X1 i_681 (.A1(n_1656), .A2(n_1645), .ZN(n_1548));
   NOR2_X1 i_682 (.A1(n_1657), .A2(n_1644), .ZN(n_1525));
   NOR2_X1 i_683 (.A1(n_1658), .A2(n_1643), .ZN(n_1502));
   NOR2_X1 i_684 (.A1(n_1655), .A2(n_1647), .ZN(n_1568));
   NOR2_X1 i_685 (.A1(n_1656), .A2(n_1646), .ZN(n_1547));
   NOR2_X1 i_686 (.A1(n_1665), .A2(n_1632), .ZN(n_1341));
   NOR2_X1 i_687 (.A1(n_1666), .A2(n_1631), .ZN(n_1318));
   NOR2_X1 i_688 (.A1(n_1667), .A2(n_1630), .ZN(n_1295));
   NOR2_X1 i_689 (.A1(n_1662), .A2(n_1639), .ZN(n_1410));
   NOR2_X1 i_690 (.A1(n_1663), .A2(n_1634), .ZN(n_1387));
   NOR2_X1 i_691 (.A1(n_1664), .A2(n_1633), .ZN(n_1364));
   NOR2_X1 i_692 (.A1(n_1659), .A2(n_1642), .ZN(n_1479));
   NOR2_X1 i_693 (.A1(n_1660), .A2(n_1641), .ZN(n_1456));
   NOR2_X1 i_694 (.A1(n_1661), .A2(n_1640), .ZN(n_1433));
   NOR2_X1 i_695 (.A1(n_1669), .A2(n_1629), .ZN(n_1248));
   NOR2_X1 i_696 (.A1(n_1670), .A2(n_1628), .ZN(n_1225));
   NOR2_X1 i_697 (.A1(n_1672), .A2(n_1625), .ZN(n_1202));
   NOR2_X1 i_698 (.A1(n_1666), .A2(n_1632), .ZN(n_1317));
   NOR2_X1 i_699 (.A1(n_1667), .A2(n_1631), .ZN(n_1294));
   NOR2_X1 i_700 (.A1(n_1668), .A2(n_1630), .ZN(n_1271));
   NOR2_X1 i_701 (.A1(n_1661), .A2(n_1649), .ZN(n_1424));
   NOR2_X1 i_702 (.A1(n_1662), .A2(n_1648), .ZN(n_1401));
   NOR2_X1 i_703 (.A1(n_1663), .A2(n_1647), .ZN(n_1378));
   NOR2_X1 i_704 (.A1(n_1658), .A2(n_1652), .ZN(n_1493));
   NOR2_X1 i_705 (.A1(n_1659), .A2(n_1651), .ZN(n_1470));
   NOR2_X1 i_706 (.A1(n_1660), .A2(n_1650), .ZN(n_1447));
   NOR2_X1 i_707 (.A1(n_1656), .A2(n_1654), .ZN(n_1539));
   NOR2_X1 i_708 (.A1(n_1657), .A2(n_1653), .ZN(n_1516));
   NOR2_X1 i_709 (.A1(n_1670), .A2(n_1640), .ZN(n_1217));
   NOR2_X1 i_710 (.A1(n_1672), .A2(n_1639), .ZN(n_1194));
   NOR2_X1 i_711 (.A1(n_1673), .A2(n_1634), .ZN(n_1171));
   NOR2_X1 i_712 (.A1(n_1667), .A2(n_1643), .ZN(n_1286));
   NOR2_X1 i_713 (.A1(n_1668), .A2(n_1642), .ZN(n_1263));
   NOR2_X1 i_714 (.A1(n_1669), .A2(n_1641), .ZN(n_1240));
   NOR2_X1 i_715 (.A1(n_1664), .A2(n_1646), .ZN(n_1355));
   NOR2_X1 i_716 (.A1(n_1665), .A2(n_1645), .ZN(n_1332));
   NOR2_X1 i_717 (.A1(n_1666), .A2(n_1644), .ZN(n_1309));
   NOR2_X1 i_718 (.A1(n_1677), .A2(n_1630), .ZN(n_1079));
   NOR2_X1 i_719 (.A1(n_1678), .A2(n_1629), .ZN(n_1056));
   NOR2_X1 i_720 (.A1(n_1654), .A2(n_1628), .ZN(n_1033));
   NOR2_X1 i_721 (.A1(n_1674), .A2(n_1633), .ZN(n_1148));
   NOR2_X1 i_722 (.A1(n_1675), .A2(n_1632), .ZN(n_1125));
   NOR2_X1 i_723 (.A1(n_1676), .A2(n_1631), .ZN(n_1102));
   NOR2_X1 i_724 (.A1(n_1658), .A2(n_1651), .ZN(n_1494));
   NOR2_X1 i_725 (.A1(n_1659), .A2(n_1650), .ZN(n_1471));
   NOR2_X1 i_726 (.A1(n_1660), .A2(n_1649), .ZN(n_1448));
   NOR2_X1 i_727 (.A1(n_1655), .A2(n_1654), .ZN(n_1561));
   NOR2_X1 i_728 (.A1(n_1656), .A2(n_1653), .ZN(n_1540));
   NOR2_X1 i_729 (.A1(n_1657), .A2(n_1652), .ZN(n_1517));
   NOR2_X1 i_730 (.A1(n_1667), .A2(n_1642), .ZN(n_1287));
   NOR2_X1 i_731 (.A1(n_1668), .A2(n_1641), .ZN(n_1264));
   NOR2_X1 i_732 (.A1(n_1669), .A2(n_1640), .ZN(n_1241));
   NOR2_X1 i_733 (.A1(n_1664), .A2(n_1645), .ZN(n_1356));
   NOR2_X1 i_734 (.A1(n_1665), .A2(n_1644), .ZN(n_1333));
   NOR2_X1 i_735 (.A1(n_1666), .A2(n_1643), .ZN(n_1310));
   NOR2_X1 i_736 (.A1(n_1661), .A2(n_1648), .ZN(n_1425));
   NOR2_X1 i_737 (.A1(n_1662), .A2(n_1647), .ZN(n_1402));
   NOR2_X1 i_738 (.A1(n_1663), .A2(n_1646), .ZN(n_1379));
   NOR2_X1 i_739 (.A1(n_1677), .A2(n_1629), .ZN(n_1080));
   NOR2_X1 i_740 (.A1(n_1678), .A2(n_1628), .ZN(n_1057));
   NOR2_X1 i_741 (.A1(n_1654), .A2(n_1625), .ZN(n_1034));
   NOR2_X1 i_742 (.A1(n_1674), .A2(n_1632), .ZN(n_1149));
   NOR2_X1 i_743 (.A1(n_1675), .A2(n_1631), .ZN(n_1126));
   NOR2_X1 i_745 (.A1(n_1676), .A2(n_1630), .ZN(n_1103));
   NOR2_X1 i_746 (.A1(n_1670), .A2(n_1639), .ZN(n_1218));
   NOR2_X1 i_747 (.A1(n_1672), .A2(n_1634), .ZN(n_1195));
   NOR2_X1 i_748 (.A1(n_1673), .A2(n_1633), .ZN(n_1172));
   NOR2_X1 i_749 (.A1(n_1676), .A2(n_1629), .ZN(n_1104));
   NOR2_X1 i_750 (.A1(n_1677), .A2(n_1628), .ZN(n_1081));
   NOR2_X1 i_751 (.A1(n_1678), .A2(n_1625), .ZN(n_1058));
   NOR2_X1 i_752 (.A1(n_1663), .A2(n_1645), .ZN(n_1380));
   NOR2_X1 i_753 (.A1(n_1664), .A2(n_1644), .ZN(n_1357));
   NOR2_X1 i_754 (.A1(n_1665), .A2(n_1643), .ZN(n_1334));
   NOR2_X1 i_755 (.A1(n_1660), .A2(n_1648), .ZN(n_1449));
   NOR2_X1 i_756 (.A1(n_1661), .A2(n_1647), .ZN(n_1426));
   NOR2_X1 i_757 (.A1(n_1662), .A2(n_1646), .ZN(n_1403));
   NOR2_X1 i_758 (.A1(n_1657), .A2(n_1651), .ZN(n_1518));
   NOR2_X1 i_759 (.A1(n_1658), .A2(n_1650), .ZN(n_1495));
   NOR2_X1 i_760 (.A1(n_1659), .A2(n_1649), .ZN(n_1472));
   NOR2_X1 i_761 (.A1(n_1673), .A2(n_1632), .ZN(n_1173));
   NOR2_X1 i_762 (.A1(n_1674), .A2(n_1631), .ZN(n_1150));
   NOR2_X1 i_763 (.A1(n_1675), .A2(n_1630), .ZN(n_1127));
   NOR2_X1 i_764 (.A1(n_1669), .A2(n_1639), .ZN(n_1242));
   NOR2_X1 i_765 (.A1(n_1670), .A2(n_1634), .ZN(n_1219));
   NOR2_X1 i_766 (.A1(n_1672), .A2(n_1633), .ZN(n_1196));
   NOR2_X1 i_768 (.A1(n_1666), .A2(n_1642), .ZN(n_1311));
   NOR2_X1 i_769 (.A1(n_1667), .A2(n_1641), .ZN(n_1288));
   NOR2_X1 i_770 (.A1(n_1668), .A2(n_1640), .ZN(n_1265));
   NOR2_X1 i_771 (.A1(n_1655), .A2(n_1653), .ZN(n_1562));
   NOR2_X1 i_772 (.A1(n_1656), .A2(n_1652), .ZN(n_1541));
   NOR2_X1 i_773 (.A1(n_1655), .A2(n_1652), .ZN(n_1563));
   NOR2_X1 i_774 (.A1(n_1658), .A2(n_1645), .ZN(n_1500));
   NOR2_X1 i_775 (.A1(n_1659), .A2(n_1644), .ZN(n_1477));
   NOR2_X1 i_776 (.A1(n_1660), .A2(n_1643), .ZN(n_1454));
   NOR2_X1 i_777 (.A1(n_1655), .A2(n_1648), .ZN(n_1567));
   NOR2_X1 i_778 (.A1(n_1656), .A2(n_1647), .ZN(n_1546));
   NOR2_X1 i_779 (.A1(n_1657), .A2(n_1646), .ZN(n_1523));
   NOR2_X1 i_780 (.A1(n_1655), .A2(n_1649), .ZN(n_1566));
   NOR2_X1 i_781 (.A1(n_1667), .A2(n_1639), .ZN(n_1290));
   NOR2_X1 i_782 (.A1(n_1668), .A2(n_1634), .ZN(n_1267));
   NOR2_X1 i_783 (.A1(n_1669), .A2(n_1633), .ZN(n_1244));
   NOR2_X1 i_784 (.A1(n_1663), .A2(n_1639), .ZN(n_1386));
   NOR2_X1 i_785 (.A1(n_1664), .A2(n_1634), .ZN(n_1363));
   NOR2_X1 i_786 (.A1(n_1665), .A2(n_1633), .ZN(n_1340));
   NOR2_X1 i_787 (.A1(n_1660), .A2(n_1642), .ZN(n_1455));
   NOR2_X1 i_788 (.A1(n_1661), .A2(n_1641), .ZN(n_1432));
   NOR2_X1 i_789 (.A1(n_1662), .A2(n_1640), .ZN(n_1409));
   NOR2_X1 i_791 (.A1(n_1657), .A2(n_1645), .ZN(n_1524));
   NOR2_X1 i_793 (.A1(n_1658), .A2(n_1644), .ZN(n_1501));
   NOR2_X1 i_794 (.A1(n_1659), .A2(n_1643), .ZN(n_1478));
   NOR2_X1 i_795 (.A1(n_1670), .A2(n_1629), .ZN(n_1224));
   NOR2_X1 i_796 (.A1(n_1672), .A2(n_1628), .ZN(n_1201));
   NOR2_X1 i_797 (.A1(n_1673), .A2(n_1625), .ZN(n_1178));
   NOR2_X1 i_798 (.A1(n_1674), .A2(n_1629), .ZN(n_1152));
   NOR2_X1 i_799 (.A1(n_1675), .A2(n_1628), .ZN(n_1129));
   NOR2_X1 i_800 (.A1(n_1676), .A2(n_1625), .ZN(n_1106));
   NOR2_X1 i_801 (.A1(n_1670), .A2(n_1632), .ZN(n_1221));
   NOR2_X1 i_802 (.A1(n_1672), .A2(n_1631), .ZN(n_1198));
   NOR2_X1 i_803 (.A1(n_1673), .A2(n_1630), .ZN(n_1175));
   NOR2_X1 i_804 (.A1(n_1675), .A2(n_1629), .ZN(n_1128));
   NOR2_X1 i_805 (.A1(n_1676), .A2(n_1628), .ZN(n_1105));
   NOR2_X1 i_806 (.A1(n_1677), .A2(n_1625), .ZN(n_1082));
   NOR2_X1 i_807 (.A1(n_1672), .A2(n_1632), .ZN(n_1197));
   NOR2_X1 i_808 (.A1(n_1673), .A2(n_1631), .ZN(n_1174));
   NOR2_X1 i_809 (.A1(n_1674), .A2(n_1630), .ZN(n_1151));
   NOR2_X1 i_810 (.A1(n_1656), .A2(n_1651), .ZN(n_1542));
   NOR2_X1 i_811 (.A1(n_1657), .A2(n_1650), .ZN(n_1519));
   NOR2_X1 i_812 (.A1(n_1658), .A2(n_1649), .ZN(n_1496));
   NOR2_X1 i_814 (.A1(n_1668), .A2(n_1639), .ZN(n_1266));
   NOR2_X1 i_817 (.A1(n_1669), .A2(n_1634), .ZN(n_1243));
   NOR2_X1 i_818 (.A1(n_1670), .A2(n_1633), .ZN(n_1220));
   NOR2_X1 i_819 (.A1(n_1665), .A2(n_1642), .ZN(n_1335));
   NOR2_X1 i_820 (.A1(n_1666), .A2(n_1641), .ZN(n_1312));
   NOR2_X1 i_821 (.A1(n_1667), .A2(n_1640), .ZN(n_1289));
   NOR2_X1 i_822 (.A1(n_1662), .A2(n_1645), .ZN(n_1404));
   NOR2_X1 i_823 (.A1(n_1663), .A2(n_1644), .ZN(n_1381));
   NOR2_X1 i_824 (.A1(n_1664), .A2(n_1643), .ZN(n_1358));
   NOR2_X1 i_825 (.A1(n_1659), .A2(n_1648), .ZN(n_1473));
   NOR2_X1 i_826 (.A1(n_1660), .A2(n_1647), .ZN(n_1450));
   NOR2_X1 i_827 (.A1(n_1661), .A2(n_1646), .ZN(n_1427));
   NOR2_X1 i_828 (.A1(n_1663), .A2(n_1642), .ZN(n_1383));
   NOR2_X1 i_829 (.A1(n_1664), .A2(n_1641), .ZN(n_1360));
   NOR2_X1 i_830 (.A1(n_1665), .A2(n_1640), .ZN(n_1337));
   NOR2_X1 i_831 (.A1(n_1660), .A2(n_1645), .ZN(n_1452));
   NOR2_X1 i_832 (.A1(n_1661), .A2(n_1644), .ZN(n_1429));
   NOR2_X1 i_833 (.A1(n_1662), .A2(n_1643), .ZN(n_1406));
   NOR2_X1 i_834 (.A1(n_1657), .A2(n_1648), .ZN(n_1521));
   NOR2_X1 i_835 (.A1(n_1658), .A2(n_1647), .ZN(n_1498));
   NOR2_X1 i_840 (.A1(n_1659), .A2(n_1646), .ZN(n_1475));
   NOR2_X1 i_841 (.A1(n_1673), .A2(n_1629), .ZN(n_1176));
   NOR2_X1 i_842 (.A1(n_1674), .A2(n_1628), .ZN(n_1153));
   NOR2_X1 i_843 (.A1(n_1675), .A2(n_1625), .ZN(n_1130));
   NOR2_X1 i_844 (.A1(n_1669), .A2(n_1632), .ZN(n_1245));
   NOR2_X1 i_845 (.A1(n_1670), .A2(n_1631), .ZN(n_1222));
   NOR2_X1 i_846 (.A1(n_1672), .A2(n_1630), .ZN(n_1199));
   NOR2_X1 i_847 (.A1(n_1666), .A2(n_1639), .ZN(n_1314));
   NOR2_X1 i_848 (.A1(n_1667), .A2(n_1634), .ZN(n_1291));
   NOR2_X1 i_849 (.A1(n_1668), .A2(n_1633), .ZN(n_1268));
   NOR2_X1 i_850 (.A1(n_1667), .A2(n_1632), .ZN(n_1293));
   NOR2_X1 i_851 (.A1(n_1668), .A2(n_1631), .ZN(n_1270));
   NOR2_X1 i_852 (.A1(n_1669), .A2(n_1630), .ZN(n_1247));
   NOR2_X1 i_853 (.A1(n_1664), .A2(n_1639), .ZN(n_1362));
   NOR2_X1 i_854 (.A1(n_1665), .A2(n_1634), .ZN(n_1339));
   NOR2_X1 i_855 (.A1(n_1666), .A2(n_1633), .ZN(n_1316));
   NOR2_X1 i_856 (.A1(n_1661), .A2(n_1642), .ZN(n_1431));
   NOR2_X1 i_857 (.A1(n_1662), .A2(n_1641), .ZN(n_1408));
   NOR2_X1 i_858 (.A1(n_1663), .A2(n_1640), .ZN(n_1385));
   NOR2_X1 i_863 (.A1(n_1672), .A2(n_1629), .ZN(n_1200));
   NOR2_X1 i_864 (.A1(n_1673), .A2(n_1628), .ZN(n_1177));
   NOR2_X1 i_865 (.A1(n_1674), .A2(n_1625), .ZN(n_1154));
   NOR2_X1 i_866 (.A1(n_1668), .A2(n_1632), .ZN(n_1269));
   NOR2_X1 i_867 (.A1(n_1669), .A2(n_1631), .ZN(n_1246));
   NOR2_X1 i_868 (.A1(n_1670), .A2(n_1630), .ZN(n_1223));
   NOR2_X1 i_869 (.A1(n_1655), .A2(n_1651), .ZN(n_1564));
   NOR2_X1 i_870 (.A1(n_1656), .A2(n_1650), .ZN(n_1543));
   NOR2_X1 i_871 (.A1(n_1657), .A2(n_1649), .ZN(n_1520));
   NOR2_X1 i_872 (.A1(n_1656), .A2(n_1648), .ZN(n_1545));
   NOR2_X1 i_873 (.A1(n_1657), .A2(n_1647), .ZN(n_1522));
   NOR2_X1 i_874 (.A1(n_1658), .A2(n_1646), .ZN(n_1499));
   NOR2_X1 i_875 (.A1(n_1655), .A2(n_1650), .ZN(n_1565));
   NOR2_X1 i_876 (.A1(n_1656), .A2(n_1649), .ZN(n_1544));
   NOR2_X1 i_877 (.A1(n_1665), .A2(n_1639), .ZN(n_1338));
   NOR2_X1 i_878 (.A1(n_1666), .A2(n_1634), .ZN(n_1315));
   NOR2_X1 i_879 (.A1(n_1667), .A2(n_1633), .ZN(n_1292));
   NOR2_X1 i_880 (.A1(n_1662), .A2(n_1642), .ZN(n_1407));
   NOR2_X1 i_881 (.A1(n_1663), .A2(n_1641), .ZN(n_1384));
   NOR2_X1 i_886 (.A1(n_1664), .A2(n_1640), .ZN(n_1361));
   NOR2_X1 i_887 (.A1(n_1659), .A2(n_1645), .ZN(n_1476));
   NOR2_X1 i_888 (.A1(n_1660), .A2(n_1644), .ZN(n_1453));
   NOR2_X1 i_889 (.A1(n_1661), .A2(n_1643), .ZN(n_1430));
   NOR2_X1 i_890 (.A1(n_1664), .A2(n_1642), .ZN(n_1359));
   NOR2_X1 i_891 (.A1(n_1665), .A2(n_1641), .ZN(n_1336));
   NOR2_X1 i_892 (.A1(n_1666), .A2(n_1640), .ZN(n_1313));
   NOR2_X1 i_893 (.A1(n_1661), .A2(n_1645), .ZN(n_1428));
   NOR2_X1 i_894 (.A1(n_1662), .A2(n_1644), .ZN(n_1405));
   NOR2_X1 i_895 (.A1(n_1663), .A2(n_1643), .ZN(n_1382));
   NOR2_X1 i_896 (.A1(n_1658), .A2(n_1648), .ZN(n_1497));
   NOR2_X1 i_897 (.A1(n_1659), .A2(n_1647), .ZN(n_1474));
   NOR2_X1 i_898 (.A1(n_1660), .A2(n_1646), .ZN(n_1451));
   XNOR2_X1 i_899 (.A(n_971), .B(n_968), .ZN(Res_imm[24]));
   OAI22_X1 i_900 (.A1(n_773), .A2(n_938), .B1(n_1584), .B2(n_973), .ZN(n_968));
   AOI21_X1 i_901 (.A(n_1586), .B1(n_775), .B2(n_900), .ZN(n_971));
   AOI21_X1 i_902 (.A(n_1583), .B1(n_1569), .B2(n_975), .ZN(n_973));
   OAI21_X1 i_903 (.A(n_1536), .B1(n_1513), .B2(n_977), .ZN(n_975));
   NAND2_X1 i_904 (.A1(n_987), .A2(n_979), .ZN(n_977));
   AOI221_X1 i_909 (.A(n_981), .B1(n_989), .B2(n_983), .C1(n_376), .C2(n_378), 
      .ZN(n_979));
   NOR3_X1 i_910 (.A1(n_1621), .A2(n_990), .A3(n_1608), .ZN(n_981));
   INV_X1 i_911 (.A(n_985), .ZN(n_983));
   AOI22_X1 i_912 (.A1(n_268), .A2(n_270), .B1(n_304), .B2(n_271), .ZN(n_985));
   OAI211_X1 i_913 (.A(n_998), .B(n_989), .C1(n_268), .C2(n_270), .ZN(n_987));
   AOI211_X1 i_914 (.A(n_991), .B(n_990), .C1(n_1621), .C2(n_1608), .ZN(n_989));
   NOR2_X1 i_915 (.A1(n_376), .A2(n_378), .ZN(n_990));
   NOR2_X1 i_916 (.A1(n_304), .A2(n_271), .ZN(n_991));
   OAI221_X1 i_917 (.A(n_1008), .B1(n_1010), .B2(n_1007), .C1(n_1011), .C2(
      n_1005), .ZN(n_998));
   AOI22_X1 i_918 (.A1(n_236), .A2(n_238), .B1(n_206), .B2(n_208), .ZN(n_1005));
   AOI22_X1 i_919 (.A1(n_152), .A2(n_154), .B1(n_178), .B2(n_180), .ZN(n_1007));
   OAI211_X1 i_920 (.A(n_1009), .B(n_1164), .C1(n_152), .C2(n_154), .ZN(n_1008));
   INV_X1 i_921 (.A(n_1010), .ZN(n_1009));
   OAI222_X1 i_922 (.A1(n_178), .A2(n_180), .B1(n_206), .B2(n_208), .C1(n_236), 
      .C2(n_238), .ZN(n_1010));
   NOR2_X1 i_923 (.A1(n_236), .A2(n_238), .ZN(n_1011));
   OAI211_X1 i_924 (.A(n_1210), .B(n_1187), .C1(n_1256), .C2(n_1226), .ZN(n_1164));
   AOI21_X1 i_925 (.A(n_1233), .B1(n_128), .B2(n_130), .ZN(n_1187));
   OAI211_X1 i_926 (.A(n_106), .B(n_108), .C1(n_128), .C2(n_130), .ZN(n_1210));
   AOI22_X1 i_927 (.A1(n_68), .A2(n_70), .B1(n_86), .B2(n_88), .ZN(n_1226));
   AOI211_X1 i_932 (.A(n_1256), .B(n_1249), .C1(n_1490), .C2(n_1272), .ZN(n_1233));
   OAI22_X1 i_933 (.A1(n_68), .A2(n_70), .B1(n_52), .B2(n_54), .ZN(n_1249));
   OAI222_X1 i_934 (.A1(n_86), .A2(n_88), .B1(n_106), .B2(n_108), .C1(n_128), 
      .C2(n_130), .ZN(n_1256));
   OAI221_X1 i_935 (.A(n_1279), .B1(n_26), .B2(n_28), .C1(n_38), .C2(n_40), 
      .ZN(n_1272));
   OAI21_X1 i_936 (.A(n_1348), .B1(n_1325), .B2(n_1302), .ZN(n_1279));
   NOR2_X1 i_937 (.A1(n_16), .A2(n_18), .ZN(n_1302));
   AOI21_X1 i_938 (.A(n_1623), .B1(n_954), .B2(n_955), .ZN(n_1325));
   AOI22_X1 i_939 (.A1(n_16), .A2(n_18), .B1(n_26), .B2(n_28), .ZN(n_1348));
   AOI22_X1 i_940 (.A1(n_52), .A2(n_54), .B1(n_38), .B2(n_40), .ZN(n_1490));
   NOR2_X1 i_941 (.A1(n_1622), .A2(n_1619), .ZN(n_1513));
   NAND2_X1 i_942 (.A1(n_1622), .A2(n_1619), .ZN(n_1536));
   NAND2_X1 i_943 (.A1(n_460), .A2(n_419), .ZN(n_1569));
   NOR2_X1 i_944 (.A1(n_460), .A2(n_419), .ZN(n_1583));
   INV_X1 i_945 (.A(n_1585), .ZN(n_1584));
   NAND2_X1 i_946 (.A1(n_773), .A2(n_938), .ZN(n_1585));
   NOR2_X1 i_947 (.A1(n_775), .A2(n_900), .ZN(n_1586));
   INV_X1 i_948 (.A(n_305), .ZN(n_1608));
   INV_X1 i_949 (.A(n_379), .ZN(n_1619));
   INV_X1 i_950 (.A(n_340), .ZN(n_1621));
   INV_X1 i_955 (.A(n_418), .ZN(n_1622));
   INV_X1 i_956 (.A(n_763), .ZN(n_1623));
   INV_X1 i_957 (.A(A_imm[0]), .ZN(n_1625));
   INV_X1 i_958 (.A(A_imm[1]), .ZN(n_1628));
   INV_X1 i_959 (.A(A_imm[2]), .ZN(n_1629));
   INV_X1 i_960 (.A(A_imm[3]), .ZN(n_1630));
   INV_X1 i_961 (.A(A_imm[4]), .ZN(n_1631));
   INV_X1 i_962 (.A(A_imm[5]), .ZN(n_1632));
   INV_X1 i_963 (.A(A_imm[6]), .ZN(n_1633));
   INV_X1 i_964 (.A(A_imm[7]), .ZN(n_1634));
   INV_X1 i_965 (.A(A_imm[8]), .ZN(n_1639));
   INV_X1 i_966 (.A(A_imm[9]), .ZN(n_1640));
   INV_X1 i_967 (.A(A_imm[10]), .ZN(n_1641));
   INV_X1 i_968 (.A(A_imm[11]), .ZN(n_1642));
   INV_X1 i_969 (.A(A_imm[12]), .ZN(n_1643));
   INV_X1 i_970 (.A(A_imm[13]), .ZN(n_1644));
   INV_X1 i_971 (.A(A_imm[14]), .ZN(n_1645));
   INV_X1 i_972 (.A(A_imm[15]), .ZN(n_1646));
   INV_X1 i_973 (.A(A_imm[16]), .ZN(n_1647));
   INV_X1 i_978 (.A(A_imm[17]), .ZN(n_1648));
   INV_X1 i_979 (.A(A_imm[18]), .ZN(n_1649));
   INV_X1 i_980 (.A(A_imm[19]), .ZN(n_1650));
   INV_X1 i_981 (.A(A_imm[20]), .ZN(n_1651));
   INV_X1 i_982 (.A(A_imm[21]), .ZN(n_1652));
   INV_X1 i_983 (.A(A_imm[22]), .ZN(n_1653));
   INV_X1 i_984 (.A(A_imm[23]), .ZN(n_1654));
   INV_X1 i_985 (.A(B_imm[0]), .ZN(n_1655));
   INV_X1 i_986 (.A(B_imm[1]), .ZN(n_1656));
   INV_X1 i_987 (.A(B_imm[2]), .ZN(n_1657));
   INV_X1 i_988 (.A(B_imm[3]), .ZN(n_1658));
   INV_X1 i_989 (.A(B_imm[4]), .ZN(n_1659));
   INV_X1 i_990 (.A(B_imm[5]), .ZN(n_1660));
   INV_X1 i_991 (.A(B_imm[6]), .ZN(n_1661));
   INV_X1 i_992 (.A(B_imm[7]), .ZN(n_1662));
   INV_X1 i_993 (.A(B_imm[8]), .ZN(n_1663));
   INV_X1 i_994 (.A(B_imm[9]), .ZN(n_1664));
   INV_X1 i_995 (.A(B_imm[10]), .ZN(n_1665));
   INV_X1 i_996 (.A(B_imm[11]), .ZN(n_1666));
   INV_X1 i_999 (.A(B_imm[12]), .ZN(n_1667));
   INV_X1 i_1001 (.A(B_imm[13]), .ZN(n_1668));
   INV_X1 i_1002 (.A(B_imm[14]), .ZN(n_1669));
   INV_X1 i_1003 (.A(B_imm[15]), .ZN(n_1670));
   INV_X1 i_1004 (.A(B_imm[16]), .ZN(n_1672));
   INV_X1 i_1005 (.A(B_imm[17]), .ZN(n_1673));
   INV_X1 i_1006 (.A(B_imm[18]), .ZN(n_1674));
   INV_X1 i_1007 (.A(B_imm[19]), .ZN(n_1675));
   INV_X1 i_1008 (.A(B_imm[20]), .ZN(n_1676));
   INV_X1 i_1009 (.A(B_imm[21]), .ZN(n_1677));
   INV_X1 i_1010 (.A(B_imm[22]), .ZN(n_1678));
   FA_X1 i_1011 (.A(n_1157), .B(n_1180), .CI(n_1203), .CO(n_945), .S(n_944));
   FA_X1 i_1012 (.A(n_1156), .B(n_1179), .CI(n_945), .CO(n_961), .S(n_960));
   FA_X1 i_1013 (.A(n_1087), .B(n_1110), .CI(n_1133), .CO(n_959), .S(n_958));
   FA_X1 i_1014 (.A(n_1018), .B(n_1041), .CI(n_1064), .CO(n_957), .S(n_956));
   FA_X1 i_1015 (.A(n_960), .B(n_958), .CI(n_956), .CO(n_965), .S(n_964));
   FA_X1 i_1016 (.A(n_1088), .B(n_1111), .CI(n_1134), .CO(n_943), .S(n_942));
   FA_X1 i_1017 (.A(n_1019), .B(n_1042), .CI(n_1065), .CO(n_941), .S(n_940));
   FA_X1 i_1018 (.A(n_1158), .B(n_1181), .CI(n_1204), .CO(n_927), .S(n_926));
   FA_X1 i_1019 (.A(n_1089), .B(n_1112), .CI(n_1135), .CO(n_925), .S(n_924));
   FA_X1 i_1022 (.A(n_1020), .B(n_1043), .CI(n_1066), .CO(n_923), .S(n_922));
   FA_X1 i_1024 (.A(n_927), .B(n_925), .CI(n_923), .CO(n_947), .S(n_946));
   FA_X1 i_1025 (.A(n_943), .B(n_941), .CI(n_947), .CO(n_963), .S(n_962));
   FA_X1 i_1026 (.A(n_1159), .B(n_1182), .CI(n_1205), .CO(n_907), .S(n_906));
   FA_X1 i_1027 (.A(n_1090), .B(n_1113), .CI(n_1136), .CO(n_905), .S(n_904));
   FA_X1 i_1028 (.A(n_1227), .B(n_907), .CI(n_905), .CO(n_929), .S(n_928));
   FA_X1 i_1029 (.A(n_929), .B(n_944), .CI(n_942), .CO(n_949), .S(n_948));
   FA_X1 i_1030 (.A(n_1021), .B(n_1044), .CI(n_1067), .CO(n_903), .S(n_902));
   FA_X1 i_1031 (.A(n_1160), .B(n_1183), .CI(n_1206), .CO(n_885), .S(n_884));
   FA_X1 i_1032 (.A(n_1091), .B(n_1114), .CI(n_1137), .CO(n_883), .S(n_882));
   FA_X1 i_1033 (.A(n_1022), .B(n_1045), .CI(n_1068), .CO(n_881), .S(n_880));
   FA_X1 i_1034 (.A(n_885), .B(n_883), .CI(n_881), .CO(n_911), .S(n_910));
   FA_X1 i_1035 (.A(n_1229), .B(n_1252), .CI(n_1275), .CO(n_887), .S(n_886));
   FA_X1 i_1036 (.A(n_1228), .B(n_1251), .CI(n_887), .CO(n_909), .S(n_908));
   FA_X1 i_1037 (.A(n_903), .B(n_911), .CI(n_909), .CO(n_931), .S(n_930));
   FA_X1 i_1038 (.A(n_940), .B(n_931), .CI(n_946), .CO(n_951), .S(n_950));
   FA_X1 i_1039 (.A(n_962), .B(n_949), .CI(n_951), .CO(n_967), .S(n_966));
   FA_X1 i_1040 (.A(n_926), .B(n_924), .CI(n_922), .CO(n_933), .S(n_932));
   FA_X1 i_1041 (.A(n_933), .B(n_948), .CI(n_950), .CO(n_953), .S(n_952));
   FA_X1 i_1042 (.A(n_964), .B(n_966), .CI(n_953), .CO(n_969), .S(n_1679));
   FA_X1 i_1044 (.A(n_1086), .B(n_1109), .CI(n_1132), .CO(n_1680), .S(n_972));
   FA_X1 i_1045 (.A(n_1017), .B(n_1040), .CI(n_1063), .CO(n_1681), .S(n_970));
   FA_X1 i_1047 (.A(n_961), .B(n_972), .CI(n_970), .CO(n_1682), .S(n_976));
   FA_X1 i_1048 (.A(n_1155), .B(n_959), .CI(n_957), .CO(n_1683), .S(n_974));
   FA_X1 i_1049 (.A(n_963), .B(n_974), .CI(n_965), .CO(n_1684), .S(n_978));
   FA_X1 i_1050 (.A(n_976), .B(n_967), .CI(n_978), .CO(n_1685), .S(n_980));
   FA_X1 i_1051 (.A(n_1230), .B(n_1253), .CI(n_1276), .CO(n_863), .S(n_862));
   FA_X1 i_1052 (.A(n_1161), .B(n_1184), .CI(n_1207), .CO(n_861), .S(n_860));
   FA_X1 i_1053 (.A(n_1092), .B(n_1115), .CI(n_1138), .CO(n_859), .S(n_858));
   FA_X1 i_1054 (.A(n_863), .B(n_861), .CI(n_859), .CO(n_889), .S(n_888));
   FA_X1 i_1055 (.A(n_889), .B(n_908), .CI(n_906), .CO(n_913), .S(n_912));
   FA_X1 i_1056 (.A(n_928), .B(n_913), .CI(n_930), .CO(n_935), .S(n_934));
   FA_X1 i_1057 (.A(n_904), .B(n_902), .CI(n_910), .CO(n_915), .S(n_914));
   FA_X1 i_1058 (.A(n_884), .B(n_882), .CI(n_880), .CO(n_893), .S(n_892));
   FA_X1 i_1059 (.A(n_1023), .B(n_1046), .CI(n_1069), .CO(n_857), .S(n_856));
   FA_X1 i_1060 (.A(n_1231), .B(n_1254), .CI(n_1277), .CO(n_837), .S(n_836));
   FA_X1 i_1061 (.A(n_1162), .B(n_1185), .CI(n_1208), .CO(n_835), .S(n_834));
   FA_X1 i_1062 (.A(n_1299), .B(n_837), .CI(n_835), .CO(n_865), .S(n_864));
   FA_X1 i_1063 (.A(n_857), .B(n_865), .CI(n_886), .CO(n_891), .S(n_890));
   FA_X1 i_1065 (.A(n_1093), .B(n_1116), .CI(n_1139), .CO(n_833), .S(n_832));
   FA_X1 i_1068 (.A(n_1024), .B(n_1047), .CI(n_1070), .CO(n_831), .S(n_830));
   FA_X1 i_1069 (.A(n_1232), .B(n_1255), .CI(n_1278), .CO(n_809), .S(n_808));
   FA_X1 i_1070 (.A(n_1163), .B(n_1186), .CI(n_1209), .CO(n_807), .S(n_806));
   FA_X1 i_1071 (.A(n_1094), .B(n_1117), .CI(n_1140), .CO(n_805), .S(n_804));
   FA_X1 i_1072 (.A(n_809), .B(n_807), .CI(n_805), .CO(n_841), .S(n_840));
   FA_X1 i_1073 (.A(n_833), .B(n_831), .CI(n_841), .CO(n_867), .S(n_866));
   FA_X1 i_1074 (.A(n_1301), .B(n_1324), .CI(n_1347), .CO(n_811), .S(n_810));
   FA_X1 i_1075 (.A(n_1300), .B(n_1323), .CI(n_811), .CO(n_839), .S(n_838));
   FA_X1 i_1076 (.A(n_839), .B(n_862), .CI(n_860), .CO(n_869), .S(n_868));
   FA_X1 i_1077 (.A(n_867), .B(n_888), .CI(n_869), .CO(n_895), .S(n_894));
   FA_X1 i_1078 (.A(n_893), .B(n_891), .CI(n_895), .CO(n_917), .S(n_916));
   FA_X1 i_1079 (.A(n_915), .B(n_932), .CI(n_917), .CO(n_937), .S(n_936));
   FA_X1 i_1080 (.A(n_935), .B(n_937), .CI(n_952), .CO(n_1687), .S(n_1686));
   FA_X1 i_1081 (.A(n_836), .B(n_834), .CI(n_832), .CO(n_845), .S(n_844));
   FA_X1 i_1082 (.A(n_1025), .B(n_1048), .CI(n_1071), .CO(n_803), .S(n_802));
   FA_X1 i_1083 (.A(n_731), .B(n_734), .CI(n_736), .CO(n_781), .S(n_1688));
   FA_X1 i_1084 (.A(n_702), .B(n_704), .CI(n_729), .CO(n_779), .S(n_1690));
   FA_X1 i_1085 (.A(n_667), .B(n_668), .CI(n_669), .CO(n_777), .S(n_1691));
   FA_X1 i_1086 (.A(n_781), .B(n_779), .CI(n_777), .CO(n_813), .S(n_812));
   FA_X1 i_1087 (.A(n_803), .B(n_813), .CI(n_838), .CO(n_843), .S(n_842));
   FA_X1 i_1088 (.A(n_864), .B(n_845), .CI(n_843), .CO(n_873), .S(n_872));
   FA_X1 i_1089 (.A(n_858), .B(n_856), .CI(n_866), .CO(n_871), .S(n_870));
   FA_X1 i_1090 (.A(n_890), .B(n_873), .CI(n_871), .CO(n_897), .S(n_896));
   FA_X1 i_1091 (.A(n_914), .B(n_912), .CI(n_897), .CO(n_919), .S(n_918));
   FA_X1 i_1092 (.A(n_934), .B(n_919), .CI(n_936), .CO(n_1693), .S(n_1692));
   FA_X1 i_1093 (.A(n_539), .B(n_537), .CI(n_543), .CO(n_815), .S(n_814));
   FA_X1 i_1094 (.A(n_830), .B(n_815), .CI(n_840), .CO(n_847), .S(n_846));
   FA_X1 i_1095 (.A(n_847), .B(n_870), .CI(n_868), .CO(n_875), .S(n_874));
   FA_X1 i_1096 (.A(n_892), .B(n_894), .CI(n_875), .CO(n_899), .S(n_898));
   FA_X1 i_1097 (.A(n_916), .B(n_899), .CI(n_918), .CO(n_1694), .S(n_920));
   FA_X1 i_1098 (.A(n_806), .B(n_804), .CI(n_802), .CO(n_819), .S(n_818));
   FA_X1 i_1099 (.A(n_541), .B(n_810), .CI(n_808), .CO(n_817), .S(n_816));
   FA_X1 i_1100 (.A(n_819), .B(n_817), .CI(n_842), .CO(n_849), .S(n_848));
   FA_X1 i_1101 (.A(n_814), .B(n_812), .CI(n_549), .CO(n_821), .S(n_820));
   FA_X1 i_1102 (.A(n_821), .B(n_844), .CI(n_846), .CO(n_851), .S(n_850));
   FA_X1 i_1103 (.A(n_849), .B(n_872), .CI(n_851), .CO(n_877), .S(n_876));
   FA_X1 i_1104 (.A(n_896), .B(n_877), .CI(n_898), .CO(n_901), .S(n_1695));
   FA_X1 i_1105 (.A(n_547), .B(n_666), .CI(n_631), .CO(n_823), .S(n_822));
   FA_X1 i_1106 (.A(n_818), .B(n_816), .CI(n_795), .CO(n_825), .S(n_824));
   FA_X1 i_1107 (.A(n_823), .B(n_848), .CI(n_825), .CO(n_853), .S(n_852));
   FA_X1 i_1108 (.A(n_853), .B(n_874), .CI(n_876), .CO(n_1697), .S(n_1696));
   FA_X1 i_1109 (.A(n_820), .B(n_822), .CI(n_797), .CO(n_827), .S(n_826));
   FA_X1 i_1110 (.A(n_850), .B(n_827), .CI(n_852), .CO(n_1699), .S(n_1698));
   FA_X1 i_1111 (.A(n_545), .B(n_527), .CI(n_531), .CO(n_795), .S(n_794));
   FA_X1 i_1112 (.A(n_511), .B(n_523), .CI(n_521), .CO(n_765), .S(n_1700));
   FA_X1 i_1113 (.A(n_513), .B(n_529), .CI(n_525), .CO(n_767), .S(n_766));
   FA_X1 i_1114 (.A(n_765), .B(n_794), .CI(n_767), .CO(n_799), .S(n_798));
   FA_X1 i_1115 (.A(n_548), .B(n_629), .CI(n_664), .CO(n_797), .S(n_796));
   FA_X1 i_1116 (.A(n_824), .B(n_799), .CI(n_826), .CO(n_1703), .S(n_1701));
   FA_X1 i_1117 (.A(n_796), .B(n_535), .CI(n_798), .CO(n_1705), .S(n_1704));
   FA_X1 i_1118 (.A(n_766), .B(n_519), .CI(n_533), .CO(n_1707), .S(n_1706));
   FA_X1 i_1119 (.A(n_505), .B(n_504), .CI(n_507), .CO(n_1709), .S(n_1708));
   FA_X1 i_1120 (.A(n_515), .B(n_509), .CI(n_517), .CO(n_1711), .S(n_1710));
   FA_X1 i_1121 (.A(n_169), .B(n_167), .CI(n_461), .CO(n_1713), .S(n_1712));
   NOR2_X1 i_1122 (.A1(n_1677), .A2(n_1642), .ZN(n_1071));
   NOR2_X1 i_1123 (.A1(n_1678), .A2(n_1641), .ZN(n_1048));
   NOR2_X1 i_1124 (.A1(n_1654), .A2(n_1640), .ZN(n_1025));
   NOR2_X1 i_1125 (.A1(n_1654), .A2(n_1664), .ZN(n_1347));
   NOR2_X1 i_1126 (.A1(n_1653), .A2(n_1665), .ZN(n_1324));
   NOR2_X1 i_1127 (.A1(n_1652), .A2(n_1666), .ZN(n_1301));
   NOR2_X1 i_1128 (.A1(n_1654), .A2(n_1665), .ZN(n_1323));
   NOR2_X1 i_1129 (.A1(n_1653), .A2(n_1666), .ZN(n_1300));
   NOR2_X1 i_1130 (.A1(n_1674), .A2(n_1645), .ZN(n_1140));
   NOR2_X1 i_1131 (.A1(n_1675), .A2(n_1644), .ZN(n_1117));
   NOR2_X1 i_1132 (.A1(n_1676), .A2(n_1643), .ZN(n_1094));
   NOR2_X1 i_1133 (.A1(n_1670), .A2(n_1648), .ZN(n_1209));
   NOR2_X1 i_1134 (.A1(n_1672), .A2(n_1647), .ZN(n_1186));
   NOR2_X1 i_1135 (.A1(n_1673), .A2(n_1646), .ZN(n_1163));
   NOR2_X1 i_1136 (.A1(n_1651), .A2(n_1667), .ZN(n_1278));
   NOR2_X1 i_1137 (.A1(n_1650), .A2(n_1668), .ZN(n_1255));
   NOR2_X1 i_1138 (.A1(n_1649), .A2(n_1669), .ZN(n_1232));
   NOR2_X1 i_1139 (.A1(n_1677), .A2(n_1643), .ZN(n_1070));
   NOR2_X1 i_1140 (.A1(n_1678), .A2(n_1642), .ZN(n_1047));
   NOR2_X1 i_1141 (.A1(n_1654), .A2(n_1641), .ZN(n_1024));
   NOR2_X1 i_1142 (.A1(n_1674), .A2(n_1646), .ZN(n_1139));
   NOR2_X1 i_1143 (.A1(n_1675), .A2(n_1645), .ZN(n_1116));
   NOR2_X1 i_1144 (.A1(n_1676), .A2(n_1644), .ZN(n_1093));
   NOR2_X1 i_1145 (.A1(n_1670), .A2(n_1649), .ZN(n_1208));
   NOR2_X1 i_1146 (.A1(n_1672), .A2(n_1648), .ZN(n_1185));
   NOR2_X1 i_1147 (.A1(n_1673), .A2(n_1647), .ZN(n_1162));
   NOR2_X1 i_1148 (.A1(n_1652), .A2(n_1667), .ZN(n_1277));
   NOR2_X1 i_1149 (.A1(n_1651), .A2(n_1668), .ZN(n_1254));
   NOR2_X1 i_1150 (.A1(n_1650), .A2(n_1669), .ZN(n_1231));
   NOR2_X1 i_1151 (.A1(n_1654), .A2(n_1666), .ZN(n_1299));
   NOR2_X1 i_1152 (.A1(n_1677), .A2(n_1644), .ZN(n_1069));
   NOR2_X1 i_1153 (.A1(n_1678), .A2(n_1643), .ZN(n_1046));
   NOR2_X1 i_1154 (.A1(n_1654), .A2(n_1642), .ZN(n_1023));
   NOR2_X1 i_1155 (.A1(n_1674), .A2(n_1647), .ZN(n_1138));
   NOR2_X1 i_1156 (.A1(n_1675), .A2(n_1646), .ZN(n_1115));
   NOR2_X1 i_1157 (.A1(n_1676), .A2(n_1645), .ZN(n_1092));
   NOR2_X1 i_1158 (.A1(n_1670), .A2(n_1650), .ZN(n_1207));
   NOR2_X1 i_1159 (.A1(n_1672), .A2(n_1649), .ZN(n_1184));
   NOR2_X1 i_1160 (.A1(n_1673), .A2(n_1648), .ZN(n_1161));
   NOR2_X1 i_1161 (.A1(n_1653), .A2(n_1667), .ZN(n_1276));
   NOR2_X1 i_1162 (.A1(n_1652), .A2(n_1668), .ZN(n_1253));
   NOR2_X1 i_1163 (.A1(n_1651), .A2(n_1669), .ZN(n_1230));
   NOR2_X1 i_1164 (.A1(n_1673), .A2(n_1654), .ZN(n_1155));
   NOR2_X1 i_1165 (.A1(n_1650), .A2(n_1677), .ZN(n_1063));
   NOR2_X1 i_1166 (.A1(n_1678), .A2(n_1649), .ZN(n_1040));
   NOR2_X1 i_1167 (.A1(n_1654), .A2(n_1648), .ZN(n_1017));
   NOR2_X1 i_1168 (.A1(n_1653), .A2(n_1674), .ZN(n_1132));
   NOR2_X1 i_1169 (.A1(n_1652), .A2(n_1675), .ZN(n_1109));
   NOR2_X1 i_1170 (.A1(n_1676), .A2(n_1651), .ZN(n_1086));
   NOR2_X1 i_1171 (.A1(n_1654), .A2(n_1667), .ZN(n_1275));
   NOR2_X1 i_1172 (.A1(n_1653), .A2(n_1668), .ZN(n_1252));
   NOR2_X1 i_1173 (.A1(n_1652), .A2(n_1669), .ZN(n_1229));
   NOR2_X1 i_1174 (.A1(n_1654), .A2(n_1668), .ZN(n_1251));
   NOR2_X1 i_1175 (.A1(n_1653), .A2(n_1669), .ZN(n_1228));
   NOR2_X1 i_1176 (.A1(n_1677), .A2(n_1645), .ZN(n_1068));
   NOR2_X1 i_1177 (.A1(n_1678), .A2(n_1644), .ZN(n_1045));
   NOR2_X1 i_1178 (.A1(n_1654), .A2(n_1643), .ZN(n_1022));
   NOR2_X1 i_1179 (.A1(n_1674), .A2(n_1648), .ZN(n_1137));
   NOR2_X1 i_1180 (.A1(n_1675), .A2(n_1647), .ZN(n_1114));
   NOR2_X1 i_1181 (.A1(n_1676), .A2(n_1646), .ZN(n_1091));
   NOR2_X1 i_1182 (.A1(n_1670), .A2(n_1651), .ZN(n_1206));
   NOR2_X1 i_1183 (.A1(n_1672), .A2(n_1650), .ZN(n_1183));
   NOR2_X1 i_1184 (.A1(n_1673), .A2(n_1649), .ZN(n_1160));
   NOR2_X1 i_1185 (.A1(n_1677), .A2(n_1646), .ZN(n_1067));
   NOR2_X1 i_1186 (.A1(n_1678), .A2(n_1645), .ZN(n_1044));
   NOR2_X1 i_1187 (.A1(n_1654), .A2(n_1644), .ZN(n_1021));
   NOR2_X1 i_1188 (.A1(n_1674), .A2(n_1649), .ZN(n_1136));
   NOR2_X1 i_1189 (.A1(n_1675), .A2(n_1648), .ZN(n_1113));
   NOR2_X1 i_1190 (.A1(n_1676), .A2(n_1647), .ZN(n_1090));
   NOR2_X1 i_1191 (.A1(n_1652), .A2(n_1670), .ZN(n_1205));
   NOR2_X1 i_1192 (.A1(n_1672), .A2(n_1651), .ZN(n_1182));
   NOR2_X1 i_1193 (.A1(n_1673), .A2(n_1650), .ZN(n_1159));
   NOR2_X1 i_1194 (.A1(n_1654), .A2(n_1669), .ZN(n_1227));
   NOR2_X1 i_1195 (.A1(n_1647), .A2(n_1677), .ZN(n_1066));
   NOR2_X1 i_1196 (.A1(n_1678), .A2(n_1646), .ZN(n_1043));
   NOR2_X1 i_1197 (.A1(n_1654), .A2(n_1645), .ZN(n_1020));
   NOR2_X1 i_1198 (.A1(n_1650), .A2(n_1674), .ZN(n_1135));
   NOR2_X1 i_1199 (.A1(n_1675), .A2(n_1649), .ZN(n_1112));
   NOR2_X1 i_1200 (.A1(n_1676), .A2(n_1648), .ZN(n_1089));
   NOR2_X1 i_1201 (.A1(n_1653), .A2(n_1670), .ZN(n_1204));
   NOR2_X1 i_1202 (.A1(n_1672), .A2(n_1652), .ZN(n_1181));
   NOR2_X1 i_1203 (.A1(n_1673), .A2(n_1651), .ZN(n_1158));
   NOR2_X1 i_1204 (.A1(n_1648), .A2(n_1677), .ZN(n_1065));
   NOR2_X1 i_1205 (.A1(n_1647), .A2(n_1678), .ZN(n_1042));
   NOR2_X1 i_1206 (.A1(n_1654), .A2(n_1646), .ZN(n_1019));
   NOR2_X1 i_1207 (.A1(n_1651), .A2(n_1674), .ZN(n_1134));
   NOR2_X1 i_1208 (.A1(n_1650), .A2(n_1675), .ZN(n_1111));
   NOR2_X1 i_1209 (.A1(n_1676), .A2(n_1649), .ZN(n_1088));
   NOR2_X1 i_1210 (.A1(n_1677), .A2(n_1649), .ZN(n_1064));
   NOR2_X1 i_1211 (.A1(n_1678), .A2(n_1648), .ZN(n_1041));
   NOR2_X1 i_1212 (.A1(n_1654), .A2(n_1647), .ZN(n_1018));
   NOR2_X1 i_1213 (.A1(n_1652), .A2(n_1674), .ZN(n_1133));
   NOR2_X1 i_1214 (.A1(n_1675), .A2(n_1651), .ZN(n_1110));
   NOR2_X1 i_1215 (.A1(n_1676), .A2(n_1650), .ZN(n_1087));
   NOR2_X1 i_1216 (.A1(n_1654), .A2(n_1670), .ZN(n_1203));
   NOR2_X1 i_1217 (.A1(n_1653), .A2(n_1672), .ZN(n_1180));
   NOR2_X1 i_1218 (.A1(n_1673), .A2(n_1652), .ZN(n_1157));
   NOR2_X1 i_1219 (.A1(n_1672), .A2(n_1654), .ZN(n_1179));
   NOR2_X1 i_1220 (.A1(n_1673), .A2(n_1653), .ZN(n_1156));
   XOR2_X1 i_1221 (.A(n_1715), .B(n_1714), .Z(Res_imm[40]));
   OAI22_X1 i_1222 (.A1(n_1679), .A2(n_1687), .B1(n_1770), .B2(n_1716), .ZN(
      n_1714));
   OR2_X1 i_1223 (.A1(n_1774), .A2(n_1772), .ZN(n_1715));
   AOI21_X1 i_1224 (.A(n_1769), .B1(n_1768), .B2(n_1717), .ZN(n_1716));
   INV_X1 i_1225 (.A(n_1718), .ZN(n_1717));
   AOI21_X1 i_1226 (.A(n_1766), .B1(n_1720), .B2(n_1719), .ZN(n_1718));
   NAND2_X1 i_1227 (.A1(n_1692), .A2(n_1694), .ZN(n_1719));
   AOI21_X1 i_1228 (.A(n_1725), .B1(n_1730), .B2(n_1727), .ZN(n_1720));
   OAI221_X1 i_1229 (.A(n_1764), .B1(n_1761), .B2(n_1760), .C1(n_1728), .C2(
      n_1726), .ZN(n_1725));
   AND2_X1 i_1230 (.A1(n_1755), .A2(n_1754), .ZN(n_1726));
   NOR2_X1 i_1231 (.A1(n_1753), .A2(n_1728), .ZN(n_1727));
   OR3_X1 i_1232 (.A1(n_1761), .A2(n_1758), .A3(n_1759), .ZN(n_1728));
   INV_X1 i_1233 (.A(n_1730), .ZN(n_1729));
   OAI221_X1 i_1234 (.A(n_1731), .B1(n_1778), .B2(n_1777), .C1(n_1752), .C2(
      n_1737), .ZN(n_1730));
   OR3_X1 i_1235 (.A1(n_770), .A2(n_1737), .A3(n_1732), .ZN(n_1731));
   NOR3_X1 i_1236 (.A1(n_1775), .A2(n_1744), .A3(n_1733), .ZN(n_1732));
   AOI21_X1 i_1237 (.A(n_1736), .B1(n_1745), .B2(n_1734), .ZN(n_1733));
   OAI21_X1 i_1238 (.A(n_1743), .B1(n_1739), .B2(n_1735), .ZN(n_1734));
   AOI21_X1 i_1239 (.A(n_1738), .B1(n_979), .B2(n_987), .ZN(n_1735));
   NOR2_X1 i_1240 (.A1(n_1709), .A2(n_1710), .ZN(n_1736));
   NOR2_X1 i_1241 (.A1(n_1701), .A2(n_1705), .ZN(n_1737));
   NAND2_X1 i_1242 (.A1(n_1536), .A2(n_771), .ZN(n_1738));
   INV_X1 i_1243 (.A(n_1740), .ZN(n_1739));
   AOI21_X1 i_1244 (.A(n_1741), .B1(n_775), .B2(n_900), .ZN(n_1740));
   OAI21_X1 i_1245 (.A(n_762), .B1(n_1586), .B2(n_1585), .ZN(n_1741));
   INV_X1 i_1246 (.A(n_1743), .ZN(n_1742));
   NOR2_X1 i_1247 (.A1(n_768), .A2(n_764), .ZN(n_1743));
   AND2_X1 i_1248 (.A1(n_1706), .A2(n_1711), .ZN(n_1744));
   AOI221_X1 i_1249 (.A(n_1746), .B1(n_1708), .B2(n_1713), .C1(n_1776), .C2(
      n_1751), .ZN(n_1745));
   AOI21_X1 i_1250 (.A(n_768), .B1(n_760), .B2(n_758), .ZN(n_1746));
   AND2_X1 i_1251 (.A1(n_1712), .A2(n_168), .ZN(n_1751));
   NAND2_X1 i_1252 (.A1(n_1704), .A2(n_1707), .ZN(n_1752));
   NOR2_X1 i_1253 (.A1(n_1698), .A2(n_1703), .ZN(n_1753));
   NAND2_X1 i_1254 (.A1(n_1696), .A2(n_1699), .ZN(n_1754));
   NAND2_X1 i_1255 (.A1(n_1698), .A2(n_1703), .ZN(n_1755));
   NOR2_X1 i_1256 (.A1(n_1696), .A2(n_1699), .ZN(n_1758));
   NOR2_X1 i_1257 (.A1(n_1695), .A2(n_1697), .ZN(n_1759));
   NAND2_X1 i_1258 (.A1(n_1695), .A2(n_1697), .ZN(n_1760));
   NOR2_X1 i_1259 (.A1(n_920), .A2(n_901), .ZN(n_1761));
   INV_X1 i_1260 (.A(n_1764), .ZN(n_1762));
   NAND2_X1 i_1261 (.A1(n_920), .A2(n_901), .ZN(n_1764));
   NOR2_X1 i_1262 (.A1(n_1692), .A2(n_1694), .ZN(n_1766));
   NAND2_X1 i_1263 (.A1(n_1686), .A2(n_1693), .ZN(n_1768));
   NOR2_X1 i_1264 (.A1(n_1686), .A2(n_1693), .ZN(n_1769));
   INV_X1 i_1265 (.A(n_1771), .ZN(n_1770));
   NAND2_X1 i_1266 (.A1(n_1679), .A2(n_1687), .ZN(n_1771));
   AND2_X1 i_1267 (.A1(n_969), .A2(n_980), .ZN(n_1772));
   NOR2_X1 i_1268 (.A1(n_969), .A2(n_980), .ZN(n_1774));
   INV_X1 i_1269 (.A(n_761), .ZN(n_1775));
   INV_X1 i_1270 (.A(n_769), .ZN(n_1776));
   INV_X1 i_1271 (.A(n_1705), .ZN(n_1777));
   INV_X1 i_1272 (.A(n_1701), .ZN(n_1778));
   FA_X1 i_1273 (.A(n_1085), .B(n_1108), .CI(n_1131), .CO(n_1779), .S(n_984));
   FA_X1 i_1274 (.A(n_1016), .B(n_1039), .CI(n_1062), .CO(n_1780), .S(n_982));
   FA_X1 i_1275 (.A(n_1680), .B(n_1681), .CI(n_1683), .CO(n_1781), .S(n_986));
   FA_X1 i_1276 (.A(n_984), .B(n_982), .CI(n_986), .CO(n_1782), .S(n_988));
   FA_X1 i_1277 (.A(n_1682), .B(n_1684), .CI(n_988), .CO(n_1784), .S(n_1783));
   NOR2_X1 i_1278 (.A1(n_1677), .A2(n_1651), .ZN(n_1062));
   NOR2_X1 i_1279 (.A1(n_1678), .A2(n_1650), .ZN(n_1039));
   NOR2_X1 i_1280 (.A1(n_1654), .A2(n_1649), .ZN(n_1016));
   NOR2_X1 i_1281 (.A1(n_1674), .A2(n_1654), .ZN(n_1131));
   NOR2_X1 i_1282 (.A1(n_1675), .A2(n_1653), .ZN(n_1108));
   NOR2_X1 i_1283 (.A1(n_1676), .A2(n_1652), .ZN(n_1085));
   XOR2_X1 i_1284 (.A(n_1787), .B(n_1785), .Z(Res_imm[41]));
   OAI21_X1 i_1285 (.A(n_1786), .B1(n_1783), .B2(n_1685), .ZN(n_1785));
   NAND2_X1 i_1286 (.A1(n_1783), .A2(n_1685), .ZN(n_1786));
   AOI211_X1 i_1287 (.A(n_1772), .B(n_1790), .C1(n_1789), .C2(n_1788), .ZN(
      n_1787));
   OAI211_X1 i_1288 (.A(n_1719), .B(n_1768), .C1(n_1766), .C2(n_1720), .ZN(
      n_1788));
   NOR3_X1 i_1289 (.A1(n_1774), .A2(n_1791), .A3(n_1769), .ZN(n_1789));
   NOR2_X1 i_1290 (.A1(n_1774), .A2(n_1771), .ZN(n_1790));
   NOR2_X1 i_1291 (.A1(n_1687), .A2(n_1679), .ZN(n_1791));
   FA_X1 i_1292 (.A(n_1014), .B(n_1037), .CI(n_1060), .CO(n_1001), .S(n_1000));
   FA_X1 i_1293 (.A(n_1015), .B(n_1038), .CI(n_1061), .CO(n_993), .S(n_992));
   FA_X1 i_1294 (.A(n_1084), .B(n_1107), .CI(n_1779), .CO(n_995), .S(n_994));
   FA_X1 i_1295 (.A(n_1083), .B(n_993), .CI(n_995), .CO(n_1003), .S(n_1002));
   FA_X1 i_1296 (.A(n_1780), .B(n_994), .CI(n_992), .CO(n_997), .S(n_996));
   FA_X1 i_1297 (.A(n_1000), .B(n_1002), .CI(n_997), .CO(n_1792), .S(n_1004));
   FA_X1 i_1298 (.A(n_1013), .B(n_1036), .CI(n_1059), .CO(n_1793), .S(n_1006));
   FA_X1 i_1299 (.A(n_1001), .B(n_1006), .CI(n_1003), .CO(n_1795), .S(n_1794));
   FA_X1 i_1300 (.A(n_1781), .B(n_1782), .CI(n_996), .CO(n_999), .S(n_1796));
   NOR2_X1 i_1301 (.A1(n_1677), .A2(n_1654), .ZN(n_1059));
   NOR2_X1 i_1302 (.A1(n_1653), .A2(n_1678), .ZN(n_1036));
   NOR2_X1 i_1303 (.A1(n_1652), .A2(n_1654), .ZN(n_1013));
   NOR2_X1 i_1304 (.A1(n_1675), .A2(n_1654), .ZN(n_1107));
   NOR2_X1 i_1305 (.A1(n_1676), .A2(n_1653), .ZN(n_1084));
   NOR2_X1 i_1306 (.A1(n_1677), .A2(n_1652), .ZN(n_1061));
   NOR2_X1 i_1307 (.A1(n_1678), .A2(n_1651), .ZN(n_1038));
   NOR2_X1 i_1308 (.A1(n_1650), .A2(n_1654), .ZN(n_1015));
   NOR2_X1 i_1309 (.A1(n_1676), .A2(n_1654), .ZN(n_1083));
   NOR2_X1 i_1310 (.A1(n_1677), .A2(n_1653), .ZN(n_1060));
   NOR2_X1 i_1311 (.A1(n_1678), .A2(n_1652), .ZN(n_1037));
   NOR2_X1 i_1312 (.A1(n_1654), .A2(n_1651), .ZN(n_1014));
   NOR2_X1 i_1313 (.A1(n_1792), .A2(n_1794), .ZN(n_1797));
   AND2_X1 i_1314 (.A1(n_1792), .A2(n_1794), .ZN(n_1798));
   NAND2_X1 i_1315 (.A1(n_1004), .A2(n_999), .ZN(n_1799));
   NOR2_X1 i_1316 (.A1(n_1004), .A2(n_999), .ZN(n_1800));
   NOR2_X1 i_1317 (.A1(n_1796), .A2(n_1784), .ZN(n_1801));
   NOR2_X1 i_1318 (.A1(n_1801), .A2(n_1800), .ZN(n_1802));
   NOR2_X1 i_1319 (.A1(n_1685), .A2(n_1783), .ZN(n_1803));
   AOI21_X1 i_1320 (.A(n_1803), .B1(n_1787), .B2(n_1786), .ZN(n_1804));
   NAND2_X1 i_1321 (.A1(n_1796), .A2(n_1784), .ZN(n_1805));
   INV_X1 i_1322 (.A(n_1805), .ZN(n_1806));
   OAI21_X1 i_1323 (.A(n_1802), .B1(n_1804), .B2(n_1806), .ZN(n_1807));
   NAND2_X1 i_1324 (.A1(n_1807), .A2(n_1799), .ZN(n_1808));
   NOR2_X1 i_1325 (.A1(n_1798), .A2(n_1797), .ZN(n_1809));
   XOR2_X1 i_1326 (.A(n_1808), .B(n_1809), .Z(Res_imm[44]));
   NOR2_X1 i_1327 (.A1(n_1806), .A2(n_1801), .ZN(n_1810));
   INV_X1 i_1328 (.A(n_1799), .ZN(n_1811));
   FA_X1 i_1329 (.A(n_1012), .B(n_1035), .CI(n_1793), .CO(n_1813), .S(n_1812));
   NOR2_X1 i_1330 (.A1(n_1654), .A2(n_1678), .ZN(n_1035));
   NOR2_X1 i_1331 (.A1(n_1654), .A2(n_1653), .ZN(n_1012));
   XNOR2_X1 i_1332 (.A(n_1815), .B(n_1814), .ZN(Res_imm[45]));
   AOI22_X1 i_1333 (.A1(n_1812), .A2(n_1819), .B1(n_1821), .B2(n_1795), .ZN(
      n_1814));
   OAI221_X1 i_1334 (.A(n_1820), .B1(n_1797), .B2(n_1799), .C1(n_1818), .C2(
      n_1816), .ZN(n_1815));
   INV_X1 i_1335 (.A(n_1817), .ZN(n_1816));
   OAI211_X1 i_1336 (.A(n_1786), .B(n_1805), .C1(n_1803), .C2(n_1787), .ZN(
      n_1817));
   OAI21_X1 i_1337 (.A(n_1802), .B1(n_1792), .B2(n_1794), .ZN(n_1818));
   INV_X1 i_1338 (.A(n_1795), .ZN(n_1819));
   INV_X1 i_1339 (.A(n_1798), .ZN(n_1820));
   INV_X1 i_1340 (.A(n_1812), .ZN(n_1821));
endmodule

module VM(Res, OVF, A, B, clk, reset, enable);
   output [63:0]Res;
   output OVF;
   input [31:0]A;
   input [31:0]B;
   input clk;
   input reset;
   input enable;

   wire [63:0]Res_imm;
   wire n_0_0__0;
   wire n_0_0__1;

   datapath__0_2 i_4 (.B_imm({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, 
      uc_8, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, 
      n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_0}), .A_imm({uc_9, 
      uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, n_46, n_24, n_25, n_26, 
      n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, 
      n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_1}), .Res_imm({uc_17, uc_18, 
      uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, 
      uc_29, uc_30, uc_31, uc_32, Res_imm[47], Res_imm[46], Res_imm[45], 
      Res_imm[44], Res_imm[43], Res_imm[42], Res_imm[41], Res_imm[40], 
      Res_imm[39], Res_imm[38], Res_imm[37], Res_imm[36], Res_imm[35], 
      Res_imm[34], Res_imm[33], Res_imm[32], Res_imm[31], Res_imm[30], 
      Res_imm[29], Res_imm[28], Res_imm[27], Res_imm[26], Res_imm[25], 
      Res_imm[24], Res_imm[23], uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, 
      uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49, 
      uc_50, uc_51, uc_52, uc_53, uc_54, uc_55}));
   DLH_X1 \Res_reg[47]  (.D(n_71), .G(n_119), .Q(Res[47]));
   DLH_X1 \Res_reg[46]  (.D(n_70), .G(n_119), .Q(Res[46]));
   DLH_X1 \Res_reg[45]  (.D(n_69), .G(n_119), .Q(Res[45]));
   DLH_X1 \Res_reg[44]  (.D(n_68), .G(n_119), .Q(Res[44]));
   DLH_X1 \Res_reg[43]  (.D(n_67), .G(n_119), .Q(Res[43]));
   DLH_X1 \Res_reg[42]  (.D(n_66), .G(n_119), .Q(Res[42]));
   DLH_X1 \Res_reg[41]  (.D(n_65), .G(n_119), .Q(Res[41]));
   DLH_X1 \Res_reg[40]  (.D(n_64), .G(n_119), .Q(Res[40]));
   DLH_X1 \Res_reg[39]  (.D(n_63), .G(n_119), .Q(Res[39]));
   DLH_X1 \Res_reg[38]  (.D(n_62), .G(n_119), .Q(Res[38]));
   DLH_X1 \Res_reg[37]  (.D(n_61), .G(n_119), .Q(Res[37]));
   DLH_X1 \Res_reg[36]  (.D(n_60), .G(n_119), .Q(Res[36]));
   DLH_X1 \Res_reg[35]  (.D(n_59), .G(n_119), .Q(Res[35]));
   DLH_X1 \Res_reg[34]  (.D(n_58), .G(n_119), .Q(Res[34]));
   DLH_X1 \Res_reg[33]  (.D(n_57), .G(n_119), .Q(Res[33]));
   DLH_X1 \Res_reg[32]  (.D(n_56), .G(n_119), .Q(Res[32]));
   DLH_X1 \Res_reg[31]  (.D(n_55), .G(n_119), .Q(Res[31]));
   DLH_X1 \Res_reg[30]  (.D(n_54), .G(n_119), .Q(Res[30]));
   DLH_X1 \Res_reg[29]  (.D(n_53), .G(n_119), .Q(Res[29]));
   DLH_X1 \Res_reg[28]  (.D(n_52), .G(n_119), .Q(Res[28]));
   DLH_X1 \Res_reg[27]  (.D(n_51), .G(n_119), .Q(Res[27]));
   DLH_X1 \Res_reg[26]  (.D(n_50), .G(n_119), .Q(Res[26]));
   DLH_X1 \Res_reg[25]  (.D(n_49), .G(n_119), .Q(Res[25]));
   DLH_X1 \Res_reg[24]  (.D(n_48), .G(n_119), .Q(Res[24]));
   DLH_X1 \Res_reg[23]  (.D(n_47), .G(n_119), .Q(Res[23]));
   DLH_X1 \B_in_reg[22]  (.D(n_118), .G(n_95), .Q(n_2));
   DLH_X1 \B_in_reg[21]  (.D(n_117), .G(n_95), .Q(n_3));
   DLH_X1 \B_in_reg[20]  (.D(n_116), .G(n_95), .Q(n_4));
   DLH_X1 \B_in_reg[19]  (.D(n_115), .G(n_95), .Q(n_5));
   DLH_X1 \B_in_reg[18]  (.D(n_114), .G(n_95), .Q(n_6));
   DLH_X1 \B_in_reg[17]  (.D(n_113), .G(n_95), .Q(n_7));
   DLH_X1 \B_in_reg[16]  (.D(n_112), .G(n_95), .Q(n_8));
   DLH_X1 \B_in_reg[15]  (.D(n_111), .G(n_95), .Q(n_9));
   DLH_X1 \B_in_reg[14]  (.D(n_110), .G(n_95), .Q(n_10));
   DLH_X1 \B_in_reg[13]  (.D(n_109), .G(n_95), .Q(n_11));
   DLH_X1 \B_in_reg[12]  (.D(n_108), .G(n_95), .Q(n_12));
   DLH_X1 \B_in_reg[11]  (.D(n_107), .G(n_95), .Q(n_13));
   DLH_X1 \B_in_reg[10]  (.D(n_106), .G(n_95), .Q(n_14));
   DLH_X1 \B_in_reg[9]  (.D(n_105), .G(n_95), .Q(n_15));
   DLH_X1 \B_in_reg[8]  (.D(n_104), .G(n_95), .Q(n_16));
   DLH_X1 \B_in_reg[7]  (.D(n_103), .G(n_95), .Q(n_17));
   DLH_X1 \B_in_reg[6]  (.D(n_102), .G(n_95), .Q(n_18));
   DLH_X1 \B_in_reg[5]  (.D(n_101), .G(n_95), .Q(n_19));
   DLH_X1 \B_in_reg[4]  (.D(n_100), .G(n_95), .Q(n_20));
   DLH_X1 \B_in_reg[3]  (.D(n_99), .G(n_95), .Q(n_21));
   DLH_X1 \B_in_reg[2]  (.D(n_98), .G(n_95), .Q(n_22));
   DLH_X1 \B_in_reg[1]  (.D(n_97), .G(n_95), .Q(n_23));
   DLH_X1 \B_in_reg[0]  (.D(n_96), .G(n_95), .Q(n_0));
   DLH_X1 \A_in_reg[22]  (.D(n_94), .G(n_95), .Q(n_24));
   DLH_X1 \A_in_reg[21]  (.D(n_93), .G(n_95), .Q(n_25));
   DLH_X1 \A_in_reg[20]  (.D(n_92), .G(n_95), .Q(n_26));
   DLH_X1 \A_in_reg[19]  (.D(n_91), .G(n_95), .Q(n_27));
   DLH_X1 \A_in_reg[18]  (.D(n_90), .G(n_95), .Q(n_28));
   DLH_X1 \A_in_reg[17]  (.D(n_89), .G(n_95), .Q(n_29));
   DLH_X1 \A_in_reg[16]  (.D(n_88), .G(n_95), .Q(n_30));
   DLH_X1 \A_in_reg[15]  (.D(n_87), .G(n_95), .Q(n_31));
   DLH_X1 \A_in_reg[14]  (.D(n_86), .G(n_95), .Q(n_32));
   DLH_X1 \A_in_reg[13]  (.D(n_85), .G(n_95), .Q(n_33));
   DLH_X1 \A_in_reg[12]  (.D(n_84), .G(n_95), .Q(n_34));
   DLH_X1 \A_in_reg[11]  (.D(n_83), .G(n_95), .Q(n_35));
   DLH_X1 \A_in_reg[10]  (.D(n_82), .G(n_95), .Q(n_36));
   DLH_X1 \A_in_reg[9]  (.D(n_81), .G(n_95), .Q(n_37));
   DLH_X1 \A_in_reg[8]  (.D(n_80), .G(n_95), .Q(n_38));
   DLH_X1 \A_in_reg[7]  (.D(n_79), .G(n_95), .Q(n_39));
   DLH_X1 \A_in_reg[6]  (.D(n_78), .G(n_95), .Q(n_40));
   DLH_X1 \A_in_reg[5]  (.D(n_77), .G(n_95), .Q(n_41));
   DLH_X1 \A_in_reg[4]  (.D(n_76), .G(n_95), .Q(n_42));
   DLH_X1 \A_in_reg[3]  (.D(n_75), .G(n_95), .Q(n_43));
   DLH_X1 \A_in_reg[2]  (.D(n_74), .G(n_95), .Q(n_44));
   DLH_X1 \A_in_reg[1]  (.D(n_73), .G(n_95), .Q(n_45));
   DLH_X1 \A_in_reg[0]  (.D(n_72), .G(n_95), .Q(n_1));
   DLH_X1 \A_in_reg[23]  (.D(n_0_0__1), .G(n_95), .Q(n_46));
   AND2_X1 i_0_0 (.A1(n_0_0__1), .A2(Res_imm[23]), .ZN(n_47));
   AND2_X1 i_0_1 (.A1(n_0_0__1), .A2(Res_imm[24]), .ZN(n_48));
   AND2_X1 i_0_2 (.A1(n_0_0__1), .A2(Res_imm[25]), .ZN(n_49));
   AND2_X1 i_0_3 (.A1(n_0_0__1), .A2(Res_imm[26]), .ZN(n_50));
   AND2_X1 i_0_4 (.A1(n_0_0__1), .A2(Res_imm[27]), .ZN(n_51));
   AND2_X1 i_0_5 (.A1(n_0_0__1), .A2(Res_imm[28]), .ZN(n_52));
   AND2_X1 i_0_6 (.A1(n_0_0__1), .A2(Res_imm[29]), .ZN(n_53));
   AND2_X1 i_0_7 (.A1(n_0_0__1), .A2(Res_imm[30]), .ZN(n_54));
   AND2_X1 i_0_8 (.A1(n_0_0__1), .A2(Res_imm[31]), .ZN(n_55));
   AND2_X1 i_0_9 (.A1(n_0_0__1), .A2(Res_imm[32]), .ZN(n_56));
   AND2_X1 i_0_10 (.A1(n_0_0__1), .A2(Res_imm[33]), .ZN(n_57));
   AND2_X1 i_0_11 (.A1(n_0_0__1), .A2(Res_imm[34]), .ZN(n_58));
   AND2_X1 i_0_12 (.A1(n_0_0__1), .A2(Res_imm[35]), .ZN(n_59));
   AND2_X1 i_0_13 (.A1(n_0_0__1), .A2(Res_imm[36]), .ZN(n_60));
   AND2_X1 i_0_14 (.A1(n_0_0__1), .A2(Res_imm[37]), .ZN(n_61));
   AND2_X1 i_0_15 (.A1(n_0_0__1), .A2(Res_imm[38]), .ZN(n_62));
   AND2_X1 i_0_16 (.A1(n_0_0__1), .A2(Res_imm[39]), .ZN(n_63));
   AND2_X1 i_0_17 (.A1(n_0_0__1), .A2(Res_imm[40]), .ZN(n_64));
   AND2_X1 i_0_18 (.A1(n_0_0__1), .A2(Res_imm[41]), .ZN(n_65));
   AND2_X1 i_0_19 (.A1(n_0_0__1), .A2(Res_imm[42]), .ZN(n_66));
   AND2_X1 i_0_20 (.A1(n_0_0__1), .A2(Res_imm[43]), .ZN(n_67));
   AND2_X1 i_0_21 (.A1(n_0_0__1), .A2(Res_imm[44]), .ZN(n_68));
   AND2_X1 i_0_22 (.A1(n_0_0__1), .A2(Res_imm[45]), .ZN(n_69));
   AND2_X1 i_0_23 (.A1(n_0_0__1), .A2(Res_imm[46]), .ZN(n_70));
   AND2_X1 i_0_24 (.A1(n_0_0__1), .A2(Res_imm[47]), .ZN(n_71));
   AND2_X1 i_0_25 (.A1(n_0_0__1), .A2(A[0]), .ZN(n_72));
   AND2_X1 i_0_26 (.A1(n_0_0__1), .A2(A[1]), .ZN(n_73));
   AND2_X1 i_0_27 (.A1(n_0_0__1), .A2(A[2]), .ZN(n_74));
   AND2_X1 i_0_28 (.A1(n_0_0__1), .A2(A[3]), .ZN(n_75));
   AND2_X1 i_0_29 (.A1(n_0_0__1), .A2(A[4]), .ZN(n_76));
   AND2_X1 i_0_30 (.A1(n_0_0__1), .A2(A[5]), .ZN(n_77));
   AND2_X1 i_0_31 (.A1(n_0_0__1), .A2(A[6]), .ZN(n_78));
   AND2_X1 i_0_32 (.A1(n_0_0__1), .A2(A[7]), .ZN(n_79));
   AND2_X1 i_0_33 (.A1(n_0_0__1), .A2(A[8]), .ZN(n_80));
   AND2_X1 i_0_34 (.A1(n_0_0__1), .A2(A[9]), .ZN(n_81));
   AND2_X1 i_0_35 (.A1(n_0_0__1), .A2(A[10]), .ZN(n_82));
   AND2_X1 i_0_36 (.A1(n_0_0__1), .A2(A[11]), .ZN(n_83));
   AND2_X1 i_0_37 (.A1(n_0_0__1), .A2(A[12]), .ZN(n_84));
   AND2_X1 i_0_38 (.A1(n_0_0__1), .A2(A[13]), .ZN(n_85));
   AND2_X1 i_0_39 (.A1(n_0_0__1), .A2(A[14]), .ZN(n_86));
   AND2_X1 i_0_40 (.A1(n_0_0__1), .A2(A[15]), .ZN(n_87));
   AND2_X1 i_0_41 (.A1(n_0_0__1), .A2(A[16]), .ZN(n_88));
   AND2_X1 i_0_42 (.A1(n_0_0__1), .A2(A[17]), .ZN(n_89));
   AND2_X1 i_0_43 (.A1(n_0_0__1), .A2(A[18]), .ZN(n_90));
   AND2_X1 i_0_44 (.A1(n_0_0__1), .A2(A[19]), .ZN(n_91));
   AND2_X1 i_0_45 (.A1(n_0_0__1), .A2(A[20]), .ZN(n_92));
   AND2_X1 i_0_46 (.A1(n_0_0__1), .A2(A[21]), .ZN(n_93));
   AND2_X1 i_0_47 (.A1(n_0_0__1), .A2(A[22]), .ZN(n_94));
   INV_X1 i_0_48 (.A(n_0_0__0), .ZN(n_95));
   AOI21_X1 i_0_49 (.A(reset), .B1(clk), .B2(enable), .ZN(n_0_0__0));
   AND2_X1 i_0_50 (.A1(n_0_0__1), .A2(B[0]), .ZN(n_96));
   AND2_X1 i_0_51 (.A1(n_0_0__1), .A2(B[1]), .ZN(n_97));
   AND2_X1 i_0_52 (.A1(n_0_0__1), .A2(B[2]), .ZN(n_98));
   AND2_X1 i_0_53 (.A1(n_0_0__1), .A2(B[3]), .ZN(n_99));
   AND2_X1 i_0_54 (.A1(n_0_0__1), .A2(B[4]), .ZN(n_100));
   AND2_X1 i_0_55 (.A1(n_0_0__1), .A2(B[5]), .ZN(n_101));
   AND2_X1 i_0_56 (.A1(n_0_0__1), .A2(B[6]), .ZN(n_102));
   AND2_X1 i_0_57 (.A1(n_0_0__1), .A2(B[7]), .ZN(n_103));
   AND2_X1 i_0_58 (.A1(n_0_0__1), .A2(B[8]), .ZN(n_104));
   AND2_X1 i_0_59 (.A1(n_0_0__1), .A2(B[9]), .ZN(n_105));
   AND2_X1 i_0_60 (.A1(n_0_0__1), .A2(B[10]), .ZN(n_106));
   AND2_X1 i_0_61 (.A1(n_0_0__1), .A2(B[11]), .ZN(n_107));
   AND2_X1 i_0_62 (.A1(n_0_0__1), .A2(B[12]), .ZN(n_108));
   AND2_X1 i_0_63 (.A1(n_0_0__1), .A2(B[13]), .ZN(n_109));
   AND2_X1 i_0_64 (.A1(n_0_0__1), .A2(B[14]), .ZN(n_110));
   AND2_X1 i_0_65 (.A1(n_0_0__1), .A2(B[15]), .ZN(n_111));
   AND2_X1 i_0_66 (.A1(n_0_0__1), .A2(B[16]), .ZN(n_112));
   AND2_X1 i_0_67 (.A1(n_0_0__1), .A2(B[17]), .ZN(n_113));
   AND2_X1 i_0_68 (.A1(n_0_0__1), .A2(B[18]), .ZN(n_114));
   AND2_X1 i_0_69 (.A1(n_0_0__1), .A2(B[19]), .ZN(n_115));
   AND2_X1 i_0_70 (.A1(n_0_0__1), .A2(B[20]), .ZN(n_116));
   AND2_X1 i_0_71 (.A1(n_0_0__1), .A2(B[21]), .ZN(n_117));
   AND2_X1 i_0_72 (.A1(n_0_0__1), .A2(B[22]), .ZN(n_118));
   NAND2_X1 i_0_73 (.A1(n_0_0__1), .A2(clk), .ZN(n_119));
   INV_X1 i_0_74 (.A(reset), .ZN(n_0_0__1));
endmodule

module datapath__0_13(M_multiplied, p_0, M_resultTruncated);
   input M_multiplied;
   input [22:0]p_0;
   output [22:0]M_resultTruncated;

   HA_X1 i_0 (.A(M_multiplied), .B(p_0[0]), .CO(n_0), .S(M_resultTruncated[0]));
   HA_X1 i_1 (.A(p_0[1]), .B(n_0), .CO(n_1), .S(M_resultTruncated[1]));
   HA_X1 i_2 (.A(p_0[2]), .B(n_1), .CO(n_2), .S(M_resultTruncated[2]));
   HA_X1 i_3 (.A(p_0[3]), .B(n_2), .CO(n_3), .S(M_resultTruncated[3]));
   HA_X1 i_4 (.A(p_0[4]), .B(n_3), .CO(n_4), .S(M_resultTruncated[4]));
   HA_X1 i_5 (.A(p_0[5]), .B(n_4), .CO(n_5), .S(M_resultTruncated[5]));
   HA_X1 i_6 (.A(p_0[6]), .B(n_5), .CO(n_6), .S(M_resultTruncated[6]));
   HA_X1 i_7 (.A(p_0[7]), .B(n_6), .CO(n_7), .S(M_resultTruncated[7]));
   HA_X1 i_8 (.A(p_0[8]), .B(n_7), .CO(n_8), .S(M_resultTruncated[8]));
   HA_X1 i_9 (.A(p_0[9]), .B(n_8), .CO(n_9), .S(M_resultTruncated[9]));
   HA_X1 i_10 (.A(p_0[10]), .B(n_9), .CO(n_10), .S(M_resultTruncated[10]));
   HA_X1 i_11 (.A(p_0[11]), .B(n_10), .CO(n_11), .S(M_resultTruncated[11]));
   HA_X1 i_12 (.A(p_0[12]), .B(n_11), .CO(n_12), .S(M_resultTruncated[12]));
   HA_X1 i_13 (.A(p_0[13]), .B(n_12), .CO(n_13), .S(M_resultTruncated[13]));
   HA_X1 i_14 (.A(p_0[14]), .B(n_13), .CO(n_14), .S(M_resultTruncated[14]));
   HA_X1 i_15 (.A(p_0[15]), .B(n_14), .CO(n_15), .S(M_resultTruncated[15]));
   HA_X1 i_16 (.A(p_0[16]), .B(n_15), .CO(n_16), .S(M_resultTruncated[16]));
   HA_X1 i_17 (.A(p_0[17]), .B(n_16), .CO(n_17), .S(M_resultTruncated[17]));
   HA_X1 i_18 (.A(p_0[18]), .B(n_17), .CO(n_18), .S(M_resultTruncated[18]));
   HA_X1 i_19 (.A(p_0[19]), .B(n_18), .CO(n_19), .S(M_resultTruncated[19]));
   HA_X1 i_20 (.A(p_0[20]), .B(n_19), .CO(n_20), .S(M_resultTruncated[20]));
   HA_X1 i_21 (.A(p_0[21]), .B(n_20), .CO(n_21), .S(M_resultTruncated[21]));
   XOR2_X1 i_22 (.A(p_0[22]), .B(n_21), .Z(M_resultTruncated[22]));
endmodule

module FPU_VM(Res, A, B, clk, reset, enable);
   output [31:0]Res;
   input [31:0]A;
   input [31:0]B;
   input clk;
   input reset;
   input enable;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire [22:0]M_resultTruncated;
   wire [7:0]EA;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire [7:0]EB;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire A_reg;
   wire B_reg;
   wire n_0_1_2;
   wire n_0_1_3;
   wire n_0_1_4;
   wire n_0_1_5;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_1_8;
   wire n_0_1_9;
   wire n_0_1_10;
   wire n_0_1_11;
   wire n_0_1_12;
   wire n_0_1_13;
   wire n_0_1_14;
   wire n_0_1_15;
   wire n_0_1_22;
   wire n_0_1_16;
   wire n_0_1_23;
   wire n_0_1_17;
   wire n_0_1_24;
   wire n_0_1_18;
   wire n_0_1_25;
   wire n_0_1_19;
   wire n_0_1_26;
   wire n_0_1_20;
   wire n_0_1_27;
   wire n_0_1_21;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_72;
   wire n_0_1_32;
   wire n_0_73;
   wire n_0_1_33;
   wire n_0_74;
   wire n_0_1_34;
   wire n_0_75;
   wire n_0_1_35;
   wire n_0_76;
   wire n_0_1_36;
   wire n_0_77;
   wire n_0_1_37;
   wire n_0_78;
   wire n_0_1_38;
   wire n_0_79;
   wire n_0_1_39;
   wire n_0_80;
   wire n_0_1_40;
   wire n_0_81;
   wire n_0_1_41;
   wire n_0_82;
   wire n_0_1_42;
   wire n_0_83;
   wire n_0_1_43;
   wire n_0_84;
   wire n_0_1_44;
   wire n_0_85;
   wire n_0_1_45;
   wire n_0_86;
   wire n_0_1_46;
   wire n_0_87;
   wire n_0_1_47;
   wire n_0_88;
   wire n_0_1_48;
   wire n_0_89;
   wire n_0_1_49;
   wire n_0_90;
   wire n_0_1_50;
   wire n_0_91;
   wire n_0_1_51;
   wire n_0_92;
   wire n_0_1_52;
   wire n_0_93;
   wire n_0_1_53;
   wire n_0_1_54;
   wire n_0_1_55;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_1_56;
   wire n_0_1_57;
   wire n_0_1_58;
   wire n_0_1_59;
   wire n_0_1_60;
   wire n_0_1_62;
   wire n_0_1_64;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_1_105;
   wire n_0_1_106;
   wire n_0_1_107;
   wire n_0_1_108;
   wire n_0_1_109;
   wire n_0_1_110;
   wire n_0_1_111;
   wire n_0_1_112;
   wire n_0_1_28;
   wire n_0_1_29;
   wire n_0_71;
   wire n_0_1_30;
   wire n_0_1_31;
   wire n_0_1_61;
   wire n_0_1_63;
   wire n_0_1_65;
   wire n_0_1_66;
   wire n_0_1_67;
   wire n_0_1_68;
   wire n_0_1_69;
   wire n_0_1_70;
   wire n_0_1_71;
   wire n_0_1_72;
   wire n_0_1_73;
   wire n_0_1_74;
   wire n_0_1_75;
   wire n_0_1_76;
   wire n_0_1_77;
   wire n_0_1_78;
   wire n_0_1_79;
   wire n_0_1_80;
   wire n_0_1_81;
   wire n_0_1_82;
   wire n_0_1_83;
   wire n_0_1_84;
   wire n_0_1_85;
   wire n_0_1_86;
   wire n_0_1_87;
   wire n_0_1_88;
   wire n_0_1_89;
   wire n_0_1_90;
   wire n_0_1_91;
   wire n_0_1_92;
   wire n_0_1_93;
   wire n_0_1_94;
   wire n_0_1_95;
   wire n_0_1_96;
   wire n_0_1_97;
   wire n_0_1_98;
   wire n_0_1_99;
   wire n_0_1_100;
   wire n_0_1_101;
   wire n_0_1_102;
   wire n_0_1_103;
   wire n_0_102;
   wire n_0_1_104;

   VM multiplier (.Res({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, 
      uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, n_0_24, n_0_23, n_0_22, 
      n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, 
      n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, 
      n_0_2, n_0_1, n_0_0, uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, 
      uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, uc_32, 
      uc_33, uc_34, uc_35, uc_36, uc_37, uc_38}), .OVF(), .A({uc_39, uc_40, 
      uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, n_0_25, n_0_26, n_0_27, 
      n_0_28, n_0_29, n_0_30, n_0_31, n_0_32, n_0_33, n_0_34, n_0_35, n_0_36, 
      n_0_37, n_0_38, n_0_39, n_0_40, n_0_41, n_0_42, n_0_43, n_0_44, n_0_45, 
      n_0_46, n_0_47}), .B({uc_48, uc_49, uc_50, uc_51, uc_52, uc_53, uc_54, 
      uc_55, uc_56, n_0_48, n_0_49, n_0_50, n_0_51, n_0_52, n_0_53, n_0_54, 
      n_0_55, n_0_56, n_0_57, n_0_58, n_0_59, n_0_60, n_0_61, n_0_62, n_0_63, 
      n_0_64, n_0_65, n_0_66, n_0_67, n_0_68, n_0_69, n_0_70}), .clk(clk), 
      .reset(reset), .enable(enable));
   datapath__0_13 i_0_0 (.M_multiplied(n_0_0), .p_0({n_0_23, n_0_22, n_0_21, 
      n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, 
      n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, 
      n_0_1}), .M_resultTruncated(M_resultTruncated));
   DLH_X1 \Res_reg[31]  (.D(n_0_102), .G(n_0_168), .Q(Res[31]));
   DLH_X1 \Res_reg[30]  (.D(n_0_101), .G(n_0_168), .Q(Res[30]));
   DLH_X1 \Res_reg[29]  (.D(n_0_100), .G(n_0_168), .Q(Res[29]));
   DLH_X1 \Res_reg[28]  (.D(n_0_99), .G(n_0_168), .Q(Res[28]));
   DLH_X1 \Res_reg[27]  (.D(n_0_98), .G(n_0_168), .Q(Res[27]));
   DLH_X1 \Res_reg[26]  (.D(n_0_97), .G(n_0_168), .Q(Res[26]));
   DLH_X1 \Res_reg[25]  (.D(n_0_96), .G(n_0_168), .Q(Res[25]));
   DLH_X1 \Res_reg[24]  (.D(n_0_95), .G(n_0_168), .Q(Res[24]));
   DLH_X1 \Res_reg[23]  (.D(n_0_94), .G(n_0_168), .Q(Res[23]));
   DLH_X1 \Res_reg[22]  (.D(n_0_93), .G(n_0_168), .Q(Res[22]));
   DLH_X1 \Res_reg[21]  (.D(n_0_92), .G(n_0_168), .Q(Res[21]));
   DLH_X1 \Res_reg[20]  (.D(n_0_91), .G(n_0_168), .Q(Res[20]));
   DLH_X1 \Res_reg[19]  (.D(n_0_90), .G(n_0_168), .Q(Res[19]));
   DLH_X1 \Res_reg[18]  (.D(n_0_89), .G(n_0_168), .Q(Res[18]));
   DLH_X1 \Res_reg[17]  (.D(n_0_88), .G(n_0_168), .Q(Res[17]));
   DLH_X1 \Res_reg[16]  (.D(n_0_87), .G(n_0_168), .Q(Res[16]));
   DLH_X1 \Res_reg[15]  (.D(n_0_86), .G(n_0_168), .Q(Res[15]));
   DLH_X1 \Res_reg[14]  (.D(n_0_85), .G(n_0_168), .Q(Res[14]));
   DLH_X1 \Res_reg[13]  (.D(n_0_84), .G(n_0_168), .Q(Res[13]));
   DLH_X1 \Res_reg[12]  (.D(n_0_83), .G(n_0_168), .Q(Res[12]));
   DLH_X1 \Res_reg[11]  (.D(n_0_82), .G(n_0_168), .Q(Res[11]));
   DLH_X1 \Res_reg[10]  (.D(n_0_81), .G(n_0_168), .Q(Res[10]));
   DLH_X1 \Res_reg[9]  (.D(n_0_80), .G(n_0_168), .Q(Res[9]));
   DLH_X1 \Res_reg[8]  (.D(n_0_79), .G(n_0_168), .Q(Res[8]));
   DLH_X1 \Res_reg[7]  (.D(n_0_78), .G(n_0_168), .Q(Res[7]));
   DLH_X1 \Res_reg[6]  (.D(n_0_77), .G(n_0_168), .Q(Res[6]));
   DLH_X1 \Res_reg[5]  (.D(n_0_76), .G(n_0_168), .Q(Res[5]));
   DLH_X1 \Res_reg[4]  (.D(n_0_75), .G(n_0_168), .Q(Res[4]));
   DLH_X1 \Res_reg[3]  (.D(n_0_74), .G(n_0_168), .Q(Res[3]));
   DLH_X1 \Res_reg[2]  (.D(n_0_73), .G(n_0_168), .Q(Res[2]));
   DLH_X1 \Res_reg[1]  (.D(n_0_72), .G(n_0_168), .Q(Res[1]));
   DLH_X1 \Res_reg[0]  (.D(n_0_71), .G(n_0_168), .Q(Res[0]));
   DLH_X1 \A_reg_reg[30]  (.D(n_0_136), .G(n_0_104), .Q(EA[7]));
   DLH_X1 \A_reg_reg[29]  (.D(n_0_135), .G(n_0_104), .Q(EA[6]));
   DLH_X1 \A_reg_reg[28]  (.D(n_0_134), .G(n_0_104), .Q(EA[5]));
   DLH_X1 \A_reg_reg[27]  (.D(n_0_133), .G(n_0_104), .Q(EA[4]));
   DLH_X1 \A_reg_reg[26]  (.D(n_0_132), .G(n_0_104), .Q(EA[3]));
   DLH_X1 \A_reg_reg[25]  (.D(n_0_131), .G(n_0_104), .Q(EA[2]));
   DLH_X1 \A_reg_reg[24]  (.D(n_0_130), .G(n_0_104), .Q(EA[1]));
   DLH_X1 \A_reg_reg[23]  (.D(n_0_129), .G(n_0_104), .Q(EA[0]));
   DLH_X1 \A_reg_reg[22]  (.D(n_0_128), .G(n_0_104), .Q(n_0_25));
   DLH_X1 \A_reg_reg[21]  (.D(n_0_127), .G(n_0_104), .Q(n_0_26));
   DLH_X1 \A_reg_reg[20]  (.D(n_0_126), .G(n_0_104), .Q(n_0_27));
   DLH_X1 \A_reg_reg[19]  (.D(n_0_125), .G(n_0_104), .Q(n_0_28));
   DLH_X1 \A_reg_reg[18]  (.D(n_0_124), .G(n_0_104), .Q(n_0_29));
   DLH_X1 \A_reg_reg[17]  (.D(n_0_123), .G(n_0_104), .Q(n_0_30));
   DLH_X1 \A_reg_reg[16]  (.D(n_0_122), .G(n_0_104), .Q(n_0_31));
   DLH_X1 \A_reg_reg[15]  (.D(n_0_121), .G(n_0_104), .Q(n_0_32));
   DLH_X1 \A_reg_reg[14]  (.D(n_0_120), .G(n_0_104), .Q(n_0_33));
   DLH_X1 \A_reg_reg[13]  (.D(n_0_119), .G(n_0_104), .Q(n_0_34));
   DLH_X1 \A_reg_reg[12]  (.D(n_0_118), .G(n_0_104), .Q(n_0_35));
   DLH_X1 \A_reg_reg[11]  (.D(n_0_117), .G(n_0_104), .Q(n_0_36));
   DLH_X1 \A_reg_reg[10]  (.D(n_0_116), .G(n_0_104), .Q(n_0_37));
   DLH_X1 \A_reg_reg[9]  (.D(n_0_115), .G(n_0_104), .Q(n_0_38));
   DLH_X1 \A_reg_reg[8]  (.D(n_0_114), .G(n_0_104), .Q(n_0_39));
   DLH_X1 \A_reg_reg[7]  (.D(n_0_113), .G(n_0_104), .Q(n_0_40));
   DLH_X1 \A_reg_reg[6]  (.D(n_0_112), .G(n_0_104), .Q(n_0_41));
   DLH_X1 \A_reg_reg[5]  (.D(n_0_111), .G(n_0_104), .Q(n_0_42));
   DLH_X1 \A_reg_reg[4]  (.D(n_0_110), .G(n_0_104), .Q(n_0_43));
   DLH_X1 \A_reg_reg[3]  (.D(n_0_109), .G(n_0_104), .Q(n_0_44));
   DLH_X1 \A_reg_reg[2]  (.D(n_0_108), .G(n_0_104), .Q(n_0_45));
   DLH_X1 \A_reg_reg[1]  (.D(n_0_107), .G(n_0_104), .Q(n_0_46));
   DLH_X1 \A_reg_reg[0]  (.D(n_0_106), .G(n_0_104), .Q(n_0_47));
   DLH_X1 \B_reg_reg[30]  (.D(n_0_167), .G(n_0_104), .Q(EB[7]));
   DLH_X1 \B_reg_reg[29]  (.D(n_0_166), .G(n_0_104), .Q(EB[6]));
   DLH_X1 \B_reg_reg[28]  (.D(n_0_165), .G(n_0_104), .Q(EB[5]));
   DLH_X1 \B_reg_reg[27]  (.D(n_0_164), .G(n_0_104), .Q(EB[4]));
   DLH_X1 \B_reg_reg[26]  (.D(n_0_163), .G(n_0_104), .Q(EB[3]));
   DLH_X1 \B_reg_reg[25]  (.D(n_0_162), .G(n_0_104), .Q(EB[2]));
   DLH_X1 \B_reg_reg[24]  (.D(n_0_161), .G(n_0_104), .Q(EB[1]));
   DLH_X1 \B_reg_reg[23]  (.D(n_0_160), .G(n_0_104), .Q(EB[0]));
   DLH_X1 \B_reg_reg[22]  (.D(n_0_159), .G(n_0_104), .Q(n_0_48));
   DLH_X1 \B_reg_reg[21]  (.D(n_0_158), .G(n_0_104), .Q(n_0_49));
   DLH_X1 \B_reg_reg[20]  (.D(n_0_157), .G(n_0_104), .Q(n_0_50));
   DLH_X1 \B_reg_reg[19]  (.D(n_0_156), .G(n_0_104), .Q(n_0_51));
   DLH_X1 \B_reg_reg[18]  (.D(n_0_155), .G(n_0_104), .Q(n_0_52));
   DLH_X1 \B_reg_reg[17]  (.D(n_0_154), .G(n_0_104), .Q(n_0_53));
   DLH_X1 \B_reg_reg[16]  (.D(n_0_153), .G(n_0_104), .Q(n_0_54));
   DLH_X1 \B_reg_reg[15]  (.D(n_0_152), .G(n_0_104), .Q(n_0_55));
   DLH_X1 \B_reg_reg[14]  (.D(n_0_151), .G(n_0_104), .Q(n_0_56));
   DLH_X1 \B_reg_reg[13]  (.D(n_0_150), .G(n_0_104), .Q(n_0_57));
   DLH_X1 \B_reg_reg[12]  (.D(n_0_149), .G(n_0_104), .Q(n_0_58));
   DLH_X1 \B_reg_reg[11]  (.D(n_0_148), .G(n_0_104), .Q(n_0_59));
   DLH_X1 \B_reg_reg[10]  (.D(n_0_147), .G(n_0_104), .Q(n_0_60));
   DLH_X1 \B_reg_reg[9]  (.D(n_0_146), .G(n_0_104), .Q(n_0_61));
   DLH_X1 \B_reg_reg[8]  (.D(n_0_145), .G(n_0_104), .Q(n_0_62));
   DLH_X1 \B_reg_reg[7]  (.D(n_0_144), .G(n_0_104), .Q(n_0_63));
   DLH_X1 \B_reg_reg[6]  (.D(n_0_143), .G(n_0_104), .Q(n_0_64));
   DLH_X1 \B_reg_reg[5]  (.D(n_0_142), .G(n_0_104), .Q(n_0_65));
   DLH_X1 \B_reg_reg[4]  (.D(n_0_141), .G(n_0_104), .Q(n_0_66));
   DLH_X1 \B_reg_reg[3]  (.D(n_0_140), .G(n_0_104), .Q(n_0_67));
   DLH_X1 \B_reg_reg[2]  (.D(n_0_139), .G(n_0_104), .Q(n_0_68));
   DLH_X1 \B_reg_reg[1]  (.D(n_0_138), .G(n_0_104), .Q(n_0_69));
   DLH_X1 \B_reg_reg[0]  (.D(n_0_137), .G(n_0_104), .Q(n_0_70));
   DLH_X1 \A_reg_reg[31]  (.D(n_0_103), .G(n_0_104), .Q(A_reg));
   DLH_X1 \B_reg_reg[31]  (.D(n_0_105), .G(n_0_104), .Q(B_reg));
   HA_X1 i_0_1_0 (.A(EB[1]), .B(EA[1]), .CO(n_0_1_3), .S(n_0_1_2));
   HA_X1 i_0_1_1 (.A(EB[2]), .B(EA[2]), .CO(n_0_1_5), .S(n_0_1_4));
   HA_X1 i_0_1_2 (.A(EB[3]), .B(EA[3]), .CO(n_0_1_7), .S(n_0_1_6));
   HA_X1 i_0_1_3 (.A(EB[4]), .B(EA[4]), .CO(n_0_1_9), .S(n_0_1_8));
   HA_X1 i_0_1_4 (.A(EB[5]), .B(EA[5]), .CO(n_0_1_11), .S(n_0_1_10));
   HA_X1 i_0_1_5 (.A(EB[6]), .B(EA[6]), .CO(n_0_1_13), .S(n_0_1_12));
   HA_X1 i_0_1_6 (.A(EA[0]), .B(n_0_1_0), .CO(n_0_1_15), .S(n_0_1_14));
   FA_X1 i_0_1_7 (.A(n_0_1_1), .B(n_0_1_2), .CI(n_0_1_15), .CO(n_0_1_16), 
      .S(n_0_1_22));
   FA_X1 i_0_1_8 (.A(n_0_1_3), .B(n_0_1_4), .CI(n_0_1_16), .CO(n_0_1_17), 
      .S(n_0_1_23));
   FA_X1 i_0_1_9 (.A(n_0_1_5), .B(n_0_1_6), .CI(n_0_1_17), .CO(n_0_1_18), 
      .S(n_0_1_24));
   FA_X1 i_0_1_10 (.A(n_0_1_7), .B(n_0_1_8), .CI(n_0_1_18), .CO(n_0_1_19), 
      .S(n_0_1_25));
   FA_X1 i_0_1_11 (.A(n_0_1_9), .B(n_0_1_10), .CI(n_0_1_19), .CO(n_0_1_20), 
      .S(n_0_1_26));
   FA_X1 i_0_1_12 (.A(n_0_1_11), .B(n_0_1_12), .CI(n_0_1_20), .CO(n_0_1_21), 
      .S(n_0_1_27));
   XNOR2_X1 i_0_1_13 (.A(EB[0]), .B(n_0_24), .ZN(n_0_1_0));
   OR2_X1 i_0_1_14 (.A1(EB[0]), .A2(n_0_24), .ZN(n_0_1_1));
   INV_X1 i_0_1_15 (.A(n_0_1_32), .ZN(n_0_72));
   AOI22_X1 i_0_1_16 (.A1(M_resultTruncated[1]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_1), .ZN(n_0_1_32));
   INV_X1 i_0_1_22 (.A(n_0_1_33), .ZN(n_0_73));
   AOI22_X1 i_0_1_23 (.A1(M_resultTruncated[2]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_2), .ZN(n_0_1_33));
   INV_X1 i_0_1_24 (.A(n_0_1_34), .ZN(n_0_74));
   AOI22_X1 i_0_1_25 (.A1(M_resultTruncated[3]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_3), .ZN(n_0_1_34));
   INV_X1 i_0_1_26 (.A(n_0_1_35), .ZN(n_0_75));
   AOI22_X1 i_0_1_27 (.A1(M_resultTruncated[4]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_4), .ZN(n_0_1_35));
   INV_X1 i_0_1_28 (.A(n_0_1_36), .ZN(n_0_76));
   AOI22_X1 i_0_1_29 (.A1(M_resultTruncated[5]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_5), .ZN(n_0_1_36));
   INV_X1 i_0_1_30 (.A(n_0_1_37), .ZN(n_0_77));
   AOI22_X1 i_0_1_31 (.A1(M_resultTruncated[6]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_6), .ZN(n_0_1_37));
   INV_X1 i_0_1_32 (.A(n_0_1_38), .ZN(n_0_78));
   AOI22_X1 i_0_1_33 (.A1(M_resultTruncated[7]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_7), .ZN(n_0_1_38));
   INV_X1 i_0_1_34 (.A(n_0_1_39), .ZN(n_0_79));
   AOI22_X1 i_0_1_35 (.A1(M_resultTruncated[8]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_8), .ZN(n_0_1_39));
   INV_X1 i_0_1_36 (.A(n_0_1_40), .ZN(n_0_80));
   AOI22_X1 i_0_1_37 (.A1(M_resultTruncated[9]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_9), .ZN(n_0_1_40));
   INV_X1 i_0_1_38 (.A(n_0_1_41), .ZN(n_0_81));
   AOI22_X1 i_0_1_39 (.A1(M_resultTruncated[10]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_10), .ZN(n_0_1_41));
   INV_X1 i_0_1_40 (.A(n_0_1_42), .ZN(n_0_82));
   AOI22_X1 i_0_1_41 (.A1(M_resultTruncated[11]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_11), .ZN(n_0_1_42));
   INV_X1 i_0_1_42 (.A(n_0_1_43), .ZN(n_0_83));
   AOI22_X1 i_0_1_43 (.A1(M_resultTruncated[12]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_12), .ZN(n_0_1_43));
   INV_X1 i_0_1_44 (.A(n_0_1_44), .ZN(n_0_84));
   AOI22_X1 i_0_1_45 (.A1(M_resultTruncated[13]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_13), .ZN(n_0_1_44));
   INV_X1 i_0_1_46 (.A(n_0_1_45), .ZN(n_0_85));
   AOI22_X1 i_0_1_47 (.A1(M_resultTruncated[14]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_14), .ZN(n_0_1_45));
   INV_X1 i_0_1_48 (.A(n_0_1_46), .ZN(n_0_86));
   AOI22_X1 i_0_1_49 (.A1(M_resultTruncated[15]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_15), .ZN(n_0_1_46));
   INV_X1 i_0_1_50 (.A(n_0_1_47), .ZN(n_0_87));
   AOI22_X1 i_0_1_51 (.A1(M_resultTruncated[16]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_16), .ZN(n_0_1_47));
   INV_X1 i_0_1_52 (.A(n_0_1_48), .ZN(n_0_88));
   AOI22_X1 i_0_1_53 (.A1(M_resultTruncated[17]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_17), .ZN(n_0_1_48));
   INV_X1 i_0_1_54 (.A(n_0_1_49), .ZN(n_0_89));
   AOI22_X1 i_0_1_55 (.A1(M_resultTruncated[18]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_18), .ZN(n_0_1_49));
   INV_X1 i_0_1_56 (.A(n_0_1_50), .ZN(n_0_90));
   AOI22_X1 i_0_1_57 (.A1(M_resultTruncated[19]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_19), .ZN(n_0_1_50));
   INV_X1 i_0_1_58 (.A(n_0_1_51), .ZN(n_0_91));
   AOI22_X1 i_0_1_59 (.A1(M_resultTruncated[20]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_20), .ZN(n_0_1_51));
   INV_X1 i_0_1_60 (.A(n_0_1_52), .ZN(n_0_92));
   AOI22_X1 i_0_1_61 (.A1(M_resultTruncated[21]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_21), .ZN(n_0_1_52));
   INV_X1 i_0_1_62 (.A(n_0_1_53), .ZN(n_0_93));
   AOI22_X1 i_0_1_63 (.A1(M_resultTruncated[22]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_0_22), .ZN(n_0_1_53));
   NOR3_X1 i_0_1_17 (.A1(n_0_1_60), .A2(n_0_24), .A3(n_0_1_64), .ZN(n_0_1_54));
   NOR3_X1 i_0_1_18 (.A1(n_0_1_29), .A2(n_0_1_64), .A3(n_0_1_60), .ZN(n_0_1_55));
   OAI21_X1 i_0_1_19 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_111), .ZN(n_0_94));
   OAI21_X1 i_0_1_67 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_110), .ZN(n_0_95));
   OAI21_X1 i_0_1_68 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_109), .ZN(n_0_96));
   OAI21_X1 i_0_1_69 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_108), .ZN(n_0_97));
   OAI21_X1 i_0_1_70 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_107), .ZN(n_0_98));
   OAI21_X1 i_0_1_71 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_106), .ZN(n_0_99));
   OAI21_X1 i_0_1_72 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_105), .ZN(n_0_100));
   OAI21_X1 i_0_1_73 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_56), .ZN(n_0_101));
   XNOR2_X1 i_0_1_74 (.A(n_0_1_58), .B(n_0_1_57), .ZN(n_0_1_56));
   XNOR2_X1 i_0_1_75 (.A(n_0_1_13), .B(n_0_1_21), .ZN(n_0_1_57));
   NOR2_X1 i_0_1_76 (.A1(n_0_1_68), .A2(n_0_1_59), .ZN(n_0_1_58));
   NOR2_X1 i_0_1_77 (.A1(EB[7]), .A2(EA[7]), .ZN(n_0_1_59));
   NAND2_X1 i_0_1_20 (.A1(n_0_1_69), .A2(n_0_1_66), .ZN(n_0_1_60));
   AOI21_X1 i_0_1_21 (.A(n_0_1_72), .B1(n_0_1_69), .B2(n_0_1_64), .ZN(n_0_1_62));
   NAND3_X1 i_0_1_64 (.A1(n_0_1_100), .A2(n_0_1_97), .A3(n_0_1_67), .ZN(n_0_1_64));
   AND2_X1 i_0_1_65 (.A1(n_0_1_112), .A2(A[31]), .ZN(n_0_103));
   OAI21_X1 i_0_1_125 (.A(n_0_1_112), .B1(n_0_1_28), .B2(clk), .ZN(n_0_104));
   AND2_X1 i_0_1_126 (.A1(n_0_1_112), .A2(B[31]), .ZN(n_0_105));
   AND2_X1 i_0_1_127 (.A1(n_0_1_112), .A2(A[0]), .ZN(n_0_106));
   AND2_X1 i_0_1_128 (.A1(n_0_1_112), .A2(A[1]), .ZN(n_0_107));
   AND2_X1 i_0_1_129 (.A1(n_0_1_112), .A2(A[2]), .ZN(n_0_108));
   AND2_X1 i_0_1_130 (.A1(n_0_1_112), .A2(A[3]), .ZN(n_0_109));
   AND2_X1 i_0_1_131 (.A1(n_0_1_112), .A2(A[4]), .ZN(n_0_110));
   AND2_X1 i_0_1_132 (.A1(n_0_1_112), .A2(A[5]), .ZN(n_0_111));
   AND2_X1 i_0_1_133 (.A1(n_0_1_112), .A2(A[6]), .ZN(n_0_112));
   AND2_X1 i_0_1_134 (.A1(n_0_1_112), .A2(A[7]), .ZN(n_0_113));
   AND2_X1 i_0_1_135 (.A1(n_0_1_112), .A2(A[8]), .ZN(n_0_114));
   AND2_X1 i_0_1_136 (.A1(n_0_1_112), .A2(A[9]), .ZN(n_0_115));
   AND2_X1 i_0_1_137 (.A1(n_0_1_112), .A2(A[10]), .ZN(n_0_116));
   AND2_X1 i_0_1_138 (.A1(n_0_1_112), .A2(A[11]), .ZN(n_0_117));
   AND2_X1 i_0_1_139 (.A1(n_0_1_112), .A2(A[12]), .ZN(n_0_118));
   AND2_X1 i_0_1_140 (.A1(n_0_1_112), .A2(A[13]), .ZN(n_0_119));
   AND2_X1 i_0_1_141 (.A1(n_0_1_112), .A2(A[14]), .ZN(n_0_120));
   AND2_X1 i_0_1_142 (.A1(n_0_1_112), .A2(A[15]), .ZN(n_0_121));
   AND2_X1 i_0_1_143 (.A1(n_0_1_112), .A2(A[16]), .ZN(n_0_122));
   AND2_X1 i_0_1_144 (.A1(n_0_1_112), .A2(A[17]), .ZN(n_0_123));
   AND2_X1 i_0_1_145 (.A1(n_0_1_112), .A2(A[18]), .ZN(n_0_124));
   AND2_X1 i_0_1_146 (.A1(n_0_1_112), .A2(A[19]), .ZN(n_0_125));
   AND2_X1 i_0_1_147 (.A1(n_0_1_112), .A2(A[20]), .ZN(n_0_126));
   AND2_X1 i_0_1_148 (.A1(n_0_1_112), .A2(A[21]), .ZN(n_0_127));
   AND2_X1 i_0_1_149 (.A1(n_0_1_112), .A2(A[22]), .ZN(n_0_128));
   AND2_X1 i_0_1_150 (.A1(n_0_1_112), .A2(A[23]), .ZN(n_0_129));
   AND2_X1 i_0_1_151 (.A1(n_0_1_112), .A2(A[24]), .ZN(n_0_130));
   AND2_X1 i_0_1_152 (.A1(n_0_1_112), .A2(A[25]), .ZN(n_0_131));
   AND2_X1 i_0_1_153 (.A1(n_0_1_112), .A2(A[26]), .ZN(n_0_132));
   AND2_X1 i_0_1_154 (.A1(n_0_1_112), .A2(A[27]), .ZN(n_0_133));
   AND2_X1 i_0_1_155 (.A1(n_0_1_112), .A2(A[28]), .ZN(n_0_134));
   AND2_X1 i_0_1_156 (.A1(n_0_1_112), .A2(A[29]), .ZN(n_0_135));
   AND2_X1 i_0_1_157 (.A1(n_0_1_112), .A2(A[30]), .ZN(n_0_136));
   AND2_X1 i_0_1_158 (.A1(n_0_1_112), .A2(B[0]), .ZN(n_0_137));
   AND2_X1 i_0_1_159 (.A1(n_0_1_112), .A2(B[1]), .ZN(n_0_138));
   AND2_X1 i_0_1_160 (.A1(n_0_1_112), .A2(B[2]), .ZN(n_0_139));
   AND2_X1 i_0_1_161 (.A1(n_0_1_112), .A2(B[3]), .ZN(n_0_140));
   AND2_X1 i_0_1_162 (.A1(n_0_1_112), .A2(B[4]), .ZN(n_0_141));
   AND2_X1 i_0_1_163 (.A1(n_0_1_112), .A2(B[5]), .ZN(n_0_142));
   AND2_X1 i_0_1_164 (.A1(n_0_1_112), .A2(B[6]), .ZN(n_0_143));
   AND2_X1 i_0_1_165 (.A1(n_0_1_112), .A2(B[7]), .ZN(n_0_144));
   AND2_X1 i_0_1_166 (.A1(n_0_1_112), .A2(B[8]), .ZN(n_0_145));
   AND2_X1 i_0_1_167 (.A1(n_0_1_112), .A2(B[9]), .ZN(n_0_146));
   AND2_X1 i_0_1_168 (.A1(n_0_1_112), .A2(B[10]), .ZN(n_0_147));
   AND2_X1 i_0_1_169 (.A1(n_0_1_112), .A2(B[11]), .ZN(n_0_148));
   AND2_X1 i_0_1_170 (.A1(n_0_1_112), .A2(B[12]), .ZN(n_0_149));
   AND2_X1 i_0_1_171 (.A1(n_0_1_112), .A2(B[13]), .ZN(n_0_150));
   AND2_X1 i_0_1_172 (.A1(n_0_1_112), .A2(B[14]), .ZN(n_0_151));
   AND2_X1 i_0_1_173 (.A1(n_0_1_112), .A2(B[15]), .ZN(n_0_152));
   AND2_X1 i_0_1_174 (.A1(n_0_1_112), .A2(B[16]), .ZN(n_0_153));
   AND2_X1 i_0_1_175 (.A1(n_0_1_112), .A2(B[17]), .ZN(n_0_154));
   AND2_X1 i_0_1_176 (.A1(n_0_1_112), .A2(B[18]), .ZN(n_0_155));
   AND2_X1 i_0_1_177 (.A1(n_0_1_112), .A2(B[19]), .ZN(n_0_156));
   AND2_X1 i_0_1_178 (.A1(n_0_1_112), .A2(B[20]), .ZN(n_0_157));
   AND2_X1 i_0_1_179 (.A1(n_0_1_112), .A2(B[21]), .ZN(n_0_158));
   AND2_X1 i_0_1_180 (.A1(n_0_1_112), .A2(B[22]), .ZN(n_0_159));
   AND2_X1 i_0_1_181 (.A1(n_0_1_112), .A2(B[23]), .ZN(n_0_160));
   AND2_X1 i_0_1_182 (.A1(n_0_1_112), .A2(B[24]), .ZN(n_0_161));
   AND2_X1 i_0_1_183 (.A1(n_0_1_112), .A2(B[25]), .ZN(n_0_162));
   AND2_X1 i_0_1_184 (.A1(n_0_1_112), .A2(B[26]), .ZN(n_0_163));
   AND2_X1 i_0_1_185 (.A1(n_0_1_112), .A2(B[27]), .ZN(n_0_164));
   AND2_X1 i_0_1_186 (.A1(n_0_1_112), .A2(B[28]), .ZN(n_0_165));
   AND2_X1 i_0_1_187 (.A1(n_0_1_112), .A2(B[29]), .ZN(n_0_166));
   AND2_X1 i_0_1_188 (.A1(n_0_1_112), .A2(B[30]), .ZN(n_0_167));
   OR2_X1 i_0_1_189 (.A1(clk), .A2(reset), .ZN(n_0_168));
   INV_X1 i_0_1_190 (.A(n_0_1_27), .ZN(n_0_1_105));
   INV_X1 i_0_1_191 (.A(n_0_1_26), .ZN(n_0_1_106));
   INV_X1 i_0_1_192 (.A(n_0_1_25), .ZN(n_0_1_107));
   INV_X1 i_0_1_193 (.A(n_0_1_24), .ZN(n_0_1_108));
   INV_X1 i_0_1_194 (.A(n_0_1_23), .ZN(n_0_1_109));
   INV_X1 i_0_1_195 (.A(n_0_1_22), .ZN(n_0_1_110));
   INV_X1 i_0_1_66 (.A(n_0_1_14), .ZN(n_0_1_111));
   INV_X1 i_0_1_78 (.A(reset), .ZN(n_0_1_112));
   INV_X1 i_0_1_198 (.A(enable), .ZN(n_0_1_28));
   INV_X1 i_0_1_79 (.A(n_0_24), .ZN(n_0_1_29));
   OAI21_X1 i_0_1_80 (.A(n_0_1_71), .B1(n_0_1_31), .B2(n_0_1_30), .ZN(n_0_71));
   OAI221_X1 i_0_1_81 (.A(n_0_1_69), .B1(n_0_1_100), .B2(n_0_1_81), .C1(n_0_1_97), 
      .C2(n_0_1_73), .ZN(n_0_1_30));
   INV_X1 i_0_1_82 (.A(n_0_1_61), .ZN(n_0_1_31));
   OAI211_X1 i_0_1_83 (.A(n_0_1_100), .B(n_0_1_97), .C1(n_0_1_65), .C2(n_0_1_63), 
      .ZN(n_0_1_61));
   NAND2_X1 i_0_1_84 (.A1(n_0_1_67), .A2(n_0_1_66), .ZN(n_0_1_63));
   AOI22_X1 i_0_1_85 (.A1(n_0_1_103), .A2(n_0_0), .B1(n_0_24), .B2(
      M_resultTruncated[0]), .ZN(n_0_1_65));
   OR4_X1 i_0_1_86 (.A1(n_0_1_101), .A2(n_0_1_98), .A3(n_0_1_92), .A4(n_0_1_95), 
      .ZN(n_0_1_66));
   OAI221_X1 i_0_1_87 (.A(n_0_1_68), .B1(EA[6]), .B2(n_0_1_98), .C1(EB[6]), 
      .C2(n_0_1_101), .ZN(n_0_1_67));
   AND2_X1 i_0_1_88 (.A1(EA[7]), .A2(EB[7]), .ZN(n_0_1_68));
   NOR2_X1 i_0_1_89 (.A1(reset), .A2(n_0_1_70), .ZN(n_0_1_69));
   OAI22_X1 i_0_1_90 (.A1(n_0_1_91), .A2(n_0_1_81), .B1(n_0_1_94), .B2(n_0_1_73), 
      .ZN(n_0_1_70));
   INV_X1 i_0_1_91 (.A(n_0_1_72), .ZN(n_0_1_71));
   NOR4_X1 i_0_1_92 (.A1(reset), .A2(n_0_1_73), .A3(n_0_1_81), .A4(n_0_1_89), 
      .ZN(n_0_1_72));
   NAND3_X1 i_0_1_93 (.A1(n_0_1_78), .A2(n_0_1_77), .A3(n_0_1_74), .ZN(n_0_1_73));
   AND4_X1 i_0_1_94 (.A1(n_0_1_80), .A2(n_0_1_79), .A3(n_0_1_76), .A4(n_0_1_75), 
      .ZN(n_0_1_74));
   NOR4_X1 i_0_1_95 (.A1(n_0_45), .A2(n_0_47), .A3(n_0_41), .A4(n_0_44), 
      .ZN(n_0_1_75));
   NOR4_X1 i_0_1_96 (.A1(n_0_37), .A2(n_0_40), .A3(n_0_34), .A4(n_0_35), 
      .ZN(n_0_1_76));
   NOR3_X1 i_0_1_97 (.A1(n_0_42), .A2(n_0_43), .A3(n_0_46), .ZN(n_0_1_77));
   NOR4_X1 i_0_1_98 (.A1(n_0_38), .A2(n_0_39), .A3(n_0_33), .A4(n_0_36), 
      .ZN(n_0_1_78));
   NOR4_X1 i_0_1_99 (.A1(n_0_25), .A2(n_0_26), .A3(n_0_27), .A4(n_0_28), 
      .ZN(n_0_1_79));
   NOR4_X1 i_0_1_100 (.A1(n_0_29), .A2(n_0_30), .A3(n_0_31), .A4(n_0_32), 
      .ZN(n_0_1_80));
   NAND3_X1 i_0_1_101 (.A1(n_0_1_86), .A2(n_0_1_85), .A3(n_0_1_82), .ZN(n_0_1_81));
   AND4_X1 i_0_1_102 (.A1(n_0_1_88), .A2(n_0_1_87), .A3(n_0_1_84), .A4(n_0_1_83), 
      .ZN(n_0_1_82));
   NOR4_X1 i_0_1_103 (.A1(n_0_68), .A2(n_0_70), .A3(n_0_64), .A4(n_0_67), 
      .ZN(n_0_1_83));
   NOR4_X1 i_0_1_104 (.A1(n_0_60), .A2(n_0_63), .A3(n_0_57), .A4(n_0_58), 
      .ZN(n_0_1_84));
   NOR3_X1 i_0_1_105 (.A1(n_0_65), .A2(n_0_66), .A3(n_0_69), .ZN(n_0_1_85));
   NOR4_X1 i_0_1_106 (.A1(n_0_61), .A2(n_0_62), .A3(n_0_56), .A4(n_0_59), 
      .ZN(n_0_1_86));
   NOR4_X1 i_0_1_107 (.A1(n_0_48), .A2(n_0_49), .A3(n_0_50), .A4(n_0_51), 
      .ZN(n_0_1_87));
   NOR4_X1 i_0_1_108 (.A1(n_0_52), .A2(n_0_53), .A3(n_0_54), .A4(n_0_55), 
      .ZN(n_0_1_88));
   INV_X1 i_0_1_109 (.A(n_0_1_90), .ZN(n_0_1_89));
   OAI22_X1 i_0_1_110 (.A1(n_0_1_100), .A2(n_0_1_94), .B1(n_0_1_97), .B2(
      n_0_1_91), .ZN(n_0_1_90));
   OR4_X1 i_0_1_111 (.A1(n_0_1_93), .A2(n_0_1_92), .A3(EB[5]), .A4(EB[4]), 
      .ZN(n_0_1_91));
   OR2_X1 i_0_1_112 (.A1(EB[7]), .A2(EB[6]), .ZN(n_0_1_92));
   OR4_X1 i_0_1_113 (.A1(EB[3]), .A2(EB[2]), .A3(EB[1]), .A4(EB[0]), .ZN(
      n_0_1_93));
   OR4_X1 i_0_1_114 (.A1(n_0_1_96), .A2(n_0_1_95), .A3(EA[5]), .A4(EA[4]), 
      .ZN(n_0_1_94));
   OR2_X1 i_0_1_115 (.A1(EA[7]), .A2(EA[6]), .ZN(n_0_1_95));
   OR4_X1 i_0_1_116 (.A1(EA[3]), .A2(EA[2]), .A3(EA[1]), .A4(EA[0]), .ZN(
      n_0_1_96));
   NAND3_X1 i_0_1_117 (.A1(EA[7]), .A2(n_0_1_98), .A3(EA[6]), .ZN(n_0_1_97));
   AND3_X1 i_0_1_118 (.A1(EA[2]), .A2(EA[1]), .A3(n_0_1_99), .ZN(n_0_1_98));
   AND4_X1 i_0_1_119 (.A1(EA[5]), .A2(EA[4]), .A3(EA[3]), .A4(EA[0]), .ZN(
      n_0_1_99));
   NAND3_X1 i_0_1_120 (.A1(EB[7]), .A2(n_0_1_101), .A3(EB[6]), .ZN(n_0_1_100));
   AND3_X1 i_0_1_121 (.A1(EB[2]), .A2(EB[1]), .A3(n_0_1_102), .ZN(n_0_1_101));
   AND4_X1 i_0_1_122 (.A1(EB[5]), .A2(EB[4]), .A3(EB[3]), .A4(EB[0]), .ZN(
      n_0_1_102));
   INV_X1 i_0_1_123 (.A(n_0_24), .ZN(n_0_1_103));
   AOI211_X1 i_0_1_124 (.A(reset), .B(n_0_1_104), .C1(B_reg), .C2(A_reg), 
      .ZN(n_0_102));
   NOR2_X1 i_0_1_196 (.A1(B_reg), .A2(A_reg), .ZN(n_0_1_104));
endmodule
