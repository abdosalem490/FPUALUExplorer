
// 	Thu Dec 22 19:44:55 2022
//	vlsi
//	192.168.126.129

module datapath__0_13 (Res_imm, p_0);

output [63:0] p_0;
input [63:0] Res_imm;
wire n_60;
wire n_0;
wire n_59;
wire n_58;
wire n_57;
wire n_1;
wire n_56;
wire n_55;
wire n_2;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_3;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_4;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire CLOCK_sgo__sro_n74;
wire n_11;
wire n_10;
wire n_5;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire sgo__n2;
wire sgo__sro_n8;
wire sgo__sro_n9;
wire sgo__sro_n10;
wire sgo__sro_n11;
wire CLOCK_sgo__sro_n71;
wire sgo__sro_n18;
wire sgo__sro_n19;
wire sgo__sro_n20;
wire sgo__sro_n21;
wire CLOCK_sgo__sro_n72;
wire sgo__sro_n28;
wire sgo__sro_n29;
wire sgo__sro_n30;
wire sgo__sro_n31;
wire CLOCK_sgo__sro_n73;
wire sgo__sro_n38;
wire sgo__sro_n39;
wire sgo__sro_n40;
wire sgo__sro_n41;
wire sgo__sro_n42;
wire sgo__sro_n52;
wire sgo__sro_n53;
wire sgo__sro_n54;
wire sgo__sro_n55;
wire sgo__sro_n56;


INV_X1 i_135 (.ZN (n_72), .A (Res_imm[62]));
INV_X1 i_134 (.ZN (n_71), .A (Res_imm[60]));
INV_X1 i_133 (.ZN (n_70), .A (Res_imm[55]));
INV_X1 i_132 (.ZN (n_69), .A (Res_imm[51]));
INV_X1 i_131 (.ZN (n_68), .A (Res_imm[42]));
INV_X1 i_130 (.ZN (n_67), .A (Res_imm[40]));
INV_X1 i_129 (.ZN (n_66), .A (Res_imm[36]));
INV_X1 i_128 (.ZN (n_65), .A (Res_imm[31]));
INV_X1 i_127 (.ZN (n_64), .A (Res_imm[26]));
INV_X1 i_126 (.ZN (n_63), .A (Res_imm[21]));
INV_X1 i_125 (.ZN (n_62), .A (Res_imm[13]));
INV_X1 i_124 (.ZN (n_61), .A (Res_imm[11]));
OR3_X4 i_123 (.ZN (n_60), .A1 (Res_imm[2]), .A2 (Res_imm[1]), .A3 (Res_imm[0]));
OR2_X4 i_122 (.ZN (n_59), .A1 (n_60), .A2 (Res_imm[3]));
OR2_X4 i_121 (.ZN (n_58), .A1 (n_59), .A2 (Res_imm[4]));
OR3_X4 i_120 (.ZN (n_57), .A1 (n_58), .A2 (Res_imm[5]), .A3 (Res_imm[6]));
OR2_X4 i_119 (.ZN (n_56), .A1 (n_57), .A2 (Res_imm[7]));
OR3_X4 i_118 (.ZN (n_55), .A1 (n_56), .A2 (Res_imm[8]), .A3 (Res_imm[9]));
NOR2_X4 i_117 (.ZN (n_54), .A1 (n_55), .A2 (Res_imm[10]));
NAND2_X4 i_116 (.ZN (n_53), .A1 (n_54), .A2 (n_61));
NOR2_X4 i_115 (.ZN (n_52), .A1 (n_53), .A2 (Res_imm[12]));
NAND2_X4 i_114 (.ZN (n_51), .A1 (n_52), .A2 (n_62));
OR3_X4 i_113 (.ZN (n_50), .A1 (n_51), .A2 (Res_imm[14]), .A3 (Res_imm[15]));
OR2_X4 i_112 (.ZN (n_49), .A1 (n_50), .A2 (Res_imm[16]));
OR2_X4 i_111 (.ZN (n_48), .A1 (n_49), .A2 (Res_imm[17]));
NOR2_X1 i_110 (.ZN (n_47), .A1 (n_48), .A2 (Res_imm[18]));
NOR3_X1 i_109 (.ZN (n_46), .A1 (n_48), .A2 (Res_imm[18]), .A3 (Res_imm[19]));
NAND2_X2 i_107 (.ZN (n_44), .A1 (sgo__sro_n52), .A2 (n_63));
OR2_X4 i_106 (.ZN (n_43), .A1 (n_44), .A2 (Res_imm[22]));
NOR2_X1 i_105 (.ZN (n_42), .A1 (n_43), .A2 (Res_imm[23]));
NOR3_X1 i_104 (.ZN (n_41), .A1 (n_43), .A2 (Res_imm[23]), .A3 (Res_imm[24]));
INV_X1 CLOCK_sgo__sro_c104 (.ZN (CLOCK_sgo__sro_n73), .A (Res_imm[49]));
NAND2_X2 i_102 (.ZN (n_39), .A1 (n_40), .A2 (n_64));
OR2_X4 i_101 (.ZN (n_38), .A1 (n_39), .A2 (Res_imm[27]));
NOR2_X1 i_100 (.ZN (n_37), .A1 (n_38), .A2 (Res_imm[28]));
NOR3_X1 i_99 (.ZN (n_36), .A1 (n_38), .A2 (Res_imm[28]), .A3 (Res_imm[29]));
NOR2_X4 CLOCK_sgo__sro_c107 (.ZN (n_16), .A1 (n_19), .A2 (CLOCK_sgo__sro_n71));
NAND2_X2 i_97 (.ZN (n_34), .A1 (n_35), .A2 (n_65));
OR2_X4 i_96 (.ZN (n_33), .A1 (n_34), .A2 (Res_imm[32]));
NOR2_X1 i_95 (.ZN (n_32), .A1 (n_33), .A2 (Res_imm[33]));
NOR3_X1 i_94 (.ZN (n_31), .A1 (n_33), .A2 (Res_imm[33]), .A3 (Res_imm[34]));
NAND2_X2 i_92 (.ZN (n_29), .A1 (n_30), .A2 (n_66));
OR2_X4 i_91 (.ZN (n_28), .A1 (n_29), .A2 (Res_imm[37]));
NOR2_X1 i_90 (.ZN (n_27), .A1 (n_28), .A2 (Res_imm[38]));
NOR3_X4 i_89 (.ZN (n_26), .A1 (n_28), .A2 (Res_imm[38]), .A3 (Res_imm[39]));
NAND2_X4 i_88 (.ZN (n_25), .A1 (n_26), .A2 (n_67));
NOR2_X4 i_87 (.ZN (n_24), .A1 (n_25), .A2 (Res_imm[41]));
NAND2_X4 i_86 (.ZN (n_23), .A1 (n_24), .A2 (n_68));
OR3_X4 i_85 (.ZN (n_22), .A1 (n_23), .A2 (Res_imm[43]), .A3 (Res_imm[44]));
OR2_X4 i_84 (.ZN (n_21), .A1 (n_22), .A2 (Res_imm[45]));
OR2_X4 i_83 (.ZN (n_20), .A1 (n_21), .A2 (Res_imm[46]));
OR2_X4 i_82 (.ZN (n_19), .A1 (n_20), .A2 (Res_imm[47]));
NOR2_X1 i_81 (.ZN (n_18), .A1 (n_19), .A2 (Res_imm[48]));
NOR3_X1 i_80 (.ZN (n_17), .A1 (n_19), .A2 (Res_imm[48]), .A3 (Res_imm[49]));
NAND2_X4 i_78 (.ZN (n_15), .A1 (n_16), .A2 (n_69));
NOR2_X1 i_77 (.ZN (n_14), .A1 (n_15), .A2 (Res_imm[52]));
NOR3_X1 i_76 (.ZN (n_13), .A1 (n_15), .A2 (Res_imm[52]), .A3 (Res_imm[53]));
NAND2_X2 i_74 (.ZN (n_11), .A1 (sgo__sro_n38), .A2 (n_70));
OR3_X4 i_73 (.ZN (n_10), .A1 (n_11), .A2 (Res_imm[56]), .A3 (Res_imm[57]));
NOR2_X1 i_72 (.ZN (n_9), .A1 (n_10), .A2 (Res_imm[58]));
NOR3_X4 i_71 (.ZN (n_8), .A1 (n_10), .A2 (Res_imm[58]), .A3 (Res_imm[59]));
NAND2_X2 i_70 (.ZN (n_7), .A1 (n_8), .A2 (n_71));
NOR2_X2 i_69 (.ZN (n_6), .A1 (n_7), .A2 (Res_imm[61]));
NAND2_X1 i_68 (.ZN (p_0[63]), .A1 (n_6), .A2 (n_72));
XNOR2_X1 i_67 (.ZN (p_0[62]), .A (Res_imm[62]), .B (n_6));
XOR2_X1 i_66 (.Z (p_0[61]), .A (Res_imm[61]), .B (n_7));
XNOR2_X1 i_65 (.ZN (p_0[60]), .A (Res_imm[60]), .B (n_8));
XNOR2_X1 i_64 (.ZN (p_0[59]), .A (Res_imm[59]), .B (n_9));
XOR2_X1 i_63 (.Z (p_0[58]), .A (Res_imm[58]), .B (n_10));
OAI21_X1 i_62 (.ZN (n_5), .A (Res_imm[57]), .B1 (n_11), .B2 (Res_imm[56]));
AND2_X1 i_61 (.ZN (p_0[57]), .A1 (n_10), .A2 (n_5));
XOR2_X1 i_60 (.Z (p_0[56]), .A (Res_imm[56]), .B (n_11));
XNOR2_X1 i_59 (.ZN (p_0[55]), .A (Res_imm[55]), .B (sgo__sro_n38));
XNOR2_X1 i_58 (.ZN (p_0[54]), .A (Res_imm[54]), .B (n_13));
XNOR2_X1 i_57 (.ZN (p_0[53]), .A (Res_imm[53]), .B (n_14));
XOR2_X1 i_56 (.Z (p_0[52]), .A (Res_imm[52]), .B (n_15));
XNOR2_X1 i_55 (.ZN (p_0[51]), .A (Res_imm[51]), .B (sgo__n2));
XNOR2_X1 i_54 (.ZN (p_0[50]), .A (Res_imm[50]), .B (n_17));
XNOR2_X1 i_53 (.ZN (p_0[49]), .A (Res_imm[49]), .B (n_18));
XOR2_X1 i_52 (.Z (p_0[48]), .A (Res_imm[48]), .B (n_19));
XOR2_X1 i_51 (.Z (p_0[47]), .A (Res_imm[47]), .B (n_20));
XOR2_X1 i_50 (.Z (p_0[46]), .A (Res_imm[46]), .B (n_21));
XOR2_X1 i_49 (.Z (p_0[45]), .A (Res_imm[45]), .B (n_22));
OAI21_X1 i_48 (.ZN (n_4), .A (Res_imm[44]), .B1 (n_23), .B2 (Res_imm[43]));
AND2_X1 i_47 (.ZN (p_0[44]), .A1 (n_22), .A2 (n_4));
XOR2_X1 i_46 (.Z (p_0[43]), .A (Res_imm[43]), .B (n_23));
XNOR2_X1 i_45 (.ZN (p_0[42]), .A (Res_imm[42]), .B (n_24));
XOR2_X1 i_44 (.Z (p_0[41]), .A (Res_imm[41]), .B (n_25));
XNOR2_X1 i_43 (.ZN (p_0[40]), .A (Res_imm[40]), .B (n_26));
XNOR2_X1 i_42 (.ZN (p_0[39]), .A (Res_imm[39]), .B (n_27));
XOR2_X1 i_41 (.Z (p_0[38]), .A (Res_imm[38]), .B (n_28));
XOR2_X1 i_40 (.Z (p_0[37]), .A (Res_imm[37]), .B (n_29));
XNOR2_X1 i_39 (.ZN (p_0[36]), .A (Res_imm[36]), .B (n_30));
XNOR2_X1 i_38 (.ZN (p_0[35]), .A (Res_imm[35]), .B (n_31));
XNOR2_X1 i_37 (.ZN (p_0[34]), .A (Res_imm[34]), .B (n_32));
XOR2_X1 i_36 (.Z (p_0[33]), .A (Res_imm[33]), .B (n_33));
XOR2_X1 i_35 (.Z (p_0[32]), .A (Res_imm[32]), .B (n_34));
XNOR2_X1 i_34 (.ZN (p_0[31]), .A (Res_imm[31]), .B (n_35));
XNOR2_X1 i_33 (.ZN (p_0[30]), .A (Res_imm[30]), .B (n_36));
XNOR2_X1 i_32 (.ZN (p_0[29]), .A (Res_imm[29]), .B (n_37));
XOR2_X1 i_31 (.Z (p_0[28]), .A (Res_imm[28]), .B (n_38));
XOR2_X1 i_30 (.Z (p_0[27]), .A (Res_imm[27]), .B (n_39));
XNOR2_X1 i_29 (.ZN (p_0[26]), .A (Res_imm[26]), .B (n_40));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (Res_imm[25]), .B (n_41));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (Res_imm[24]), .B (n_42));
XOR2_X1 i_26 (.Z (p_0[23]), .A (Res_imm[23]), .B (n_43));
XOR2_X1 i_25 (.Z (p_0[22]), .A (Res_imm[22]), .B (n_44));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (Res_imm[21]), .B (sgo__sro_n52));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (Res_imm[20]), .B (n_46));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (Res_imm[19]), .B (n_47));
XOR2_X1 i_21 (.Z (p_0[18]), .A (Res_imm[18]), .B (n_48));
XOR2_X1 i_20 (.Z (p_0[17]), .A (Res_imm[17]), .B (n_49));
XOR2_X1 i_19 (.Z (p_0[16]), .A (Res_imm[16]), .B (n_50));
OAI21_X1 i_18 (.ZN (n_3), .A (Res_imm[15]), .B1 (n_51), .B2 (Res_imm[14]));
AND2_X1 i_17 (.ZN (p_0[15]), .A1 (n_50), .A2 (n_3));
XOR2_X1 i_16 (.Z (p_0[14]), .A (Res_imm[14]), .B (n_51));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (Res_imm[13]), .B (n_52));
XOR2_X1 i_14 (.Z (p_0[12]), .A (Res_imm[12]), .B (n_53));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (Res_imm[11]), .B (n_54));
XOR2_X1 i_12 (.Z (p_0[10]), .A (Res_imm[10]), .B (n_55));
OAI21_X1 i_11 (.ZN (n_2), .A (Res_imm[9]), .B1 (n_56), .B2 (Res_imm[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_55), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (Res_imm[8]), .B (n_56));
XOR2_X1 i_8 (.Z (p_0[7]), .A (Res_imm[7]), .B (n_57));
OAI21_X1 i_7 (.ZN (n_1), .A (Res_imm[6]), .B1 (n_58), .B2 (Res_imm[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_57), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (Res_imm[5]), .B (n_58));
XOR2_X1 i_4 (.Z (p_0[4]), .A (Res_imm[4]), .B (n_59));
XOR2_X1 i_3 (.Z (p_0[3]), .A (Res_imm[3]), .B (n_60));
OAI21_X1 i_2 (.ZN (n_0), .A (Res_imm[2]), .B1 (Res_imm[1]), .B2 (Res_imm[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_60), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (Res_imm[1]), .B (Res_imm[0]));
CLKBUF_X1 sgo__L1_c1 (.Z (sgo__n2), .A (n_16));
INV_X1 CLOCK_sgo__sro_c103 (.ZN (CLOCK_sgo__sro_n74), .A (Res_imm[48]));
INV_X1 sgo__sro_c13 (.ZN (sgo__sro_n11), .A (Res_imm[23]));
INV_X1 sgo__sro_c14 (.ZN (sgo__sro_n10), .A (Res_imm[24]));
INV_X1 sgo__sro_c15 (.ZN (sgo__sro_n9), .A (Res_imm[25]));
NAND3_X1 sgo__sro_c16 (.ZN (sgo__sro_n8), .A1 (sgo__sro_n11), .A2 (sgo__sro_n9), .A3 (sgo__sro_n10));
NOR2_X4 sgo__sro_c17 (.ZN (n_40), .A1 (n_43), .A2 (sgo__sro_n8));
INV_X1 CLOCK_sgo__sro_c105 (.ZN (CLOCK_sgo__sro_n72), .A (Res_imm[50]));
NAND3_X1 CLOCK_sgo__sro_c106 (.ZN (CLOCK_sgo__sro_n71), .A1 (CLOCK_sgo__sro_n74), .A2 (CLOCK_sgo__sro_n72), .A3 (CLOCK_sgo__sro_n73));
INV_X1 sgo__sro_c30 (.ZN (sgo__sro_n21), .A (Res_imm[28]));
INV_X1 sgo__sro_c31 (.ZN (sgo__sro_n20), .A (Res_imm[29]));
INV_X1 sgo__sro_c32 (.ZN (sgo__sro_n19), .A (Res_imm[30]));
NAND3_X1 sgo__sro_c33 (.ZN (sgo__sro_n18), .A1 (sgo__sro_n21), .A2 (sgo__sro_n19), .A3 (sgo__sro_n20));
NOR2_X4 sgo__sro_c34 (.ZN (n_35), .A1 (n_38), .A2 (sgo__sro_n18));
INV_X1 sgo__sro_c47 (.ZN (sgo__sro_n31), .A (Res_imm[33]));
INV_X1 sgo__sro_c48 (.ZN (sgo__sro_n30), .A (Res_imm[34]));
INV_X1 sgo__sro_c49 (.ZN (sgo__sro_n29), .A (Res_imm[35]));
NAND3_X1 sgo__sro_c50 (.ZN (sgo__sro_n28), .A1 (sgo__sro_n31), .A2 (sgo__sro_n29), .A3 (sgo__sro_n30));
NOR2_X4 sgo__sro_c51 (.ZN (n_30), .A1 (n_33), .A2 (sgo__sro_n28));
INV_X1 sgo__sro_c64 (.ZN (sgo__sro_n42), .A (Res_imm[52]));
INV_X1 sgo__sro_c65 (.ZN (sgo__sro_n41), .A (Res_imm[53]));
INV_X1 sgo__sro_c66 (.ZN (sgo__sro_n40), .A (Res_imm[54]));
NAND3_X1 sgo__sro_c67 (.ZN (sgo__sro_n39), .A1 (sgo__sro_n42), .A2 (sgo__sro_n40), .A3 (sgo__sro_n41));
NOR2_X4 sgo__sro_c68 (.ZN (sgo__sro_n38), .A1 (n_15), .A2 (sgo__sro_n39));
INV_X1 sgo__sro_c81 (.ZN (sgo__sro_n56), .A (Res_imm[18]));
INV_X1 sgo__sro_c82 (.ZN (sgo__sro_n55), .A (Res_imm[19]));
INV_X1 sgo__sro_c83 (.ZN (sgo__sro_n54), .A (Res_imm[20]));
NAND3_X1 sgo__sro_c84 (.ZN (sgo__sro_n53), .A1 (sgo__sro_n56), .A2 (sgo__sro_n54), .A3 (sgo__sro_n55));
NOR2_X4 sgo__sro_c85 (.ZN (sgo__sro_n52), .A1 (n_48), .A2 (sgo__sro_n53));

endmodule //datapath__0_13

module datapath__0_6 (p_0, B);

output [31:0] p_0;
input [31:0] B;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (B[25]));
INV_X1 i_63 (.ZN (n_32), .A (B[21]));
INV_X1 i_62 (.ZN (n_31), .A (B[14]));
INV_X1 i_61 (.ZN (n_30), .A (B[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (B[2]), .A2 (B[1]), .A3 (B[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (B[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (B[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (B[5]), .A3 (B[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (B[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (B[8]), .A3 (B[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (B[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (B[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (B[12]), .A3 (B[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (B[15]), .A3 (B[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (B[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (B[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (B[18]), .A3 (B[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (B[18]), .A3 (B[19]), .A4 (B[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (B[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (B[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (B[23]), .A3 (B[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (B[26]), .A3 (B[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (B[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (B[28]), .A3 (B[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (B[28]), .A3 (B[29]), .A4 (B[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (B[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (B[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (B[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (B[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (B[27]), .B1 (n_9), .B2 (B[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (B[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (B[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (B[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (B[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (B[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (B[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (B[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (B[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (B[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (B[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (B[16]), .B1 (n_19), .B2 (B[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (B[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (B[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (B[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (B[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (B[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (B[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (B[9]), .B1 (n_25), .B2 (B[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (B[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (B[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (B[6]), .B1 (n_27), .B2 (B[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (B[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (B[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (B[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (B[2]), .B1 (B[1]), .B2 (B[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (B[1]), .B (B[0]));

endmodule //datapath__0_6

module datapath__0_4 (p_0, A);

output [31:0] p_0;
input [31:0] A;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (A[25]));
INV_X1 i_63 (.ZN (n_32), .A (A[21]));
INV_X1 i_62 (.ZN (n_31), .A (A[14]));
INV_X1 i_61 (.ZN (n_30), .A (A[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (A[2]), .A2 (A[1]), .A3 (A[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (A[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (A[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (A[5]), .A3 (A[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (A[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (A[8]), .A3 (A[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (A[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (A[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (A[12]), .A3 (A[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (A[15]), .A3 (A[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (A[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (A[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (A[18]), .A3 (A[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (A[18]), .A3 (A[19]), .A4 (A[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (A[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (A[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (A[23]), .A3 (A[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (A[26]), .A3 (A[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (A[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (A[28]), .A3 (A[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (A[28]), .A3 (A[29]), .A4 (A[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (A[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (A[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (A[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (A[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (A[27]), .B1 (n_9), .B2 (A[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (A[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (A[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (A[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (A[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (A[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (A[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (A[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (A[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (A[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (A[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (A[16]), .B1 (n_19), .B2 (A[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (A[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (A[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (A[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (A[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (A[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (A[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (A[9]), .B1 (n_25), .B2 (A[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (A[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (A[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (A[6]), .B1 (n_27), .B2 (A[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (A[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (A[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (A[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (A[2]), .B1 (A[1]), .B2 (A[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (A[1]), .B (A[0]));

endmodule //datapath__0_4

module datapath (p_0, accumulator, p_1);

output [31:0] p_1;
input [31:0] accumulator;
input [31:0] p_0;
wire n_0;
wire n_159;
wire n_1;
wire n_158;
wire n_157;
wire n_2;
wire n_162;
wire n_156;
wire n_3;
wire n_163;
wire n_168;
wire n_165;
wire n_154;
wire n_10;
wire n_9;
wire n_6;
wire n_7;
wire n_4;
wire n_151;
wire n_142;
wire n_11;
wire n_5;
wire n_152;
wire n_146;
wire n_8;
wire n_149;
wire n_147;
wire n_153;
wire n_144;
wire n_140;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_12;
wire n_137;
wire n_128;
wire n_19;
wire n_13;
wire n_138;
wire n_132;
wire n_16;
wire n_135;
wire n_133;
wire n_139;
wire n_130;
wire n_126;
wire n_26;
wire n_25;
wire n_22;
wire n_23;
wire n_20;
wire n_123;
wire n_114;
wire n_27;
wire n_21;
wire n_124;
wire n_118;
wire n_24;
wire n_121;
wire n_119;
wire n_125;
wire n_116;
wire n_112;
wire n_34;
wire n_33;
wire n_30;
wire n_31;
wire n_28;
wire n_109;
wire n_100;
wire n_35;
wire n_29;
wire n_110;
wire n_104;
wire n_32;
wire n_107;
wire n_105;
wire n_111;
wire n_102;
wire n_98;
wire n_42;
wire n_41;
wire n_38;
wire n_39;
wire n_36;
wire n_87;
wire n_77;
wire n_43;
wire n_37;
wire n_86;
wire n_89;
wire n_79;
wire n_40;
wire n_88;
wire n_84;
wire n_81;
wire n_91;
wire n_52;
wire n_51;
wire n_49;
wire n_48;
wire n_45;
wire n_44;
wire n_72;
wire n_95;
wire n_68;
wire n_53;
wire n_46;
wire n_47;
wire n_94;
wire n_69;
wire n_50;
wire n_96;
wire n_73;
wire n_74;
wire n_76;
wire n_83;
wire n_97;
wire n_66;
wire n_65;
wire n_63;
wire n_59;
wire n_64;
wire n_58;
wire n_55;
wire n_54;
wire n_60;
wire n_62;
wire n_56;
wire n_57;
wire n_61;
wire n_170;
wire n_167;
wire n_164;
wire n_70;
wire n_67;
wire n_75;
wire n_82;
wire n_169;
wire n_166;
wire n_71;
wire n_93;
wire n_92;
wire n_78;
wire n_90;
wire n_85;
wire n_80;
wire n_99;
wire n_103;
wire n_106;
wire n_101;
wire n_108;
wire n_113;
wire n_117;
wire n_120;
wire n_115;
wire n_122;
wire n_127;
wire n_131;
wire n_134;
wire n_129;
wire n_136;
wire n_141;
wire n_145;
wire n_148;
wire n_143;
wire n_150;
wire n_155;
wire n_161;
wire n_160;


INV_X1 i_202 (.ZN (n_170), .A (p_0[29]));
INV_X1 i_201 (.ZN (n_169), .A (p_0[27]));
INV_X1 i_200 (.ZN (n_168), .A (p_0[3]));
INV_X1 i_199 (.ZN (n_167), .A (accumulator[29]));
INV_X1 i_198 (.ZN (n_166), .A (accumulator[27]));
INV_X1 i_197 (.ZN (n_165), .A (accumulator[3]));
NOR2_X1 i_196 (.ZN (n_164), .A1 (p_0[28]), .A2 (accumulator[28]));
NAND2_X1 i_195 (.ZN (n_163), .A1 (n_168), .A2 (n_165));
NAND2_X1 i_194 (.ZN (n_162), .A1 (p_0[2]), .A2 (accumulator[2]));
INV_X1 i_193 (.ZN (n_161), .A (n_162));
NOR2_X1 i_192 (.ZN (n_160), .A1 (p_0[1]), .A2 (accumulator[1]));
NAND2_X1 i_191 (.ZN (n_159), .A1 (p_0[0]), .A2 (accumulator[0]));
NAND2_X1 i_190 (.ZN (n_158), .A1 (p_0[1]), .A2 (accumulator[1]));
AOI21_X1 i_189 (.ZN (n_157), .A (n_160), .B1 (n_159), .B2 (n_158));
OAI22_X1 i_188 (.ZN (n_156), .A1 (p_0[2]), .A2 (accumulator[2]), .B1 (n_161), .B2 (n_157));
OAI21_X1 i_187 (.ZN (n_155), .A (n_156), .B1 (n_168), .B2 (n_165));
NAND2_X1 i_186 (.ZN (n_154), .A1 (n_163), .A2 (n_155));
NOR2_X1 i_185 (.ZN (n_153), .A1 (p_0[7]), .A2 (accumulator[7]));
NOR2_X1 i_184 (.ZN (n_152), .A1 (p_0[5]), .A2 (accumulator[5]));
NOR2_X1 i_183 (.ZN (n_151), .A1 (p_0[6]), .A2 (accumulator[6]));
OR3_X1 i_182 (.ZN (n_150), .A1 (n_153), .A2 (n_151), .A3 (n_152));
NOR2_X1 i_181 (.ZN (n_149), .A1 (p_0[4]), .A2 (accumulator[4]));
NOR3_X1 i_180 (.ZN (n_148), .A1 (n_150), .A2 (n_149), .A3 (n_154));
NAND2_X1 i_179 (.ZN (n_147), .A1 (p_0[4]), .A2 (accumulator[4]));
NAND2_X1 i_178 (.ZN (n_146), .A1 (p_0[5]), .A2 (accumulator[5]));
AOI21_X1 i_177 (.ZN (n_145), .A (n_150), .B1 (n_147), .B2 (n_146));
AND2_X1 i_176 (.ZN (n_144), .A1 (p_0[7]), .A2 (accumulator[7]));
NAND2_X1 i_175 (.ZN (n_143), .A1 (p_0[6]), .A2 (accumulator[6]));
INV_X1 i_174 (.ZN (n_142), .A (n_143));
NOR2_X1 i_173 (.ZN (n_141), .A1 (n_153), .A2 (n_143));
NOR4_X1 i_172 (.ZN (n_140), .A1 (n_144), .A2 (n_141), .A3 (n_145), .A4 (n_148));
NOR2_X1 i_171 (.ZN (n_139), .A1 (p_0[11]), .A2 (accumulator[11]));
NOR2_X1 i_170 (.ZN (n_138), .A1 (p_0[9]), .A2 (accumulator[9]));
NOR2_X1 i_169 (.ZN (n_137), .A1 (p_0[10]), .A2 (accumulator[10]));
OR3_X1 i_168 (.ZN (n_136), .A1 (n_139), .A2 (n_137), .A3 (n_138));
NOR2_X1 i_167 (.ZN (n_135), .A1 (p_0[8]), .A2 (accumulator[8]));
NOR3_X1 i_166 (.ZN (n_134), .A1 (n_136), .A2 (n_135), .A3 (n_140));
NAND2_X1 i_165 (.ZN (n_133), .A1 (p_0[8]), .A2 (accumulator[8]));
NAND2_X1 i_164 (.ZN (n_132), .A1 (p_0[9]), .A2 (accumulator[9]));
AOI21_X1 i_163 (.ZN (n_131), .A (n_136), .B1 (n_133), .B2 (n_132));
AND2_X1 i_162 (.ZN (n_130), .A1 (p_0[11]), .A2 (accumulator[11]));
NAND2_X1 i_161 (.ZN (n_129), .A1 (p_0[10]), .A2 (accumulator[10]));
INV_X1 i_160 (.ZN (n_128), .A (n_129));
NOR2_X1 i_159 (.ZN (n_127), .A1 (n_139), .A2 (n_129));
NOR4_X1 i_158 (.ZN (n_126), .A1 (n_130), .A2 (n_127), .A3 (n_131), .A4 (n_134));
NOR2_X1 i_157 (.ZN (n_125), .A1 (p_0[15]), .A2 (accumulator[15]));
NOR2_X1 i_156 (.ZN (n_124), .A1 (p_0[13]), .A2 (accumulator[13]));
NOR2_X1 i_155 (.ZN (n_123), .A1 (p_0[14]), .A2 (accumulator[14]));
OR3_X1 i_154 (.ZN (n_122), .A1 (n_125), .A2 (n_123), .A3 (n_124));
NOR2_X1 i_153 (.ZN (n_121), .A1 (p_0[12]), .A2 (accumulator[12]));
NOR3_X1 i_152 (.ZN (n_120), .A1 (n_122), .A2 (n_121), .A3 (n_126));
NAND2_X1 i_151 (.ZN (n_119), .A1 (p_0[12]), .A2 (accumulator[12]));
NAND2_X1 i_150 (.ZN (n_118), .A1 (p_0[13]), .A2 (accumulator[13]));
AOI21_X1 i_149 (.ZN (n_117), .A (n_122), .B1 (n_119), .B2 (n_118));
AND2_X1 i_148 (.ZN (n_116), .A1 (p_0[15]), .A2 (accumulator[15]));
NAND2_X1 i_147 (.ZN (n_115), .A1 (p_0[14]), .A2 (accumulator[14]));
INV_X1 i_146 (.ZN (n_114), .A (n_115));
NOR2_X1 i_145 (.ZN (n_113), .A1 (n_125), .A2 (n_115));
NOR4_X1 i_144 (.ZN (n_112), .A1 (n_116), .A2 (n_113), .A3 (n_117), .A4 (n_120));
NOR2_X1 i_143 (.ZN (n_111), .A1 (p_0[19]), .A2 (accumulator[19]));
NOR2_X1 i_142 (.ZN (n_110), .A1 (p_0[17]), .A2 (accumulator[17]));
NOR2_X1 i_141 (.ZN (n_109), .A1 (p_0[18]), .A2 (accumulator[18]));
OR3_X1 i_140 (.ZN (n_108), .A1 (n_111), .A2 (n_109), .A3 (n_110));
NOR2_X1 i_139 (.ZN (n_107), .A1 (p_0[16]), .A2 (accumulator[16]));
NOR3_X1 i_138 (.ZN (n_106), .A1 (n_108), .A2 (n_107), .A3 (n_112));
NAND2_X1 i_137 (.ZN (n_105), .A1 (p_0[16]), .A2 (accumulator[16]));
NAND2_X1 i_136 (.ZN (n_104), .A1 (p_0[17]), .A2 (accumulator[17]));
AOI21_X1 i_135 (.ZN (n_103), .A (n_108), .B1 (n_105), .B2 (n_104));
AND2_X1 i_134 (.ZN (n_102), .A1 (p_0[19]), .A2 (accumulator[19]));
NAND2_X1 i_133 (.ZN (n_101), .A1 (p_0[18]), .A2 (accumulator[18]));
INV_X1 i_132 (.ZN (n_100), .A (n_101));
NOR2_X1 i_131 (.ZN (n_99), .A1 (n_111), .A2 (n_101));
NOR4_X1 i_130 (.ZN (n_98), .A1 (n_102), .A2 (n_99), .A3 (n_103), .A4 (n_106));
NOR2_X1 i_129 (.ZN (n_97), .A1 (p_0[27]), .A2 (accumulator[27]));
NOR2_X1 i_128 (.ZN (n_96), .A1 (p_0[25]), .A2 (accumulator[25]));
NOR2_X1 i_127 (.ZN (n_95), .A1 (p_0[26]), .A2 (accumulator[26]));
NOR2_X1 i_126 (.ZN (n_94), .A1 (n_96), .A2 (n_95));
NOR3_X1 i_125 (.ZN (n_93), .A1 (n_97), .A2 (n_95), .A3 (n_96));
OAI21_X1 i_124 (.ZN (n_92), .A (n_93), .B1 (p_0[24]), .B2 (accumulator[24]));
NOR2_X1 i_123 (.ZN (n_91), .A1 (p_0[23]), .A2 (accumulator[23]));
INV_X1 i_122 (.ZN (n_90), .A (n_91));
NOR2_X1 i_121 (.ZN (n_89), .A1 (p_0[21]), .A2 (accumulator[21]));
INV_X1 i_120 (.ZN (n_88), .A (n_89));
NOR2_X1 i_119 (.ZN (n_87), .A1 (p_0[22]), .A2 (accumulator[22]));
INV_X1 i_118 (.ZN (n_86), .A (n_87));
NAND3_X1 i_117 (.ZN (n_85), .A1 (n_90), .A2 (n_86), .A3 (n_88));
NOR2_X1 i_116 (.ZN (n_84), .A1 (p_0[20]), .A2 (accumulator[20]));
OR2_X1 i_115 (.ZN (n_83), .A1 (n_85), .A2 (n_84));
NOR3_X1 i_114 (.ZN (n_82), .A1 (n_92), .A2 (n_83), .A3 (n_98));
NAND2_X1 i_113 (.ZN (n_81), .A1 (p_0[20]), .A2 (accumulator[20]));
NAND2_X1 i_112 (.ZN (n_80), .A1 (p_0[21]), .A2 (accumulator[21]));
INV_X1 i_111 (.ZN (n_79), .A (n_80));
AOI21_X1 i_110 (.ZN (n_78), .A (n_85), .B1 (n_81), .B2 (n_80));
AND2_X1 i_109 (.ZN (n_77), .A1 (p_0[22]), .A2 (accumulator[22]));
AOI221_X1 i_108 (.ZN (n_76), .A (n_78), .B1 (p_0[23]), .B2 (accumulator[23]), .C1 (n_90), .C2 (n_77));
NOR2_X1 i_107 (.ZN (n_75), .A1 (n_92), .A2 (n_76));
NAND2_X1 i_106 (.ZN (n_74), .A1 (p_0[24]), .A2 (accumulator[24]));
INV_X1 i_105 (.ZN (n_73), .A (n_74));
AND2_X1 i_104 (.ZN (n_72), .A1 (p_0[25]), .A2 (accumulator[25]));
OAI21_X1 i_103 (.ZN (n_71), .A (n_93), .B1 (n_73), .B2 (n_72));
INV_X1 i_102 (.ZN (n_70), .A (n_71));
NAND2_X1 i_101 (.ZN (n_69), .A1 (p_0[26]), .A2 (accumulator[26]));
INV_X1 i_100 (.ZN (n_68), .A (n_69));
OAI22_X1 i_99 (.ZN (n_67), .A1 (n_169), .A2 (n_166), .B1 (n_97), .B2 (n_69));
NOR4_X1 i_98 (.ZN (n_66), .A1 (n_70), .A2 (n_67), .A3 (n_75), .A4 (n_82));
AOI21_X1 i_97 (.ZN (n_65), .A (n_164), .B1 (p_0[28]), .B2 (accumulator[28]));
AOI21_X1 i_96 (.ZN (n_64), .A (n_164), .B1 (n_66), .B2 (n_65));
INV_X1 i_95 (.ZN (n_63), .A (n_64));
NAND2_X1 i_94 (.ZN (n_62), .A1 (p_0[30]), .A2 (accumulator[30]));
INV_X1 i_93 (.ZN (n_61), .A (n_62));
NAND2_X1 i_92 (.ZN (n_60), .A1 (n_170), .A2 (n_167));
OAI21_X1 i_91 (.ZN (n_59), .A (n_60), .B1 (n_170), .B2 (n_167));
INV_X1 i_90 (.ZN (n_58), .A (n_59));
NAND3_X1 i_89 (.ZN (n_57), .A1 (n_62), .A2 (n_58), .A3 (n_63));
OAI221_X1 i_88 (.ZN (n_56), .A (n_57), .B1 (p_0[30]), .B2 (accumulator[30]), .C1 (n_61), .C2 (n_60));
XNOR2_X1 i_87 (.ZN (p_1[31]), .A (p_0[31]), .B (n_56));
OAI21_X1 i_86 (.ZN (n_55), .A (n_62), .B1 (p_0[30]), .B2 (accumulator[30]));
AOI22_X1 i_85 (.ZN (n_54), .A1 (p_0[29]), .A2 (accumulator[29]), .B1 (n_64), .B2 (n_60));
XOR2_X1 i_84 (.Z (p_1[30]), .A (n_55), .B (n_54));
AOI22_X1 i_83 (.ZN (p_1[29]), .A1 (n_63), .A2 (n_59), .B1 (n_64), .B2 (n_58));
XNOR2_X1 i_82 (.ZN (p_1[28]), .A (n_66), .B (n_65));
AOI21_X1 i_81 (.ZN (n_53), .A (n_97), .B1 (p_0[27]), .B2 (accumulator[27]));
OAI21_X1 i_80 (.ZN (n_52), .A (n_76), .B1 (n_98), .B2 (n_83));
OAI21_X1 i_79 (.ZN (n_51), .A (n_74), .B1 (p_0[24]), .B2 (accumulator[24]));
OAI22_X1 i_78 (.ZN (n_50), .A1 (p_0[24]), .A2 (accumulator[24]), .B1 (n_73), .B2 (n_52));
INV_X1 i_77 (.ZN (n_49), .A (n_50));
NOR2_X1 i_76 (.ZN (n_48), .A1 (n_96), .A2 (n_72));
NAND3_X1 i_75 (.ZN (n_47), .A1 (n_69), .A2 (n_48), .A3 (n_50));
OAI21_X1 i_74 (.ZN (n_46), .A (n_47), .B1 (n_94), .B2 (n_68));
XNOR2_X1 i_73 (.ZN (p_1[27]), .A (n_53), .B (n_46));
NOR2_X1 i_72 (.ZN (n_45), .A1 (n_95), .A2 (n_68));
OAI22_X1 i_71 (.ZN (n_44), .A1 (p_0[25]), .A2 (accumulator[25]), .B1 (n_72), .B2 (n_49));
XNOR2_X1 i_70 (.ZN (p_1[26]), .A (n_45), .B (n_44));
XOR2_X1 i_69 (.Z (p_1[25]), .A (n_49), .B (n_48));
XNOR2_X1 i_68 (.ZN (p_1[24]), .A (n_52), .B (n_51));
AOI21_X1 i_67 (.ZN (n_43), .A (n_91), .B1 (p_0[23]), .B2 (accumulator[23]));
OAI21_X1 i_66 (.ZN (n_42), .A (n_81), .B1 (p_0[20]), .B2 (accumulator[20]));
AOI21_X1 i_65 (.ZN (n_41), .A (n_84), .B1 (n_98), .B2 (n_81));
OAI21_X1 i_64 (.ZN (n_40), .A (n_88), .B1 (n_79), .B2 (n_41));
INV_X1 i_63 (.ZN (n_39), .A (n_40));
NOR2_X1 i_62 (.ZN (n_38), .A1 (n_89), .A2 (n_79));
OAI21_X1 i_61 (.ZN (n_37), .A (n_86), .B1 (n_77), .B2 (n_39));
XNOR2_X1 i_60 (.ZN (p_1[23]), .A (n_43), .B (n_37));
NOR2_X1 i_59 (.ZN (n_36), .A1 (n_87), .A2 (n_77));
XOR2_X1 i_58 (.Z (p_1[22]), .A (n_39), .B (n_36));
XOR2_X1 i_57 (.Z (p_1[21]), .A (n_41), .B (n_38));
XOR2_X1 i_56 (.Z (p_1[20]), .A (n_98), .B (n_42));
NOR2_X1 i_55 (.ZN (n_35), .A1 (n_111), .A2 (n_102));
OAI21_X1 i_54 (.ZN (n_34), .A (n_105), .B1 (p_0[16]), .B2 (accumulator[16]));
AOI21_X1 i_53 (.ZN (n_33), .A (n_107), .B1 (n_112), .B2 (n_105));
INV_X1 i_52 (.ZN (n_32), .A (n_33));
AOI21_X1 i_51 (.ZN (n_31), .A (n_110), .B1 (n_104), .B2 (n_32));
AOI21_X1 i_50 (.ZN (n_30), .A (n_110), .B1 (p_0[17]), .B2 (accumulator[17]));
OAI22_X1 i_49 (.ZN (n_29), .A1 (p_0[18]), .A2 (accumulator[18]), .B1 (n_100), .B2 (n_31));
XNOR2_X1 i_48 (.ZN (p_1[19]), .A (n_35), .B (n_29));
NOR2_X1 i_47 (.ZN (n_28), .A1 (n_109), .A2 (n_100));
XOR2_X1 i_46 (.Z (p_1[18]), .A (n_31), .B (n_28));
XOR2_X1 i_45 (.Z (p_1[17]), .A (n_33), .B (n_30));
XOR2_X1 i_44 (.Z (p_1[16]), .A (n_112), .B (n_34));
NOR2_X1 i_43 (.ZN (n_27), .A1 (n_125), .A2 (n_116));
OAI21_X1 i_42 (.ZN (n_26), .A (n_119), .B1 (p_0[12]), .B2 (accumulator[12]));
AOI21_X1 i_41 (.ZN (n_25), .A (n_121), .B1 (n_126), .B2 (n_119));
INV_X1 i_40 (.ZN (n_24), .A (n_25));
AOI21_X1 i_39 (.ZN (n_23), .A (n_124), .B1 (n_118), .B2 (n_24));
AOI21_X1 i_38 (.ZN (n_22), .A (n_124), .B1 (p_0[13]), .B2 (accumulator[13]));
OAI22_X1 i_37 (.ZN (n_21), .A1 (p_0[14]), .A2 (accumulator[14]), .B1 (n_114), .B2 (n_23));
XNOR2_X1 i_36 (.ZN (p_1[15]), .A (n_27), .B (n_21));
NOR2_X1 i_35 (.ZN (n_20), .A1 (n_123), .A2 (n_114));
XOR2_X1 i_34 (.Z (p_1[14]), .A (n_23), .B (n_20));
XOR2_X1 i_33 (.Z (p_1[13]), .A (n_25), .B (n_22));
XOR2_X1 i_32 (.Z (p_1[12]), .A (n_126), .B (n_26));
NOR2_X1 i_31 (.ZN (n_19), .A1 (n_139), .A2 (n_130));
AOI21_X1 i_30 (.ZN (n_18), .A (n_135), .B1 (p_0[8]), .B2 (accumulator[8]));
AOI21_X1 i_29 (.ZN (n_17), .A (n_135), .B1 (n_140), .B2 (n_133));
INV_X1 i_28 (.ZN (n_16), .A (n_17));
AOI21_X1 i_27 (.ZN (n_15), .A (n_138), .B1 (n_132), .B2 (n_16));
AOI21_X1 i_26 (.ZN (n_14), .A (n_138), .B1 (p_0[9]), .B2 (accumulator[9]));
OAI22_X1 i_25 (.ZN (n_13), .A1 (p_0[10]), .A2 (accumulator[10]), .B1 (n_128), .B2 (n_15));
XNOR2_X1 i_24 (.ZN (p_1[11]), .A (n_19), .B (n_13));
NOR2_X1 i_23 (.ZN (n_12), .A1 (n_137), .A2 (n_128));
XOR2_X1 i_22 (.Z (p_1[10]), .A (n_15), .B (n_12));
XOR2_X1 i_21 (.Z (p_1[9]), .A (n_17), .B (n_14));
XNOR2_X1 i_20 (.ZN (p_1[8]), .A (n_140), .B (n_18));
NOR2_X1 i_19 (.ZN (n_11), .A1 (n_153), .A2 (n_144));
OAI21_X1 i_18 (.ZN (n_10), .A (n_147), .B1 (p_0[4]), .B2 (accumulator[4]));
AOI21_X1 i_17 (.ZN (n_9), .A (n_149), .B1 (n_154), .B2 (n_147));
INV_X1 i_16 (.ZN (n_8), .A (n_9));
AOI21_X1 i_15 (.ZN (n_7), .A (n_152), .B1 (n_146), .B2 (n_8));
AOI21_X1 i_14 (.ZN (n_6), .A (n_152), .B1 (p_0[5]), .B2 (accumulator[5]));
OAI22_X1 i_13 (.ZN (n_5), .A1 (p_0[6]), .A2 (accumulator[6]), .B1 (n_142), .B2 (n_7));
XNOR2_X1 i_12 (.ZN (p_1[7]), .A (n_11), .B (n_5));
NOR2_X1 i_11 (.ZN (n_4), .A1 (n_151), .A2 (n_142));
XOR2_X1 i_10 (.Z (p_1[6]), .A (n_7), .B (n_4));
XOR2_X1 i_9 (.Z (p_1[5]), .A (n_9), .B (n_6));
XOR2_X1 i_8 (.Z (p_1[4]), .A (n_154), .B (n_10));
OAI21_X1 i_7 (.ZN (n_3), .A (n_163), .B1 (n_168), .B2 (n_165));
XOR2_X1 i_6 (.Z (p_1[3]), .A (n_156), .B (n_3));
OAI21_X1 i_5 (.ZN (n_2), .A (n_162), .B1 (p_0[2]), .B2 (accumulator[2]));
XNOR2_X1 i_4 (.ZN (p_1[2]), .A (n_157), .B (n_2));
OAI21_X1 i_3 (.ZN (n_1), .A (n_158), .B1 (p_0[1]), .B2 (accumulator[1]));
XOR2_X1 i_2 (.Z (p_1[1]), .A (n_159), .B (n_1));
OAI21_X1 i_1 (.ZN (n_0), .A (n_159), .B1 (p_0[0]), .B2 (accumulator[0]));
INV_X1 i_0 (.ZN (p_1[0]), .A (n_0));

endmodule //datapath

module sequentialMultiplier (Res, OVF, A, B, clk, reset, enable);

output OVF;
output [63:0] Res;
input [31:0] A;
input [31:0] B;
input clk;
input enable;
input reset;
wire drc_ipo_n18;
wire CTS_n_tid1_102;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire \isNeg[1] ;
wire \isNeg[0] ;
wire \accumulator[30] ;
wire \accumulator[29] ;
wire \accumulator[28] ;
wire \accumulator[27] ;
wire \accumulator[26] ;
wire \accumulator[25] ;
wire \accumulator[24] ;
wire \accumulator[23] ;
wire \accumulator[22] ;
wire \accumulator[21] ;
wire \accumulator[20] ;
wire \accumulator[19] ;
wire \accumulator[18] ;
wire \accumulator[17] ;
wire \accumulator[16] ;
wire \accumulator[15] ;
wire \accumulator[14] ;
wire \accumulator[13] ;
wire \accumulator[12] ;
wire \accumulator[11] ;
wire \accumulator[10] ;
wire \accumulator[9] ;
wire \accumulator[8] ;
wire \accumulator[7] ;
wire \accumulator[6] ;
wire \accumulator[5] ;
wire \accumulator[4] ;
wire \accumulator[3] ;
wire \accumulator[2] ;
wire \accumulator[1] ;
wire \accumulator[0] ;
wire \multiplier[31] ;
wire \multiplier[30] ;
wire \multiplier[29] ;
wire \multiplier[28] ;
wire \multiplier[27] ;
wire \multiplier[26] ;
wire \multiplier[25] ;
wire \multiplier[24] ;
wire \multiplier[23] ;
wire \multiplier[22] ;
wire \multiplier[21] ;
wire \multiplier[20] ;
wire \multiplier[19] ;
wire \multiplier[18] ;
wire \multiplier[17] ;
wire \multiplier[16] ;
wire \multiplier[15] ;
wire \multiplier[14] ;
wire \multiplier[13] ;
wire \multiplier[12] ;
wire \multiplier[11] ;
wire \multiplier[10] ;
wire \multiplier[9] ;
wire \multiplier[8] ;
wire \multiplier[7] ;
wire \multiplier[6] ;
wire \multiplier[5] ;
wire \multiplier[4] ;
wire \multiplier[3] ;
wire \multiplier[2] ;
wire \multiplier[1] ;
wire \multiplier[0] ;
wire \multiplicand[31] ;
wire \multiplicand[30] ;
wire \multiplicand[29] ;
wire \multiplicand[28] ;
wire \multiplicand[27] ;
wire \multiplicand[26] ;
wire \multiplicand[25] ;
wire \multiplicand[24] ;
wire \multiplicand[23] ;
wire \multiplicand[22] ;
wire \multiplicand[21] ;
wire \multiplicand[20] ;
wire \multiplicand[19] ;
wire \multiplicand[18] ;
wire \multiplicand[17] ;
wire \multiplicand[16] ;
wire \multiplicand[15] ;
wire \multiplicand[14] ;
wire \multiplicand[13] ;
wire \multiplicand[12] ;
wire \multiplicand[11] ;
wire \multiplicand[10] ;
wire \multiplicand[9] ;
wire \multiplicand[8] ;
wire \multiplicand[7] ;
wire \multiplicand[6] ;
wire \multiplicand[5] ;
wire \multiplicand[4] ;
wire \multiplicand[3] ;
wire \multiplicand[2] ;
wire \multiplicand[1] ;
wire ready;
wire n_0_159;
wire \counter[4] ;
wire \counter[3] ;
wire \counter[2] ;
wire \counter[1] ;
wire \counter[0] ;
wire CTS_n_tid1_103;
wire n_0_0_0;
wire n_0_0_1;
wire n_0_0_2;
wire n_0_0_3;
wire n_0_0_4;
wire n_0_0_5;
wire n_0_0_6;
wire n_0_0_7;
wire n_0_0_8;
wire n_0_0_9;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_0_12;
wire n_0_0_13;
wire n_0_0_14;
wire n_0_0_15;
wire n_0_0_16;
wire n_0_0_17;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_0_20;
wire n_0_0_21;
wire n_0_0_22;
wire \counter_in[4] ;
wire \counter_in[3] ;
wire \counter_in[2] ;
wire \counter_in[1] ;
wire \counter_in[0] ;
wire n_0_0_23;
wire n_0_0_24;
wire n_0_0_25;
wire n_0_0_26;
wire n_0_0_27;
wire n_0_160;
wire n_0_161;
wire n_0_0_28;
wire n_0_0_29;
wire n_0_0_30;
wire \multiplicand_in[31] ;
wire \multiplicand_in[30] ;
wire \multiplicand_in[29] ;
wire \multiplicand_in[28] ;
wire \multiplicand_in[27] ;
wire \multiplicand_in[26] ;
wire \multiplicand_in[25] ;
wire \multiplicand_in[24] ;
wire \multiplicand_in[23] ;
wire \multiplicand_in[22] ;
wire \multiplicand_in[21] ;
wire \multiplicand_in[20] ;
wire \multiplicand_in[19] ;
wire \multiplicand_in[18] ;
wire \multiplicand_in[17] ;
wire \multiplicand_in[16] ;
wire \multiplicand_in[15] ;
wire \multiplicand_in[14] ;
wire \multiplicand_in[13] ;
wire \multiplicand_in[12] ;
wire \multiplicand_in[11] ;
wire \multiplicand_in[10] ;
wire \multiplicand_in[9] ;
wire \multiplicand_in[8] ;
wire \multiplicand_in[7] ;
wire \multiplicand_in[6] ;
wire \multiplicand_in[5] ;
wire \multiplicand_in[4] ;
wire \multiplicand_in[3] ;
wire \multiplicand_in[2] ;
wire \multiplicand_in[1] ;
wire \multiplicand_in[0] ;
wire n_0_0_32;
wire n_0_0_33;
wire n_0_0_34;
wire n_0_0_35;
wire n_0_0_36;
wire n_0_0_37;
wire n_0_0_38;
wire n_0_0_39;
wire n_0_0_40;
wire n_0_0_41;
wire n_0_0_42;
wire n_0_0_43;
wire n_0_0_44;
wire n_0_0_45;
wire n_0_0_46;
wire n_0_0_47;
wire n_0_0_48;
wire n_0_0_49;
wire n_0_0_50;
wire n_0_0_51;
wire n_0_0_52;
wire n_0_0_53;
wire n_0_0_54;
wire n_0_0_55;
wire n_0_0_56;
wire n_0_0_57;
wire n_0_0_58;
wire n_0_0_59;
wire n_0_0_60;
wire n_0_0_61;
wire n_0_0_62;
wire n_0_0_63;
wire n_0_0_64;
wire n_0_162;
wire n_0_163;
wire n_0_0_65;
wire n_0_164;
wire n_0_0_66;
wire n_0_165;
wire n_0_0_67;
wire n_0_166;
wire n_0_0_68;
wire n_0_167;
wire n_0_0_69;
wire n_0_168;
wire n_0_0_70;
wire n_0_169;
wire n_0_0_71;
wire n_0_170;
wire n_0_0_72;
wire n_0_171;
wire n_0_0_73;
wire n_0_172;
wire n_0_0_74;
wire n_0_173;
wire n_0_0_75;
wire n_0_174;
wire n_0_0_76;
wire n_0_175;
wire n_0_0_77;
wire n_0_176;
wire n_0_0_78;
wire n_0_177;
wire n_0_0_79;
wire n_0_178;
wire n_0_0_80;
wire n_0_179;
wire n_0_0_81;
wire n_0_180;
wire n_0_0_82;
wire n_0_181;
wire n_0_0_83;
wire n_0_182;
wire n_0_0_84;
wire n_0_183;
wire n_0_0_85;
wire n_0_184;
wire n_0_0_86;
wire n_0_185;
wire n_0_0_87;
wire n_0_186;
wire n_0_0_88;
wire n_0_187;
wire n_0_0_89;
wire n_0_188;
wire n_0_0_90;
wire n_0_189;
wire n_0_0_91;
wire n_0_190;
wire n_0_0_92;
wire n_0_191;
wire n_0_0_93;
wire n_0_192;
wire n_0_0_94;
wire n_0_0_95;
wire n_0_0_96;
wire n_0_193;
wire n_0_0_98;
wire n_0_194;
wire n_0_195;
wire n_0_196;
wire n_0_197;
wire n_0_198;
wire n_0_199;
wire n_0_200;
wire n_0_201;
wire n_0_202;
wire n_0_203;
wire n_0_204;
wire n_0_205;
wire n_0_206;
wire n_0_207;
wire n_0_208;
wire n_0_209;
wire n_0_210;
wire n_0_211;
wire n_0_212;
wire n_0_213;
wire n_0_214;
wire n_0_215;
wire n_0_216;
wire n_0_217;
wire n_0_218;
wire n_0_219;
wire n_0_220;
wire n_0_221;
wire n_0_222;
wire n_0_223;
wire n_0_224;
wire n_0_225;
wire n_0_226;
wire n_0_227;
wire n_0_228;
wire n_0_229;
wire n_0_230;
wire n_0_231;
wire n_0_232;
wire n_0_233;
wire n_0_234;
wire n_0_235;
wire n_0_236;
wire n_0_237;
wire n_0_238;
wire n_0_239;
wire n_0_240;
wire n_0_241;
wire n_0_242;
wire n_0_243;
wire n_0_244;
wire n_0_245;
wire n_0_246;
wire n_0_247;
wire n_0_248;
wire n_0_249;
wire n_0_250;
wire n_0_251;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_255;
wire n_0_256;
wire n_0_257;
wire \isNeg_in[1] ;
wire \isNeg_in[0] ;
wire n_0_258;
wire n_0_0_101;
wire n_0_0_102;
wire n_0_0_103;
wire n_0_0_104;
wire n_0_0_105;
wire n_0_0_106;
wire n_0_0_107;
wire n_0_0_31;
wire n_0_0_97;
wire n_0_0_99;
wire n_0_0_100;
wire n_0_0_108;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire hfn_ipo_n14;
wire hfn_ipo_n15;
wire hfn_ipo_n16;
wire hfn_ipo_n13;
wire sgo__n20;
wire sgo__n21;
wire CTS_n_tid1_28;
wire CTS_n_tid0_29;
wire CTS_n_tid0_30;
wire CTS_n_tid1_31;
wire CTS_n_tid1_32;
wire CTS_n_tid0_92;


NOR2_X1 i_0_0_310 (.ZN (n_0_0_108), .A1 (ready), .A2 (reset));
NAND2_X1 i_0_0_309 (.ZN (n_0_0_100), .A1 (ready), .A2 (enable));
NOR2_X1 i_0_0_308 (.ZN (n_0_0_99), .A1 (reset), .A2 (n_0_0_100));
INV_X1 i_0_0_307 (.ZN (n_0_0_97), .A (n_0_0_99));
AOI22_X1 i_0_0_306 (.ZN (n_0_0_31), .A1 (\multiplicand[1] ), .A2 (hfn_ipo_n16), .B1 (B[0]), .B2 (n_0_0_99));
INV_X1 i_0_0_304 (.ZN (\multiplicand_in[0] ), .A (n_0_0_31));
INV_X1 i_0_0_303 (.ZN (n_0_0_107), .A (n_0_0_100));
INV_X1 i_0_0_302 (.ZN (n_0_0_106), .A (hfn_ipo_n16));
INV_X1 i_0_0_301 (.ZN (n_0_0_105), .A (ready));
INV_X1 i_0_0_299 (.ZN (n_0_0_104), .A (A[31]));
INV_X1 i_0_0_305 (.ZN (n_0_0_103), .A (A[0]));
INV_X1 i_0_0_298 (.ZN (n_0_0_102), .A (B[31]));
INV_X1 i_0_0_265 (.ZN (n_0_0_101), .A (\isNeg[0] ));
OR2_X1 i_0_0_231 (.ZN (n_0_258), .A1 (reset), .A2 (n_0_0_107));
NOR2_X1 i_0_0_300 (.ZN (\isNeg_in[1] ), .A1 (n_0_0_104), .A2 (reset));
NOR2_X1 i_0_0_230 (.ZN (\isNeg_in[0] ), .A1 (n_0_0_102), .A2 (reset));
OR3_X1 i_0_0_229 (.ZN (n_0_257), .A1 (n_0_0_105), .A2 (reset), .A3 (enable));
AND2_X1 i_0_0_297 (.ZN (n_0_256), .A1 (\multiplier[31] ), .A2 (sgo__n21));
AND2_X1 i_0_0_296 (.ZN (n_0_255), .A1 (\multiplier[30] ), .A2 (sgo__n21));
AND2_X1 i_0_0_295 (.ZN (n_0_254), .A1 (\multiplier[29] ), .A2 (sgo__n21));
AND2_X1 i_0_0_294 (.ZN (n_0_253), .A1 (\multiplier[28] ), .A2 (sgo__n20));
AND2_X1 i_0_0_293 (.ZN (n_0_252), .A1 (\multiplier[27] ), .A2 (sgo__n20));
AND2_X1 i_0_0_292 (.ZN (n_0_251), .A1 (\multiplier[26] ), .A2 (sgo__n21));
AND2_X1 i_0_0_291 (.ZN (n_0_250), .A1 (\multiplier[25] ), .A2 (sgo__n20));
AND2_X1 i_0_0_290 (.ZN (n_0_249), .A1 (\multiplier[24] ), .A2 (sgo__n20));
AND2_X1 i_0_0_289 (.ZN (n_0_248), .A1 (\multiplier[23] ), .A2 (sgo__n20));
AND2_X1 i_0_0_288 (.ZN (n_0_247), .A1 (\multiplier[22] ), .A2 (sgo__n20));
AND2_X1 i_0_0_287 (.ZN (n_0_246), .A1 (\multiplier[21] ), .A2 (sgo__n20));
AND2_X1 i_0_0_286 (.ZN (n_0_245), .A1 (\multiplier[20] ), .A2 (sgo__n20));
AND2_X1 i_0_0_285 (.ZN (n_0_244), .A1 (\multiplier[19] ), .A2 (sgo__n20));
AND2_X1 i_0_0_284 (.ZN (n_0_243), .A1 (\multiplier[18] ), .A2 (sgo__n20));
AND2_X1 i_0_0_283 (.ZN (n_0_242), .A1 (\multiplier[17] ), .A2 (sgo__n20));
AND2_X1 i_0_0_282 (.ZN (n_0_241), .A1 (\multiplier[16] ), .A2 (sgo__n20));
AND2_X1 i_0_0_281 (.ZN (n_0_240), .A1 (\multiplier[15] ), .A2 (sgo__n20));
AND2_X1 i_0_0_280 (.ZN (n_0_239), .A1 (\multiplier[14] ), .A2 (sgo__n20));
AND2_X1 i_0_0_279 (.ZN (n_0_238), .A1 (\multiplier[13] ), .A2 (sgo__n20));
AND2_X1 i_0_0_278 (.ZN (n_0_237), .A1 (\multiplier[12] ), .A2 (sgo__n20));
AND2_X1 i_0_0_277 (.ZN (n_0_236), .A1 (\multiplier[11] ), .A2 (sgo__n21));
AND2_X1 i_0_0_276 (.ZN (n_0_235), .A1 (\multiplier[10] ), .A2 (sgo__n21));
AND2_X1 i_0_0_275 (.ZN (n_0_234), .A1 (\multiplier[9] ), .A2 (sgo__n21));
AND2_X1 i_0_0_274 (.ZN (n_0_233), .A1 (\multiplier[8] ), .A2 (sgo__n21));
AND2_X1 i_0_0_273 (.ZN (n_0_232), .A1 (\multiplier[7] ), .A2 (sgo__n21));
AND2_X1 i_0_0_272 (.ZN (n_0_231), .A1 (\multiplier[6] ), .A2 (sgo__n21));
AND2_X1 i_0_0_271 (.ZN (n_0_230), .A1 (\multiplier[5] ), .A2 (sgo__n21));
AND2_X1 i_0_0_270 (.ZN (n_0_229), .A1 (\multiplier[4] ), .A2 (sgo__n21));
AND2_X1 i_0_0_269 (.ZN (n_0_228), .A1 (\multiplier[3] ), .A2 (sgo__n21));
AND2_X1 i_0_0_268 (.ZN (n_0_227), .A1 (\multiplier[2] ), .A2 (sgo__n21));
AND2_X1 i_0_0_267 (.ZN (n_0_226), .A1 (\multiplier[1] ), .A2 (sgo__n21));
AND2_X1 i_0_0_266 (.ZN (n_0_225), .A1 (\multiplier[0] ), .A2 (sgo__n21));
AND2_X1 i_0_0_264 (.ZN (n_0_224), .A1 (n_0_33), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_263 (.ZN (n_0_223), .A1 (n_0_32), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_262 (.ZN (n_0_222), .A1 (n_0_31), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_261 (.ZN (n_0_221), .A1 (n_0_30), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_260 (.ZN (n_0_220), .A1 (n_0_29), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_259 (.ZN (n_0_219), .A1 (n_0_28), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_258 (.ZN (n_0_218), .A1 (n_0_27), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_257 (.ZN (n_0_217), .A1 (n_0_26), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_256 (.ZN (n_0_216), .A1 (n_0_25), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_255 (.ZN (n_0_215), .A1 (n_0_24), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_254 (.ZN (n_0_214), .A1 (n_0_23), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_253 (.ZN (n_0_213), .A1 (n_0_22), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_252 (.ZN (n_0_212), .A1 (n_0_21), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_251 (.ZN (n_0_211), .A1 (n_0_20), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_250 (.ZN (n_0_210), .A1 (n_0_19), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_249 (.ZN (n_0_209), .A1 (n_0_18), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_248 (.ZN (n_0_208), .A1 (n_0_17), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_247 (.ZN (n_0_207), .A1 (n_0_16), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_246 (.ZN (n_0_206), .A1 (n_0_15), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_245 (.ZN (n_0_205), .A1 (n_0_14), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_244 (.ZN (n_0_204), .A1 (n_0_13), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_243 (.ZN (n_0_203), .A1 (n_0_12), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_242 (.ZN (n_0_202), .A1 (n_0_11), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_241 (.ZN (n_0_201), .A1 (n_0_10), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_240 (.ZN (n_0_200), .A1 (n_0_9), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_239 (.ZN (n_0_199), .A1 (n_0_8), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_238 (.ZN (n_0_198), .A1 (n_0_7), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_237 (.ZN (n_0_197), .A1 (n_0_6), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_236 (.ZN (n_0_196), .A1 (n_0_5), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_235 (.ZN (n_0_195), .A1 (n_0_4), .A2 (hfn_ipo_n15));
AND2_X1 i_0_0_234 (.ZN (n_0_194), .A1 (n_0_3), .A2 (hfn_ipo_n15));
NOR2_X1 i_0_0_233 (.ZN (n_0_0_98), .A1 (n_0_0_100), .A2 (n_0_64));
NOR3_X1 i_0_0_232 (.ZN (n_0_193), .A1 (reset), .A2 (n_0_0_98), .A3 (n_0_0_104));
NOR2_X4 i_0_0_198 (.ZN (n_0_0_96), .A1 (n_0_0_104), .A2 (n_0_0_97));
AOI21_X4 i_0_0_197 (.ZN (n_0_0_95), .A (reset), .B1 (A[31]), .B2 (n_0_0_107));
AOI22_X1 i_0_0_228 (.ZN (n_0_0_94), .A1 (n_0_63), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[30]));
INV_X1 i_0_0_227 (.ZN (n_0_192), .A (n_0_0_94));
AOI22_X1 i_0_0_226 (.ZN (n_0_0_93), .A1 (n_0_62), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[29]));
INV_X1 i_0_0_225 (.ZN (n_0_191), .A (n_0_0_93));
AOI22_X1 i_0_0_224 (.ZN (n_0_0_92), .A1 (n_0_61), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[28]));
INV_X1 i_0_0_223 (.ZN (n_0_190), .A (n_0_0_92));
AOI22_X1 i_0_0_222 (.ZN (n_0_0_91), .A1 (n_0_60), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[27]));
INV_X1 i_0_0_221 (.ZN (n_0_189), .A (n_0_0_91));
AOI22_X1 i_0_0_220 (.ZN (n_0_0_90), .A1 (n_0_59), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[26]));
INV_X1 i_0_0_219 (.ZN (n_0_188), .A (n_0_0_90));
AOI22_X1 i_0_0_218 (.ZN (n_0_0_89), .A1 (n_0_58), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[25]));
INV_X1 i_0_0_217 (.ZN (n_0_187), .A (n_0_0_89));
AOI22_X1 i_0_0_216 (.ZN (n_0_0_88), .A1 (n_0_57), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[24]));
INV_X1 i_0_0_215 (.ZN (n_0_186), .A (n_0_0_88));
AOI22_X1 i_0_0_214 (.ZN (n_0_0_87), .A1 (n_0_56), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[23]));
INV_X1 i_0_0_213 (.ZN (n_0_185), .A (n_0_0_87));
AOI22_X1 i_0_0_212 (.ZN (n_0_0_86), .A1 (n_0_55), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[22]));
INV_X1 i_0_0_211 (.ZN (n_0_184), .A (n_0_0_86));
AOI22_X1 i_0_0_210 (.ZN (n_0_0_85), .A1 (n_0_54), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[21]));
INV_X1 i_0_0_209 (.ZN (n_0_183), .A (n_0_0_85));
AOI22_X1 i_0_0_208 (.ZN (n_0_0_84), .A1 (n_0_53), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[20]));
INV_X1 i_0_0_207 (.ZN (n_0_182), .A (n_0_0_84));
AOI22_X1 i_0_0_206 (.ZN (n_0_0_83), .A1 (n_0_52), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[19]));
INV_X1 i_0_0_205 (.ZN (n_0_181), .A (n_0_0_83));
AOI22_X1 i_0_0_204 (.ZN (n_0_0_82), .A1 (n_0_51), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[18]));
INV_X1 i_0_0_203 (.ZN (n_0_180), .A (n_0_0_82));
AOI22_X1 i_0_0_202 (.ZN (n_0_0_81), .A1 (n_0_50), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[17]));
INV_X1 i_0_0_201 (.ZN (n_0_179), .A (n_0_0_81));
AOI22_X1 i_0_0_200 (.ZN (n_0_0_80), .A1 (n_0_49), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[16]));
INV_X1 i_0_0_199 (.ZN (n_0_178), .A (n_0_0_80));
AOI22_X1 i_0_0_167 (.ZN (n_0_0_79), .A1 (n_0_48), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[15]));
INV_X1 i_0_0_164 (.ZN (n_0_177), .A (n_0_0_79));
AOI22_X1 i_0_0_196 (.ZN (n_0_0_78), .A1 (n_0_47), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[14]));
INV_X1 i_0_0_195 (.ZN (n_0_176), .A (n_0_0_78));
AOI22_X1 i_0_0_194 (.ZN (n_0_0_77), .A1 (n_0_46), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[13]));
INV_X1 i_0_0_193 (.ZN (n_0_175), .A (n_0_0_77));
AOI22_X1 i_0_0_192 (.ZN (n_0_0_76), .A1 (n_0_45), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[12]));
INV_X1 i_0_0_191 (.ZN (n_0_174), .A (n_0_0_76));
AOI22_X1 i_0_0_190 (.ZN (n_0_0_75), .A1 (n_0_44), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[11]));
INV_X1 i_0_0_189 (.ZN (n_0_173), .A (n_0_0_75));
AOI22_X1 i_0_0_188 (.ZN (n_0_0_74), .A1 (n_0_43), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[10]));
INV_X1 i_0_0_187 (.ZN (n_0_172), .A (n_0_0_74));
AOI22_X1 i_0_0_186 (.ZN (n_0_0_73), .A1 (n_0_42), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[9]));
INV_X1 i_0_0_185 (.ZN (n_0_171), .A (n_0_0_73));
AOI22_X1 i_0_0_184 (.ZN (n_0_0_72), .A1 (n_0_41), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[8]));
INV_X1 i_0_0_183 (.ZN (n_0_170), .A (n_0_0_72));
AOI22_X1 i_0_0_182 (.ZN (n_0_0_71), .A1 (n_0_40), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[7]));
INV_X1 i_0_0_181 (.ZN (n_0_169), .A (n_0_0_71));
AOI22_X1 i_0_0_180 (.ZN (n_0_0_70), .A1 (n_0_39), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[6]));
INV_X1 i_0_0_179 (.ZN (n_0_168), .A (n_0_0_70));
AOI22_X1 i_0_0_178 (.ZN (n_0_0_69), .A1 (n_0_38), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[5]));
INV_X1 i_0_0_177 (.ZN (n_0_167), .A (n_0_0_69));
AOI22_X1 i_0_0_176 (.ZN (n_0_0_68), .A1 (n_0_37), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[4]));
INV_X1 i_0_0_175 (.ZN (n_0_166), .A (n_0_0_68));
AOI22_X1 i_0_0_174 (.ZN (n_0_0_67), .A1 (n_0_36), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[3]));
INV_X1 i_0_0_173 (.ZN (n_0_165), .A (n_0_0_67));
AOI22_X1 i_0_0_172 (.ZN (n_0_0_66), .A1 (n_0_35), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[2]));
INV_X1 i_0_0_171 (.ZN (n_0_164), .A (n_0_0_66));
AOI22_X1 i_0_0_170 (.ZN (n_0_0_65), .A1 (n_0_34), .A2 (n_0_0_96), .B1 (n_0_0_95), .B2 (A[1]));
INV_X1 i_0_0_169 (.ZN (n_0_163), .A (n_0_0_65));
NOR2_X1 i_0_0_168 (.ZN (n_0_162), .A1 (n_0_0_103), .A2 (reset));
NOR2_X4 i_0_0_105 (.ZN (n_0_0_64), .A1 (n_0_0_102), .A2 (n_0_0_97));
AOI22_X1 i_0_0_166 (.ZN (n_0_0_63), .A1 (n_0_2), .A2 (hfn_ipo_n16), .B1 (n_0_0_64), .B2 (n_0_95));
INV_X1 i_0_0_165 (.ZN (\multiplicand_in[31] ), .A (n_0_0_63));
NOR2_X4 i_0_0_104 (.ZN (n_0_0_62), .A1 (n_0_0_97), .A2 (B[31]));
AOI222_X1 i_0_0_163 (.ZN (n_0_0_61), .A1 (\multiplicand[31] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_94), .C1 (n_0_0_62), .C2 (B[30]));
INV_X1 i_0_0_162 (.ZN (\multiplicand_in[30] ), .A (n_0_0_61));
AOI222_X1 i_0_0_161 (.ZN (n_0_0_60), .A1 (\multiplicand[30] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_93), .C1 (n_0_0_62), .C2 (B[29]));
INV_X1 i_0_0_160 (.ZN (\multiplicand_in[29] ), .A (n_0_0_60));
AOI222_X1 i_0_0_159 (.ZN (n_0_0_59), .A1 (\multiplicand[29] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_92), .C1 (n_0_0_62), .C2 (B[28]));
INV_X1 i_0_0_158 (.ZN (\multiplicand_in[28] ), .A (n_0_0_59));
AOI222_X1 i_0_0_157 (.ZN (n_0_0_58), .A1 (\multiplicand[28] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_91), .C1 (n_0_0_62), .C2 (B[27]));
INV_X1 i_0_0_156 (.ZN (\multiplicand_in[27] ), .A (n_0_0_58));
AOI222_X1 i_0_0_155 (.ZN (n_0_0_57), .A1 (\multiplicand[27] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_90), .C1 (n_0_0_62), .C2 (B[26]));
INV_X1 i_0_0_154 (.ZN (\multiplicand_in[26] ), .A (n_0_0_57));
AOI222_X1 i_0_0_153 (.ZN (n_0_0_56), .A1 (\multiplicand[26] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_89), .C1 (n_0_0_62), .C2 (B[25]));
INV_X1 i_0_0_152 (.ZN (\multiplicand_in[25] ), .A (n_0_0_56));
AOI222_X1 i_0_0_151 (.ZN (n_0_0_55), .A1 (\multiplicand[25] ), .A2 (hfn_ipo_n15), .B1 (n_0_0_64)
    , .B2 (n_0_88), .C1 (n_0_0_62), .C2 (B[24]));
INV_X1 i_0_0_150 (.ZN (\multiplicand_in[24] ), .A (n_0_0_55));
AOI222_X1 i_0_0_149 (.ZN (n_0_0_54), .A1 (\multiplicand[24] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_87), .C1 (n_0_0_62), .C2 (B[23]));
INV_X1 i_0_0_148 (.ZN (\multiplicand_in[23] ), .A (n_0_0_54));
AOI222_X1 i_0_0_147 (.ZN (n_0_0_53), .A1 (\multiplicand[23] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_86), .C1 (n_0_0_62), .C2 (B[22]));
INV_X1 i_0_0_146 (.ZN (\multiplicand_in[22] ), .A (n_0_0_53));
AOI222_X1 i_0_0_145 (.ZN (n_0_0_52), .A1 (\multiplicand[22] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_85), .C1 (n_0_0_62), .C2 (B[21]));
INV_X1 i_0_0_144 (.ZN (\multiplicand_in[21] ), .A (n_0_0_52));
AOI222_X1 i_0_0_143 (.ZN (n_0_0_51), .A1 (\multiplicand[21] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_84), .C1 (n_0_0_62), .C2 (B[20]));
INV_X1 i_0_0_142 (.ZN (\multiplicand_in[20] ), .A (n_0_0_51));
AOI222_X1 i_0_0_141 (.ZN (n_0_0_50), .A1 (\multiplicand[20] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_83), .C1 (n_0_0_62), .C2 (B[19]));
INV_X1 i_0_0_140 (.ZN (\multiplicand_in[19] ), .A (n_0_0_50));
AOI222_X1 i_0_0_139 (.ZN (n_0_0_49), .A1 (\multiplicand[19] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_82), .C1 (n_0_0_62), .C2 (B[18]));
INV_X1 i_0_0_138 (.ZN (\multiplicand_in[18] ), .A (n_0_0_49));
AOI222_X1 i_0_0_137 (.ZN (n_0_0_48), .A1 (\multiplicand[18] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_81), .C1 (n_0_0_62), .C2 (B[17]));
INV_X1 i_0_0_136 (.ZN (\multiplicand_in[17] ), .A (n_0_0_48));
AOI222_X1 i_0_0_135 (.ZN (n_0_0_47), .A1 (\multiplicand[17] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_80), .C1 (n_0_0_62), .C2 (B[16]));
INV_X1 i_0_0_134 (.ZN (\multiplicand_in[16] ), .A (n_0_0_47));
AOI222_X1 i_0_0_133 (.ZN (n_0_0_46), .A1 (\multiplicand[16] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_79), .C1 (n_0_0_62), .C2 (B[15]));
INV_X1 i_0_0_132 (.ZN (\multiplicand_in[15] ), .A (n_0_0_46));
AOI222_X1 i_0_0_131 (.ZN (n_0_0_45), .A1 (\multiplicand[15] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_78), .C1 (n_0_0_62), .C2 (B[14]));
INV_X1 i_0_0_130 (.ZN (\multiplicand_in[14] ), .A (n_0_0_45));
AOI222_X1 i_0_0_129 (.ZN (n_0_0_44), .A1 (\multiplicand[14] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_77), .C1 (n_0_0_62), .C2 (B[13]));
INV_X1 i_0_0_128 (.ZN (\multiplicand_in[13] ), .A (n_0_0_44));
AOI222_X1 i_0_0_127 (.ZN (n_0_0_43), .A1 (\multiplicand[13] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_76), .C1 (n_0_0_62), .C2 (B[12]));
INV_X1 i_0_0_126 (.ZN (\multiplicand_in[12] ), .A (n_0_0_43));
AOI222_X1 i_0_0_125 (.ZN (n_0_0_42), .A1 (\multiplicand[12] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_75), .C1 (n_0_0_62), .C2 (B[11]));
INV_X1 i_0_0_124 (.ZN (\multiplicand_in[11] ), .A (n_0_0_42));
AOI222_X1 i_0_0_123 (.ZN (n_0_0_41), .A1 (\multiplicand[11] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_74), .C1 (n_0_0_62), .C2 (B[10]));
INV_X1 i_0_0_122 (.ZN (\multiplicand_in[10] ), .A (n_0_0_41));
AOI222_X1 i_0_0_121 (.ZN (n_0_0_40), .A1 (\multiplicand[10] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_73), .C1 (n_0_0_62), .C2 (B[9]));
INV_X1 i_0_0_120 (.ZN (\multiplicand_in[9] ), .A (n_0_0_40));
AOI222_X1 i_0_0_119 (.ZN (n_0_0_39), .A1 (\multiplicand[9] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_72), .C1 (n_0_0_62), .C2 (B[8]));
INV_X1 i_0_0_118 (.ZN (\multiplicand_in[8] ), .A (n_0_0_39));
AOI222_X1 i_0_0_117 (.ZN (n_0_0_38), .A1 (\multiplicand[8] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_71), .C1 (n_0_0_62), .C2 (B[7]));
INV_X1 i_0_0_116 (.ZN (\multiplicand_in[7] ), .A (n_0_0_38));
AOI222_X1 i_0_0_115 (.ZN (n_0_0_37), .A1 (\multiplicand[7] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_70), .C1 (n_0_0_62), .C2 (B[6]));
INV_X1 i_0_0_114 (.ZN (\multiplicand_in[6] ), .A (n_0_0_37));
AOI222_X1 i_0_0_113 (.ZN (n_0_0_36), .A1 (\multiplicand[6] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_69), .C1 (n_0_0_62), .C2 (B[5]));
INV_X1 i_0_0_112 (.ZN (\multiplicand_in[5] ), .A (n_0_0_36));
AOI222_X1 i_0_0_111 (.ZN (n_0_0_35), .A1 (\multiplicand[5] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_68), .C1 (n_0_0_62), .C2 (B[4]));
INV_X1 i_0_0_110 (.ZN (\multiplicand_in[4] ), .A (n_0_0_35));
AOI222_X1 i_0_0_109 (.ZN (n_0_0_34), .A1 (\multiplicand[4] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_67), .C1 (n_0_0_62), .C2 (B[3]));
INV_X1 i_0_0_108 (.ZN (\multiplicand_in[3] ), .A (n_0_0_34));
AOI222_X1 i_0_0_107 (.ZN (n_0_0_33), .A1 (\multiplicand[3] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_66), .C1 (n_0_0_62), .C2 (B[2]));
INV_X1 i_0_0_106 (.ZN (\multiplicand_in[2] ), .A (n_0_0_33));
AOI222_X1 i_0_0_103 (.ZN (n_0_0_32), .A1 (\multiplicand[2] ), .A2 (hfn_ipo_n16), .B1 (n_0_0_64)
    , .B2 (n_0_65), .C1 (n_0_0_62), .C2 (B[1]));
INV_X1 i_0_0_102 (.ZN (\multiplicand_in[1] ), .A (n_0_0_32));
OR3_X1 i_0_0_101 (.ZN (n_0_0_30), .A1 (\counter[2] ), .A2 (\counter[1] ), .A3 (\counter[0] ));
OR2_X1 i_0_0_100 (.ZN (n_0_0_29), .A1 (n_0_0_30), .A2 (\counter[3] ));
NOR3_X1 i_0_0_99 (.ZN (n_0_0_28), .A1 (n_0_0_29), .A2 (ready), .A3 (\counter[4] ));
OR2_X1 i_0_0_98 (.ZN (n_0_161), .A1 (n_0_0_28), .A2 (n_0_258));
OR2_X1 i_0_0_97 (.ZN (n_0_160), .A1 (reset), .A2 (n_0_0_28));
XOR2_X1 i_0_0_96 (.Z (n_0_0_27), .A (\counter[4] ), .B (n_0_0_29));
OAI21_X1 i_0_0_95 (.ZN (\counter_in[4] ), .A (n_0_0_97), .B1 (n_0_0_27), .B2 (n_0_0_106));
XOR2_X1 i_0_0_94 (.Z (n_0_0_26), .A (\counter[3] ), .B (n_0_0_30));
OAI21_X1 i_0_0_93 (.ZN (\counter_in[3] ), .A (n_0_0_97), .B1 (n_0_0_26), .B2 (n_0_0_106));
OAI21_X1 i_0_0_92 (.ZN (n_0_0_25), .A (\counter[2] ), .B1 (\counter[1] ), .B2 (\counter[0] ));
AND2_X1 i_0_0_91 (.ZN (n_0_0_24), .A1 (n_0_0_30), .A2 (n_0_0_25));
OAI21_X1 i_0_0_90 (.ZN (\counter_in[2] ), .A (n_0_0_97), .B1 (n_0_0_24), .B2 (n_0_0_106));
XOR2_X1 i_0_0_89 (.Z (n_0_0_23), .A (\counter[1] ), .B (\counter[0] ));
OAI21_X1 i_0_0_88 (.ZN (\counter_in[1] ), .A (n_0_0_97), .B1 (n_0_0_23), .B2 (n_0_0_106));
OAI21_X1 i_0_0_87 (.ZN (\counter_in[0] ), .A (n_0_0_97), .B1 (n_0_0_106), .B2 (\counter[0] ));
NOR4_X1 i_0_0_86 (.ZN (n_0_0_22), .A1 (\multiplicand[7] ), .A2 (\multiplicand[6] )
    , .A3 (\multiplicand[5] ), .A4 (\multiplicand[4] ));
NOR4_X1 i_0_0_85 (.ZN (n_0_0_21), .A1 (\multiplicand[31] ), .A2 (\multiplicand[3] )
    , .A3 (\multiplicand[2] ), .A4 (\multiplicand[1] ));
NOR4_X1 i_0_0_84 (.ZN (n_0_0_20), .A1 (\multiplicand[14] ), .A2 (\multiplicand[13] )
    , .A3 (\multiplicand[12] ), .A4 (\multiplicand[8] ));
NOR4_X1 i_0_0_83 (.ZN (n_0_0_19), .A1 (\multiplicand[15] ), .A2 (\multiplicand[11] )
    , .A3 (\multiplicand[10] ), .A4 (\multiplicand[9] ));
NAND4_X1 i_0_0_82 (.ZN (n_0_0_18), .A1 (n_0_0_22), .A2 (n_0_0_21), .A3 (n_0_0_20), .A4 (n_0_0_19));
NOR4_X1 i_0_0_81 (.ZN (n_0_0_17), .A1 (\multiplicand[30] ), .A2 (\multiplicand[29] )
    , .A3 (\multiplicand[28] ), .A4 (\multiplicand[24] ));
NOR4_X1 i_0_0_80 (.ZN (n_0_0_16), .A1 (\multiplicand[27] ), .A2 (\multiplicand[26] )
    , .A3 (\multiplicand[25] ), .A4 (\multiplicand[16] ));
NOR4_X1 i_0_0_79 (.ZN (n_0_0_15), .A1 (\multiplicand[23] ), .A2 (\multiplicand[22] )
    , .A3 (\multiplicand[21] ), .A4 (\multiplicand[20] ));
NOR3_X1 i_0_0_78 (.ZN (n_0_0_14), .A1 (\multiplicand[19] ), .A2 (\multiplicand[18] ), .A3 (\multiplicand[17] ));
NAND4_X1 i_0_0_77 (.ZN (n_0_0_13), .A1 (n_0_0_17), .A2 (n_0_0_16), .A3 (n_0_0_15), .A4 (n_0_0_14));
NOR4_X1 i_0_0_76 (.ZN (n_0_0_12), .A1 (\accumulator[23] ), .A2 (\accumulator[22] )
    , .A3 (\accumulator[21] ), .A4 (\accumulator[20] ));
NOR4_X1 i_0_0_75 (.ZN (n_0_0_11), .A1 (\accumulator[19] ), .A2 (\accumulator[18] )
    , .A3 (\accumulator[17] ), .A4 (sgo__n20));
NOR4_X1 i_0_0_74 (.ZN (n_0_0_10), .A1 (\accumulator[30] ), .A2 (\accumulator[29] )
    , .A3 (\accumulator[28] ), .A4 (\accumulator[24] ));
NOR4_X1 i_0_0_73 (.ZN (n_0_0_9), .A1 (\accumulator[27] ), .A2 (\accumulator[26] )
    , .A3 (\accumulator[25] ), .A4 (\accumulator[16] ));
NAND4_X1 i_0_0_72 (.ZN (n_0_0_8), .A1 (n_0_0_12), .A2 (n_0_0_11), .A3 (n_0_0_10), .A4 (n_0_0_9));
NOR4_X1 i_0_0_71 (.ZN (n_0_0_7), .A1 (\accumulator[7] ), .A2 (\accumulator[6] ), .A3 (\accumulator[5] ), .A4 (\accumulator[4] ));
NOR4_X1 i_0_0_70 (.ZN (n_0_0_6), .A1 (\accumulator[3] ), .A2 (\accumulator[2] ), .A3 (\accumulator[1] ), .A4 (\accumulator[0] ));
NOR4_X1 i_0_0_69 (.ZN (n_0_0_5), .A1 (\accumulator[14] ), .A2 (\accumulator[13] )
    , .A3 (\accumulator[12] ), .A4 (\accumulator[8] ));
NOR4_X1 i_0_0_68 (.ZN (n_0_0_4), .A1 (\accumulator[15] ), .A2 (\accumulator[11] )
    , .A3 (\accumulator[10] ), .A4 (\accumulator[9] ));
NAND4_X1 i_0_0_67 (.ZN (n_0_0_3), .A1 (n_0_0_7), .A2 (n_0_0_6), .A3 (n_0_0_5), .A4 (n_0_0_4));
OR4_X1 i_0_0_66 (.ZN (n_0_0_2), .A1 (n_0_0_18), .A2 (n_0_0_13), .A3 (n_0_0_8), .A4 (n_0_0_3));
XNOR2_X1 i_0_0_65 (.ZN (n_0_0_1), .A (\isNeg[1] ), .B (n_0_0_101));
NAND2_X1 i_0_0_64 (.ZN (n_0_0_0), .A1 (n_0_0_2), .A2 (n_0_0_1));
AND3_X4 i_0_0_63 (.ZN (Res[63]), .A1 (n_0_0_2), .A2 (n_0_0_1), .A3 (n_0_158));
MUX2_X2 i_0_0_62 (.Z (Res[62]), .A (n_0_157), .B (\accumulator[30] ), .S (hfn_ipo_n13));
MUX2_X2 i_0_0_61 (.Z (Res[61]), .A (n_0_156), .B (\accumulator[29] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_60 (.Z (Res[60]), .A (n_0_155), .B (\accumulator[28] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_59 (.Z (Res[59]), .A (n_0_154), .B (\accumulator[27] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_58 (.Z (Res[58]), .A (n_0_153), .B (\accumulator[26] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_57 (.Z (Res[57]), .A (n_0_152), .B (\accumulator[25] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_56 (.Z (Res[56]), .A (n_0_151), .B (\accumulator[24] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_55 (.Z (Res[55]), .A (n_0_150), .B (\accumulator[23] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_54 (.Z (Res[54]), .A (n_0_149), .B (\accumulator[22] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_53 (.Z (Res[53]), .A (n_0_148), .B (\accumulator[21] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_52 (.Z (Res[52]), .A (n_0_147), .B (\accumulator[20] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_51 (.Z (Res[51]), .A (n_0_146), .B (\accumulator[19] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_50 (.Z (Res[50]), .A (n_0_145), .B (\accumulator[18] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_49 (.Z (Res[49]), .A (n_0_144), .B (\accumulator[17] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_48 (.Z (Res[48]), .A (n_0_143), .B (\accumulator[16] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_47 (.Z (Res[47]), .A (n_0_142), .B (\accumulator[15] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_46 (.Z (Res[46]), .A (n_0_141), .B (\accumulator[14] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_45 (.Z (Res[45]), .A (n_0_140), .B (\accumulator[13] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_44 (.Z (Res[44]), .A (n_0_139), .B (\accumulator[12] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_43 (.Z (Res[43]), .A (n_0_138), .B (\accumulator[11] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_42 (.Z (Res[42]), .A (n_0_137), .B (\accumulator[10] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_41 (.Z (Res[41]), .A (n_0_136), .B (\accumulator[9] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_40 (.Z (Res[40]), .A (n_0_135), .B (\accumulator[8] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_39 (.Z (Res[39]), .A (n_0_134), .B (\accumulator[7] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_38 (.Z (Res[38]), .A (n_0_133), .B (\accumulator[6] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_37 (.Z (Res[37]), .A (n_0_132), .B (\accumulator[5] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_36 (.Z (Res[36]), .A (n_0_131), .B (\accumulator[4] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_35 (.Z (Res[35]), .A (n_0_130), .B (\accumulator[3] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_34 (.Z (Res[34]), .A (n_0_129), .B (\accumulator[2] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_33 (.Z (Res[33]), .A (n_0_128), .B (\accumulator[1] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_32 (.Z (Res[32]), .A (n_0_127), .B (\accumulator[0] ), .S (hfn_ipo_n13));
MUX2_X1 i_0_0_31 (.Z (Res[31]), .A (n_0_126), .B (\multiplicand[31] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_30 (.Z (Res[30]), .A (n_0_125), .B (\multiplicand[30] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_29 (.Z (Res[29]), .A (n_0_124), .B (\multiplicand[29] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_28 (.Z (Res[28]), .A (n_0_123), .B (\multiplicand[28] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_27 (.Z (Res[27]), .A (n_0_122), .B (\multiplicand[27] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_26 (.Z (Res[26]), .A (n_0_121), .B (\multiplicand[26] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_25 (.Z (Res[25]), .A (n_0_120), .B (\multiplicand[25] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_24 (.Z (Res[24]), .A (n_0_119), .B (\multiplicand[24] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_23 (.Z (Res[23]), .A (n_0_118), .B (\multiplicand[23] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_22 (.Z (Res[22]), .A (n_0_117), .B (\multiplicand[22] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_21 (.Z (Res[21]), .A (n_0_116), .B (\multiplicand[21] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_20 (.Z (Res[20]), .A (n_0_115), .B (\multiplicand[20] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_19 (.Z (Res[19]), .A (n_0_114), .B (\multiplicand[19] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_18 (.Z (Res[18]), .A (n_0_113), .B (\multiplicand[18] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_17 (.Z (Res[17]), .A (n_0_112), .B (\multiplicand[17] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_16 (.Z (Res[16]), .A (n_0_111), .B (\multiplicand[16] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_15 (.Z (Res[15]), .A (n_0_110), .B (\multiplicand[15] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_14 (.Z (Res[14]), .A (n_0_109), .B (\multiplicand[14] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_13 (.Z (Res[13]), .A (n_0_108), .B (\multiplicand[13] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_12 (.Z (Res[12]), .A (n_0_107), .B (\multiplicand[12] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_11 (.Z (Res[11]), .A (n_0_106), .B (\multiplicand[11] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_10 (.Z (Res[10]), .A (n_0_105), .B (\multiplicand[10] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_9 (.Z (Res[9]), .A (n_0_104), .B (\multiplicand[9] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_8 (.Z (Res[8]), .A (n_0_103), .B (\multiplicand[8] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_7 (.Z (Res[7]), .A (n_0_102), .B (\multiplicand[7] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_6 (.Z (Res[6]), .A (n_0_101), .B (\multiplicand[6] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_5 (.Z (Res[5]), .A (n_0_100), .B (\multiplicand[5] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_4 (.Z (Res[4]), .A (n_0_99), .B (\multiplicand[4] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_3 (.Z (Res[3]), .A (n_0_98), .B (\multiplicand[3] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_2 (.Z (Res[2]), .A (n_0_97), .B (\multiplicand[2] ), .S (hfn_ipo_n14));
MUX2_X1 i_0_0_1 (.Z (Res[1]), .A (n_0_96), .B (\multiplicand[1] ), .S (hfn_ipo_n14));
NOR2_X4 i_0_0_0 (.ZN (OVF), .A1 (Res[63]), .A2 (n_0_0_101));
CLKGATETST_X4 clk_gate_isNeg_reg (.GCK (CTS_n_tid1_28), .CK (clk), .E (n_0_258), .SE (1'b0 ));
CLKGATETST_X8 clk_gate_accumulator_reg (.GCK (CTS_n_tid0_92), .CK (clk), .E (n_0_257), .SE (1'b0 ));
DFF_X1 \counter_reg[0]  (.Q (\counter[0] ), .CK (CTS_n_tid0_30), .D (\counter_in[0] ));
DFF_X1 \counter_reg[1]  (.Q (\counter[1] ), .CK (CTS_n_tid0_30), .D (\counter_in[1] ));
DFF_X1 \counter_reg[2]  (.Q (\counter[2] ), .CK (CTS_n_tid0_30), .D (\counter_in[2] ));
DFF_X1 \counter_reg[3]  (.Q (\counter[3] ), .CK (CTS_n_tid0_30), .D (\counter_in[3] ));
DFF_X1 \counter_reg[4]  (.Q (\counter[4] ), .CK (CTS_n_tid0_30), .D (\counter_in[4] ));
MUX2_X1 ready_reg_enable_mux_0 (.Z (n_0_159), .A (ready), .B (n_0_160), .S (n_0_161));
DFF_X1 ready_reg (.Q (ready), .CK (CTS_n_tid1_102), .D (n_0_159));
DFF_X1 \multiplicand_reg[0]  (.Q (drc_ipo_n18), .CK (CTS_n_tid0_30), .D (\multiplicand_in[0] ));
DFF_X1 \multiplicand_reg[1]  (.Q (\multiplicand[1] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[1] ));
DFF_X1 \multiplicand_reg[2]  (.Q (\multiplicand[2] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[2] ));
DFF_X1 \multiplicand_reg[3]  (.Q (\multiplicand[3] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[3] ));
DFF_X1 \multiplicand_reg[4]  (.Q (\multiplicand[4] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[4] ));
DFF_X1 \multiplicand_reg[5]  (.Q (\multiplicand[5] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[5] ));
DFF_X1 \multiplicand_reg[6]  (.Q (\multiplicand[6] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[6] ));
DFF_X1 \multiplicand_reg[7]  (.Q (\multiplicand[7] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[7] ));
DFF_X1 \multiplicand_reg[8]  (.Q (\multiplicand[8] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[8] ));
DFF_X1 \multiplicand_reg[9]  (.Q (\multiplicand[9] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[9] ));
DFF_X1 \multiplicand_reg[10]  (.Q (\multiplicand[10] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[10] ));
DFF_X1 \multiplicand_reg[11]  (.Q (\multiplicand[11] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[11] ));
DFF_X1 \multiplicand_reg[12]  (.Q (\multiplicand[12] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[12] ));
DFF_X1 \multiplicand_reg[13]  (.Q (\multiplicand[13] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[13] ));
DFF_X1 \multiplicand_reg[14]  (.Q (\multiplicand[14] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[14] ));
DFF_X1 \multiplicand_reg[15]  (.Q (\multiplicand[15] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[15] ));
DFF_X1 \multiplicand_reg[16]  (.Q (\multiplicand[16] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[16] ));
DFF_X1 \multiplicand_reg[17]  (.Q (\multiplicand[17] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[17] ));
DFF_X1 \multiplicand_reg[18]  (.Q (\multiplicand[18] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[18] ));
DFF_X1 \multiplicand_reg[19]  (.Q (\multiplicand[19] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[19] ));
DFF_X1 \multiplicand_reg[20]  (.Q (\multiplicand[20] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[20] ));
DFF_X1 \multiplicand_reg[21]  (.Q (\multiplicand[21] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[21] ));
DFF_X1 \multiplicand_reg[22]  (.Q (\multiplicand[22] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[22] ));
DFF_X1 \multiplicand_reg[23]  (.Q (\multiplicand[23] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[23] ));
DFF_X1 \multiplicand_reg[24]  (.Q (\multiplicand[24] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[24] ));
DFF_X1 \multiplicand_reg[25]  (.Q (\multiplicand[25] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[25] ));
DFF_X1 \multiplicand_reg[26]  (.Q (\multiplicand[26] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[26] ));
DFF_X1 \multiplicand_reg[27]  (.Q (\multiplicand[27] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[27] ));
DFF_X1 \multiplicand_reg[28]  (.Q (\multiplicand[28] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[28] ));
DFF_X1 \multiplicand_reg[29]  (.Q (\multiplicand[29] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[29] ));
DFF_X1 \multiplicand_reg[30]  (.Q (\multiplicand[30] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[30] ));
DFF_X1 \multiplicand_reg[31]  (.Q (\multiplicand[31] ), .CK (CTS_n_tid0_30), .D (\multiplicand_in[31] ));
DFF_X1 \multiplier_reg[0]  (.Q (\multiplier[0] ), .CK (CTS_n_tid1_31), .D (n_0_162));
DFF_X1 \multiplier_reg[1]  (.Q (\multiplier[1] ), .CK (CTS_n_tid1_31), .D (n_0_163));
DFF_X1 \multiplier_reg[2]  (.Q (\multiplier[2] ), .CK (CTS_n_tid1_31), .D (n_0_164));
DFF_X1 \multiplier_reg[3]  (.Q (\multiplier[3] ), .CK (CTS_n_tid1_31), .D (n_0_165));
DFF_X1 \multiplier_reg[4]  (.Q (\multiplier[4] ), .CK (CTS_n_tid1_31), .D (n_0_166));
DFF_X1 \multiplier_reg[5]  (.Q (\multiplier[5] ), .CK (CTS_n_tid1_31), .D (n_0_167));
DFF_X1 \multiplier_reg[6]  (.Q (\multiplier[6] ), .CK (CTS_n_tid1_31), .D (n_0_168));
DFF_X1 \multiplier_reg[7]  (.Q (\multiplier[7] ), .CK (CTS_n_tid1_31), .D (n_0_169));
DFF_X1 \multiplier_reg[8]  (.Q (\multiplier[8] ), .CK (CTS_n_tid1_31), .D (n_0_170));
DFF_X1 \multiplier_reg[9]  (.Q (\multiplier[9] ), .CK (CTS_n_tid1_31), .D (n_0_171));
DFF_X1 \multiplier_reg[10]  (.Q (\multiplier[10] ), .CK (CTS_n_tid1_31), .D (n_0_172));
DFF_X1 \multiplier_reg[11]  (.Q (\multiplier[11] ), .CK (CTS_n_tid1_31), .D (n_0_173));
DFF_X1 \multiplier_reg[12]  (.Q (\multiplier[12] ), .CK (CTS_n_tid1_31), .D (n_0_174));
DFF_X1 \multiplier_reg[13]  (.Q (\multiplier[13] ), .CK (CTS_n_tid1_31), .D (n_0_175));
DFF_X1 \multiplier_reg[14]  (.Q (\multiplier[14] ), .CK (CTS_n_tid1_31), .D (n_0_176));
DFF_X1 \multiplier_reg[15]  (.Q (\multiplier[15] ), .CK (CTS_n_tid1_31), .D (n_0_177));
DFF_X1 \multiplier_reg[16]  (.Q (\multiplier[16] ), .CK (CTS_n_tid1_32), .D (n_0_178));
DFF_X1 \multiplier_reg[17]  (.Q (\multiplier[17] ), .CK (CTS_n_tid1_32), .D (n_0_179));
DFF_X1 \multiplier_reg[18]  (.Q (\multiplier[18] ), .CK (CTS_n_tid1_32), .D (n_0_180));
DFF_X1 \multiplier_reg[19]  (.Q (\multiplier[19] ), .CK (CTS_n_tid1_32), .D (n_0_181));
DFF_X1 \multiplier_reg[20]  (.Q (\multiplier[20] ), .CK (CTS_n_tid1_32), .D (n_0_182));
DFF_X1 \multiplier_reg[21]  (.Q (\multiplier[21] ), .CK (CTS_n_tid1_32), .D (n_0_183));
DFF_X1 \multiplier_reg[22]  (.Q (\multiplier[22] ), .CK (CTS_n_tid1_32), .D (n_0_184));
DFF_X1 \multiplier_reg[23]  (.Q (\multiplier[23] ), .CK (CTS_n_tid1_32), .D (n_0_185));
DFF_X1 \multiplier_reg[24]  (.Q (\multiplier[24] ), .CK (CTS_n_tid1_32), .D (n_0_186));
DFF_X1 \multiplier_reg[25]  (.Q (\multiplier[25] ), .CK (CTS_n_tid1_32), .D (n_0_187));
DFF_X1 \multiplier_reg[26]  (.Q (\multiplier[26] ), .CK (CTS_n_tid1_32), .D (n_0_188));
DFF_X1 \multiplier_reg[27]  (.Q (\multiplier[27] ), .CK (CTS_n_tid1_32), .D (n_0_189));
DFF_X1 \multiplier_reg[28]  (.Q (\multiplier[28] ), .CK (CTS_n_tid1_32), .D (n_0_190));
DFF_X1 \multiplier_reg[29]  (.Q (\multiplier[29] ), .CK (CTS_n_tid1_32), .D (n_0_191));
DFF_X1 \multiplier_reg[30]  (.Q (\multiplier[30] ), .CK (CTS_n_tid1_32), .D (n_0_192));
DFF_X1 \multiplier_reg[31]  (.Q (\multiplier[31] ), .CK (CTS_n_tid1_32), .D (n_0_193));
DFF_X1 \accumulator_reg[0]  (.Q (\accumulator[0] ), .CK (CTS_n_tid0_29), .D (n_0_194));
DFF_X1 \accumulator_reg[1]  (.Q (\accumulator[1] ), .CK (CTS_n_tid0_29), .D (n_0_195));
DFF_X1 \accumulator_reg[2]  (.Q (\accumulator[2] ), .CK (CTS_n_tid0_29), .D (n_0_196));
DFF_X1 \accumulator_reg[3]  (.Q (\accumulator[3] ), .CK (CTS_n_tid0_29), .D (n_0_197));
DFF_X1 \accumulator_reg[4]  (.Q (\accumulator[4] ), .CK (CTS_n_tid0_29), .D (n_0_198));
DFF_X1 \accumulator_reg[5]  (.Q (\accumulator[5] ), .CK (CTS_n_tid0_29), .D (n_0_199));
DFF_X1 \accumulator_reg[6]  (.Q (\accumulator[6] ), .CK (CTS_n_tid0_29), .D (n_0_200));
DFF_X1 \accumulator_reg[7]  (.Q (\accumulator[7] ), .CK (CTS_n_tid0_29), .D (n_0_201));
DFF_X1 \accumulator_reg[8]  (.Q (\accumulator[8] ), .CK (CTS_n_tid0_29), .D (n_0_202));
DFF_X1 \accumulator_reg[9]  (.Q (\accumulator[9] ), .CK (CTS_n_tid0_29), .D (n_0_203));
DFF_X1 \accumulator_reg[10]  (.Q (\accumulator[10] ), .CK (CTS_n_tid0_29), .D (n_0_204));
DFF_X1 \accumulator_reg[11]  (.Q (\accumulator[11] ), .CK (CTS_n_tid0_29), .D (n_0_205));
DFF_X1 \accumulator_reg[12]  (.Q (\accumulator[12] ), .CK (CTS_n_tid0_29), .D (n_0_206));
DFF_X1 \accumulator_reg[13]  (.Q (\accumulator[13] ), .CK (CTS_n_tid0_29), .D (n_0_207));
DFF_X1 \accumulator_reg[14]  (.Q (\accumulator[14] ), .CK (CTS_n_tid0_29), .D (n_0_208));
DFF_X1 \accumulator_reg[15]  (.Q (\accumulator[15] ), .CK (CTS_n_tid0_29), .D (n_0_209));
DFF_X1 \accumulator_reg[16]  (.Q (\accumulator[16] ), .CK (CTS_n_tid0_29), .D (n_0_210));
DFF_X1 \accumulator_reg[17]  (.Q (\accumulator[17] ), .CK (CTS_n_tid0_29), .D (n_0_211));
DFF_X1 \accumulator_reg[18]  (.Q (\accumulator[18] ), .CK (CTS_n_tid0_29), .D (n_0_212));
DFF_X1 \accumulator_reg[19]  (.Q (\accumulator[19] ), .CK (CTS_n_tid0_29), .D (n_0_213));
DFF_X1 \accumulator_reg[20]  (.Q (\accumulator[20] ), .CK (CTS_n_tid0_29), .D (n_0_214));
DFF_X1 \accumulator_reg[21]  (.Q (\accumulator[21] ), .CK (CTS_n_tid0_29), .D (n_0_215));
DFF_X1 \accumulator_reg[22]  (.Q (\accumulator[22] ), .CK (CTS_n_tid0_29), .D (n_0_216));
DFF_X1 \accumulator_reg[23]  (.Q (\accumulator[23] ), .CK (CTS_n_tid0_29), .D (n_0_217));
DFF_X1 \accumulator_reg[24]  (.Q (\accumulator[24] ), .CK (CTS_n_tid0_29), .D (n_0_218));
DFF_X1 \accumulator_reg[25]  (.Q (\accumulator[25] ), .CK (CTS_n_tid0_29), .D (n_0_219));
DFF_X1 \accumulator_reg[26]  (.Q (\accumulator[26] ), .CK (CTS_n_tid0_29), .D (n_0_220));
DFF_X1 \accumulator_reg[27]  (.Q (\accumulator[27] ), .CK (CTS_n_tid0_29), .D (n_0_221));
DFF_X1 \accumulator_reg[28]  (.Q (\accumulator[28] ), .CK (CTS_n_tid0_29), .D (n_0_222));
DFF_X1 \accumulator_reg[29]  (.Q (\accumulator[29] ), .CK (CTS_n_tid0_30), .D (n_0_223));
DFF_X1 \accumulator_reg[30]  (.Q (\accumulator[30] ), .CK (CTS_n_tid0_30), .D (n_0_224));
DFF_X1 \isNeg_reg[0]  (.Q (\isNeg[0] ), .CK (CTS_n_tid1_32), .D (\isNeg_in[0] ));
DFF_X1 \isNeg_reg[1]  (.Q (\isNeg[1] ), .CK (CTS_n_tid1_32), .D (\isNeg_in[1] ));
datapath__0_13 i_0_16 (.p_0 ({n_0_158, n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, 
    n_0_152, n_0_151, n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, 
    n_0_143, n_0_142, n_0_141, n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, 
    n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, n_0_126, 
    n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, n_0_117, 
    n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, n_0_108, 
    n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, 
    n_0_98, n_0_97, n_0_96, uc_4}), .Res_imm ({uc_3, \accumulator[30] , \accumulator[29] , 
    \accumulator[28] , \accumulator[27] , \accumulator[26] , \accumulator[25] , \accumulator[24] , 
    \accumulator[23] , \accumulator[22] , \accumulator[21] , \accumulator[20] , \accumulator[19] , 
    \accumulator[18] , \accumulator[17] , \accumulator[16] , \accumulator[15] , \accumulator[14] , 
    \accumulator[13] , \accumulator[12] , \accumulator[11] , \accumulator[10] , \accumulator[9] , 
    \accumulator[8] , \accumulator[7] , \accumulator[6] , \accumulator[5] , \accumulator[4] , 
    \accumulator[3] , \accumulator[2] , \accumulator[1] , \accumulator[0] , \multiplicand[31] , 
    \multiplicand[30] , \multiplicand[29] , \multiplicand[28] , \multiplicand[27] , 
    \multiplicand[26] , \multiplicand[25] , \multiplicand[24] , \multiplicand[23] , 
    \multiplicand[22] , \multiplicand[21] , \multiplicand[20] , \multiplicand[19] , 
    \multiplicand[18] , \multiplicand[17] , \multiplicand[16] , \multiplicand[15] , 
    \multiplicand[14] , \multiplicand[13] , \multiplicand[12] , \multiplicand[11] , 
    \multiplicand[10] , \multiplicand[9] , \multiplicand[8] , \multiplicand[7] , 
    \multiplicand[6] , \multiplicand[5] , \multiplicand[4] , \multiplicand[3] , \multiplicand[2] , 
    \multiplicand[1] , sgo__n21}));
datapath__0_6 i_0_9 (.p_0 ({n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, 
    n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, 
    n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, 
    n_0_68, n_0_67, n_0_66, n_0_65, uc_2}), .B ({B[31], B[30], B[29], B[28], B[27], 
    B[26], B[25], B[24], B[23], B[22], B[21], B[20], B[19], B[18], B[17], B[16], 
    B[15], B[14], B[13], B[12], B[11], B[10], B[9], B[8], B[7], B[6], B[5], B[4], 
    B[3], B[2], B[1], B[0]}));
datapath__0_4 i_0_7 (.p_0 ({n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, 
    n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, 
    n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, 
    n_0_37, n_0_36, n_0_35, n_0_34, uc_1}), .A ({A[31], A[30], A[29], A[28], A[27], 
    A[26], A[25], A[24], A[23], A[22], A[21], A[20], A[19], A[18], A[17], A[16], 
    A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], 
    A[3], A[2], A[1], A[0]}));
datapath i_0_5 (.p_1 ({n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, 
    n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
    n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, 
    n_0_4, n_0_3, n_0_2}), .accumulator ({uc_0, \accumulator[30] , \accumulator[29] , 
    \accumulator[28] , \accumulator[27] , \accumulator[26] , \accumulator[25] , \accumulator[24] , 
    \accumulator[23] , \accumulator[22] , \accumulator[21] , \accumulator[20] , \accumulator[19] , 
    \accumulator[18] , \accumulator[17] , \accumulator[16] , \accumulator[15] , \accumulator[14] , 
    \accumulator[13] , \accumulator[12] , \accumulator[11] , \accumulator[10] , \accumulator[9] , 
    \accumulator[8] , \accumulator[7] , \accumulator[6] , \accumulator[5] , \accumulator[4] , 
    \accumulator[3] , \accumulator[2] , \accumulator[1] , \accumulator[0] }), .p_0 ({
    n_0_256, n_0_255, n_0_254, n_0_253, n_0_252, n_0_251, n_0_250, n_0_249, n_0_248, 
    n_0_247, n_0_246, n_0_245, n_0_244, n_0_243, n_0_242, n_0_241, n_0_240, n_0_239, 
    n_0_238, n_0_237, n_0_236, n_0_235, n_0_234, n_0_233, n_0_232, n_0_231, n_0_230, 
    n_0_229, n_0_228, n_0_227, n_0_226, n_0_225}));
CLKBUF_X2 hfn_ipo_c12 (.Z (hfn_ipo_n14), .A (n_0_0_0));
CLKBUF_X1 hfn_ipo_c13 (.Z (hfn_ipo_n15), .A (n_0_0_108));
CLKBUF_X2 hfn_ipo_c14 (.Z (hfn_ipo_n16), .A (n_0_0_108));
BUF_X8 drc_ipo_c15 (.Z (sgo__n21), .A (drc_ipo_n18));
CLKBUF_X2 hfn_ipo_c11 (.Z (hfn_ipo_n13), .A (n_0_0_0));
CLKBUF_X1 sgo__L2_c2_c16 (.Z (Res[0]), .A (sgo__n20));
CLKBUF_X1 sgo__L1_c1_c17 (.Z (sgo__n20), .A (sgo__n21));
CLKBUF_X3 CTS_L2_c_tid0_23 (.Z (CTS_n_tid0_29), .A (CTS_n_tid0_92));
CLKBUF_X3 CTS_L2_c_tid0_24 (.Z (CTS_n_tid0_30), .A (CTS_n_tid0_92));
CLKBUF_X3 CTS_L2_c_tid1_25 (.Z (CTS_n_tid1_31), .A (CTS_n_tid1_28));
CLKBUF_X3 CTS_L2_c_tid1_26 (.Z (CTS_n_tid1_32), .A (CTS_n_tid1_28));
CLKBUF_X1 CTS_L2_c_tid1_75 (.Z (CTS_n_tid1_102), .A (CTS_n_tid1_103));
CLKBUF_X1 CTS_L1_c_tid1_78 (.Z (CTS_n_tid1_103), .A (clk));

endmodule //sequentialMultiplier


