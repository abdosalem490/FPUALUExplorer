/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 16 23:31:31 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 532782118 */

module FA__1_917(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__1_913(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_909(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_905(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_901(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_897(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_893(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_889(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_885(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_881(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_877(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_873(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_869(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_865(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_861(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_857(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_853(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_849(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_845(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_841(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_837(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_833(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_829(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_825(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__1_1006(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__1_917 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__1_913 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__1_909 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__1_905 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__1_901 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__1_897 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__1_893 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__1_889 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__1_885 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__1_881 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__1_877 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__1_873 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__1_869 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__1_865 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__1_861 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(C[36]), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__1_857 genblk1_37_fa (.A(A[37]), .B(B[37]), .CIN(C[37]), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__1_853 genblk1_38_fa (.A(A[38]), .B(B[38]), .CIN(C[38]), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__1_849 genblk1_39_fa (.A(A[39]), .B(B[39]), .CIN(C[39]), .SUM(result[39]), 
      .COUT(carry[40]));
   FA__1_845 genblk1_40_fa (.A(A[40]), .B(B[40]), .CIN(C[40]), .SUM(result[40]), 
      .COUT(carry[41]));
   FA__1_841 genblk1_41_fa (.A(A[41]), .B(B[41]), .CIN(C[41]), .SUM(result[41]), 
      .COUT(carry[42]));
   FA__1_837 genblk1_42_fa (.A(A[42]), .B(B[42]), .CIN(C[42]), .SUM(result[42]), 
      .COUT(carry[43]));
   FA__1_833 genblk1_43_fa (.A(A[43]), .B(B[43]), .CIN(C[43]), .SUM(result[43]), 
      .COUT(carry[44]));
   FA__1_829 genblk1_44_fa (.A(A[44]), .B(B[44]), .CIN(C[44]), .SUM(result[44]), 
      .COUT(carry[45]));
   FA__1_825 genblk1_45_fa (.A(), .B(B[45]), .CIN(C[45]), .SUM(result[45]), 
      .COUT(carry[46]));
endmodule

module FA__1_1182(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__1_1178(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1174(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1170(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1166(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1162(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1158(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1154(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1150(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1146(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1142(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1138(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1134(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1130(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1126(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1122(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1118(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1114(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1110(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1106(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1102(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1098(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1094(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1090(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__1_1259(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__1_1182 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__1_1178 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__1_1174 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__1_1170 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__1_1166 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__1_1162 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__1_1158 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__1_1154 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__1_1150 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__1_1146 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__1_1142 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__1_1138 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__1_1134 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__1_1130 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__1_1126 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__1_1122 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__1_1118 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__1_1114 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(C[36]), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__1_1110 genblk1_37_fa (.A(A[37]), .B(B[37]), .CIN(C[37]), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__1_1106 genblk1_38_fa (.A(A[38]), .B(B[38]), .CIN(C[38]), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__1_1102 genblk1_39_fa (.A(A[39]), .B(B[39]), .CIN(C[39]), .SUM(result[39]), 
      .COUT(carry[40]));
   FA__1_1098 genblk1_40_fa (.A(A[40]), .B(B[40]), .CIN(C[40]), .SUM(result[40]), 
      .COUT(carry[41]));
   FA__1_1094 genblk1_41_fa (.A(A[41]), .B(B[41]), .CIN(C[41]), .SUM(result[41]), 
      .COUT(carry[42]));
   FA__1_1090 genblk1_42_fa (.A(), .B(B[42]), .CIN(C[42]), .SUM(result[42]), 
      .COUT(carry[43]));
endmodule

module FA__1_1447(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__1_1443(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1439(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1435(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1431(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1427(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1423(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1419(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1415(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1411(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1407(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1403(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1399(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1395(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1391(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1387(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1383(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1379(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1375(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1371(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1367(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1363(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1359(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1355(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__1_1512(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__1_1447 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__1_1443 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__1_1439 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__1_1435 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__1_1431 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__1_1427 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__1_1423 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__1_1419 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__1_1415 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__1_1411 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__1_1407 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__1_1403 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__1_1399 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__1_1395 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__1_1391 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__1_1387 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__1_1383 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__1_1379 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__1_1375 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__1_1371 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__1_1367 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(C[36]), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__1_1363 genblk1_37_fa (.A(A[37]), .B(B[37]), .CIN(C[37]), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__1_1359 genblk1_38_fa (.A(A[38]), .B(B[38]), .CIN(C[38]), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__1_1355 genblk1_39_fa (.A(), .B(B[39]), .CIN(C[39]), .SUM(result[39]), 
      .COUT(carry[40]));
endmodule

module FA__1_1712(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__1_1708(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1704(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1700(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1696(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1692(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1688(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1684(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1680(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1676(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1672(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1668(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1664(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1660(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1656(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1652(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1648(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1644(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1640(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1636(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1632(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1628(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1624(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1620(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__1_1765(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__1_1712 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__1_1708 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(C[14]), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__1_1704 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__1_1700 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__1_1696 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__1_1692 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__1_1688 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__1_1684 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__1_1680 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__1_1676 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__1_1672 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__1_1668 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__1_1664 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__1_1660 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__1_1656 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__1_1652 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__1_1648 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__1_1644 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__1_1640 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__1_1636 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__1_1632 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__1_1628 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__1_1624 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__1_1620 genblk1_36_fa (.A(), .B(B[36]), .CIN(C[36]), .SUM(result[36]), 
      .COUT(carry[37]));
endmodule

module FA__1_1977(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__1_1973(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1969(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1965(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1961(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1957(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1953(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1949(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1945(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1941(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1937(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1933(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1929(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1925(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1921(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1917(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1913(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1909(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1905(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1901(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1897(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1893(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1889(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_1885(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__1_2018(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__1_1977 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__1_1973 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(C[11]), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__1_1969 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(C[12]), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__1_1965 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(C[13]), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__1_1961 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(C[14]), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__1_1957 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__1_1953 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__1_1949 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__1_1945 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__1_1941 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__1_1937 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__1_1933 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__1_1929 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__1_1925 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__1_1921 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__1_1917 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__1_1913 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__1_1909 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__1_1905 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__1_1901 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__1_1897 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__1_1893 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__1_1889 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__1_1885 genblk1_33_fa (.A(), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
endmodule

module FA__1_2242(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__1_2238(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2234(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2230(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2226(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2222(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2218(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2214(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2210(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2206(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2202(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2198(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2194(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2190(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2186(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2182(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2178(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2174(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2170(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2166(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2162(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2158(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2154(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2150(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__1_2271(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__1_2242 genblk1_7_fa (.A(A[7]), .B(B[7]), .CIN(), .SUM(result[7]), 
      .COUT(carry[8]));
   FA__1_2238 genblk1_8_fa (.A(A[8]), .B(B[8]), .CIN(C[8]), .SUM(result[8]), 
      .COUT(carry[9]));
   FA__1_2234 genblk1_9_fa (.A(A[9]), .B(B[9]), .CIN(C[9]), .SUM(result[9]), 
      .COUT(carry[10]));
   FA__1_2230 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(C[10]), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__1_2226 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(C[11]), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__1_2222 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(C[12]), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__1_2218 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(C[13]), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__1_2214 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(C[14]), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__1_2210 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__1_2206 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__1_2202 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__1_2198 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__1_2194 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__1_2190 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__1_2186 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__1_2182 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__1_2178 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__1_2174 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__1_2170 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__1_2166 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__1_2162 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__1_2158 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__1_2154 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__1_2150 genblk1_30_fa (.A(), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
endmodule

module FA__1_2507(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__1_2503(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2499(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2495(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2491(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2487(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2483(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2479(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2475(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2471(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2467(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2463(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2459(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2455(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2451(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2447(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2443(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2439(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2435(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2431(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2427(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2423(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2419(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_2415(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__1_2524(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__1_2507 genblk1_4_fa (.A(A[4]), .B(B[4]), .CIN(), .SUM(result[4]), 
      .COUT(carry[5]));
   FA__1_2503 genblk1_5_fa (.A(A[5]), .B(B[5]), .CIN(C[5]), .SUM(result[5]), 
      .COUT(carry[6]));
   FA__1_2499 genblk1_6_fa (.A(A[6]), .B(B[6]), .CIN(C[6]), .SUM(result[6]), 
      .COUT(carry[7]));
   FA__1_2495 genblk1_7_fa (.A(A[7]), .B(B[7]), .CIN(C[7]), .SUM(result[7]), 
      .COUT(carry[8]));
   FA__1_2491 genblk1_8_fa (.A(A[8]), .B(B[8]), .CIN(C[8]), .SUM(result[8]), 
      .COUT(carry[9]));
   FA__1_2487 genblk1_9_fa (.A(A[9]), .B(B[9]), .CIN(C[9]), .SUM(result[9]), 
      .COUT(carry[10]));
   FA__1_2483 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(C[10]), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__1_2479 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(C[11]), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__1_2475 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(C[12]), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__1_2471 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(C[13]), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__1_2467 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(C[14]), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__1_2463 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__1_2459 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__1_2455 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__1_2451 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__1_2447 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__1_2443 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__1_2439 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__1_2435 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__1_2431 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__1_2427 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__1_2423 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__1_2419 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__1_2415 genblk1_27_fa (.A(), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
endmodule

module FA__1_7(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__1_11(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_15(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_19(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_23(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_27(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_31(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_35(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_39(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_43(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_47(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_51(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_55(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_59(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_63(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_67(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_71(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_75(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_79(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_83(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_87(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_91(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_95(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__1_99(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__0_108(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__1_7 genblk1_1_fa (.A(A[1]), .B(B[1]), .CIN(), .SUM(), .COUT(carry[2]));
   FA__1_11 genblk1_2_fa (.A(A[2]), .B(B[2]), .CIN(C[2]), .SUM(result[2]), 
      .COUT(carry[3]));
   FA__1_15 genblk1_3_fa (.A(A[3]), .B(B[3]), .CIN(C[3]), .SUM(result[3]), 
      .COUT(carry[4]));
   FA__1_19 genblk1_4_fa (.A(A[4]), .B(B[4]), .CIN(C[4]), .SUM(result[4]), 
      .COUT(carry[5]));
   FA__1_23 genblk1_5_fa (.A(A[5]), .B(B[5]), .CIN(C[5]), .SUM(result[5]), 
      .COUT(carry[6]));
   FA__1_27 genblk1_6_fa (.A(A[6]), .B(B[6]), .CIN(C[6]), .SUM(result[6]), 
      .COUT(carry[7]));
   FA__1_31 genblk1_7_fa (.A(A[7]), .B(B[7]), .CIN(C[7]), .SUM(result[7]), 
      .COUT(carry[8]));
   FA__1_35 genblk1_8_fa (.A(A[8]), .B(B[8]), .CIN(C[8]), .SUM(result[8]), 
      .COUT(carry[9]));
   FA__1_39 genblk1_9_fa (.A(A[9]), .B(B[9]), .CIN(C[9]), .SUM(result[9]), 
      .COUT(carry[10]));
   FA__1_43 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(C[10]), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__1_47 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(C[11]), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__1_51 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(C[12]), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__1_55 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(C[13]), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__1_59 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(C[14]), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__1_63 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__1_67 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__1_71 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__1_75 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__1_79 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__1_83 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__1_87 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__1_91 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__1_95 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__1_99 genblk1_24_fa (.A(), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
endmodule

module FA__2_925(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__2_921(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_917(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_913(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_909(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_905(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_901(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_897(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_893(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_889(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_885(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_881(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_877(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_873(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_869(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_865(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_861(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_857(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_853(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_849(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_845(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_841(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_837(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_833(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module CSAlike__2_1006(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__2_925 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__2_921 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__2_917 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__2_913 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__2_909 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__2_905 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__2_901 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__2_897 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__2_893 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__2_889 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__2_885 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__2_881 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__2_877 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__2_873 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__2_869 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__2_865 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__2_861 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(C[36]), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__2_857 genblk1_37_fa (.A(A[37]), .B(B[37]), .CIN(C[37]), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__2_853 genblk1_38_fa (.A(A[38]), .B(B[38]), .CIN(C[38]), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__2_849 genblk1_39_fa (.A(A[39]), .B(B[39]), .CIN(C[39]), .SUM(result[39]), 
      .COUT(carry[40]));
   FA__2_845 genblk1_40_fa (.A(A[40]), .B(B[40]), .CIN(C[40]), .SUM(result[40]), 
      .COUT(carry[41]));
   FA__2_841 genblk1_41_fa (.A(A[41]), .B(B[41]), .CIN(C[41]), .SUM(result[41]), 
      .COUT(carry[42]));
   FA__2_837 genblk1_42_fa (.A(A[42]), .B(B[42]), .CIN(C[42]), .SUM(result[42]), 
      .COUT(carry[43]));
   FA__2_833 genblk1_43_fa (.A(A[43]), .B(B[43]), .CIN(C[43]), .SUM(result[43]), 
      .COUT(carry[44]));
endmodule

module FA__2_1198(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__2_1194(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__2_1190(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1186(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1182(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1178(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1174(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1170(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1166(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1162(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1158(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1154(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1150(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1146(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1142(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1138(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1134(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1130(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1126(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1122(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1118(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1114(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1110(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1106(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__2_1102(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__2_1098(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__2_1259(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__2_1198 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__2_1194 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__2_1190 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__2_1186 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__2_1182 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__2_1178 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__2_1174 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__2_1170 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__2_1166 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__2_1162 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__2_1158 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__2_1154 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__2_1150 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__2_1146 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__2_1142 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__2_1138 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__2_1134 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__2_1130 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__2_1126 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__2_1122 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__2_1118 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__2_1114 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(C[36]), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__2_1110 genblk1_37_fa (.A(A[37]), .B(B[37]), .CIN(C[37]), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__2_1106 genblk1_38_fa (.A(), .B(B[38]), .CIN(C[38]), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__2_1102 genblk1_39_fa (.A(), .B(B[39]), .CIN(C[39]), .SUM(result[39]), 
      .COUT(carry[40]));
   FA__2_1098 genblk1_40_fa (.A(), .B(B[40]), .CIN(C[40]), .SUM(result[40]), 
      .COUT(carry[41]));
endmodule

module FA__2_1467(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__2_1463(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1459(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1455(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1451(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1447(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1443(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1439(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1435(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1431(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1427(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1423(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1419(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1415(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1411(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1407(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1403(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1399(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1395(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1391(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1387(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1383(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1379(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1375(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module CSAlike__2_1512(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__2_1467 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__2_1463 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(C[12]), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__2_1459 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(C[13]), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__2_1455 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(C[14]), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__2_1451 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__2_1447 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__2_1443 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__2_1439 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__2_1435 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__2_1431 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__2_1427 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__2_1423 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__2_1419 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__2_1415 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__2_1411 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__2_1407 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__2_1403 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__2_1399 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__2_1395 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__2_1391 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__2_1387 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__2_1383 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__2_1379 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__2_1375 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
endmodule

module FA__2_1740(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__2_1736(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__2_1732(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1728(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1724(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1720(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1716(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1712(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1708(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1704(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1700(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1696(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1692(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1688(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1684(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1680(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1676(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1672(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1668(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1664(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1660(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1656(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1652(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_1648(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__2_1644(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__2_1640(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__2_1765(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__2_1740 genblk1_6_fa (.A(A[6]), .B(B[6]), .CIN(), .SUM(result[6]), 
      .COUT(carry[7]));
   FA__2_1736 genblk1_7_fa (.A(A[7]), .B(B[7]), .CIN(), .SUM(result[7]), 
      .COUT(carry[8]));
   FA__2_1732 genblk1_8_fa (.A(A[8]), .B(B[8]), .CIN(C[8]), .SUM(result[8]), 
      .COUT(carry[9]));
   FA__2_1728 genblk1_9_fa (.A(A[9]), .B(B[9]), .CIN(C[9]), .SUM(result[9]), 
      .COUT(carry[10]));
   FA__2_1724 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(C[10]), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__2_1720 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(C[11]), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__2_1716 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(C[12]), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__2_1712 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(C[13]), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__2_1708 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(C[14]), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__2_1704 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__2_1700 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__2_1696 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__2_1692 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__2_1688 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__2_1684 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__2_1680 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__2_1676 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__2_1672 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__2_1668 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__2_1664 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__2_1660 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__2_1656 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__2_1652 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__2_1648 genblk1_29_fa (.A(), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__2_1644 genblk1_30_fa (.A(), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__2_1640 genblk1_31_fa (.A(), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
endmodule

module FA__2_11(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__2_15(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_19(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_23(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_27(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_31(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_35(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_39(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_43(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_47(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_51(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_55(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_59(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_63(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_67(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_71(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_75(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_79(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_83(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_87(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_91(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_95(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_99(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__2_103(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module CSAlike__0_113(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__2_11 genblk1_2_fa (.A(A[2]), .B(B[2]), .CIN(), .SUM(), .COUT(carry[3]));
   FA__2_15 genblk1_3_fa (.A(A[3]), .B(B[3]), .CIN(C[3]), .SUM(result[3]), 
      .COUT(carry[4]));
   FA__2_19 genblk1_4_fa (.A(A[4]), .B(B[4]), .CIN(C[4]), .SUM(result[4]), 
      .COUT(carry[5]));
   FA__2_23 genblk1_5_fa (.A(A[5]), .B(B[5]), .CIN(C[5]), .SUM(result[5]), 
      .COUT(carry[6]));
   FA__2_27 genblk1_6_fa (.A(A[6]), .B(B[6]), .CIN(C[6]), .SUM(result[6]), 
      .COUT(carry[7]));
   FA__2_31 genblk1_7_fa (.A(A[7]), .B(B[7]), .CIN(C[7]), .SUM(result[7]), 
      .COUT(carry[8]));
   FA__2_35 genblk1_8_fa (.A(A[8]), .B(B[8]), .CIN(C[8]), .SUM(result[8]), 
      .COUT(carry[9]));
   FA__2_39 genblk1_9_fa (.A(A[9]), .B(B[9]), .CIN(C[9]), .SUM(result[9]), 
      .COUT(carry[10]));
   FA__2_43 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(C[10]), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__2_47 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(C[11]), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__2_51 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(C[12]), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__2_55 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(C[13]), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__2_59 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(C[14]), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__2_63 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__2_67 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__2_71 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__2_75 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__2_79 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__2_83 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__2_87 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__2_91 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__2_95 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__2_99 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__2_103 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
endmodule

module FA__3_660(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__3_656(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__3_652(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_648(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_644(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_640(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_636(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_632(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_628(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_624(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_620(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_616(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_612(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_608(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_604(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_600(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_596(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_592(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_588(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_584(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_580(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__3_576(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module CSAlike__3_753(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__3_660 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__3_656 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__3_652 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__3_648 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__3_644 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__3_640 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__3_636 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__3_632 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__3_628 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__3_624 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__3_620 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__3_616 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__3_612 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__3_608 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__3_604 genblk1_37_fa (.A(A[37]), .B(B[37]), .CIN(), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__3_600 genblk1_38_fa (.A(A[38]), .B(B[38]), .CIN(), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__3_596 genblk1_39_fa (.A(A[39]), .B(B[39]), .CIN(), .SUM(result[39]), 
      .COUT(carry[40]));
   FA__3_592 genblk1_40_fa (.A(A[40]), .B(B[40]), .CIN(), .SUM(result[40]), 
      .COUT(carry[41]));
   FA__3_588 genblk1_41_fa (.A(A[41]), .B(B[41]), .CIN(), .SUM(result[41]), 
      .COUT(carry[42]));
   FA__3_584 genblk1_42_fa (.A(A[42]), .B(B[42]), .CIN(), .SUM(result[42]), 
      .COUT(carry[43]));
   FA__3_580 genblk1_43_fa (.A(A[43]), .B(B[43]), .CIN(), .SUM(result[43]), 
      .COUT(carry[44]));
   FA__3_576 genblk1_44_fa (.A(A[44]), .B(B[44]), .CIN(), .SUM(result[44]), 
      .COUT(carry[45]));
endmodule

module FA__3_941(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__3_937(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__3_933(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_929(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_925(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_921(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_917(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_913(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_909(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_905(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_901(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_897(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_893(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_889(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_885(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_881(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_877(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_873(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_869(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_865(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_861(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_857(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_853(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_849(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_845(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_841(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__3_1006(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__3_941 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__3_937 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__3_933 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__3_929 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__3_925 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__3_921 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__3_917 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__3_913 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__3_909 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__3_905 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__3_901 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__3_897 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__3_893 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__3_889 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__3_885 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__3_881 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__3_877 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__3_873 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__3_869 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__3_865 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__3_861 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(C[36]), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__3_857 genblk1_37_fa (.A(A[37]), .B(B[37]), .CIN(C[37]), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__3_853 genblk1_38_fa (.A(A[38]), .B(B[38]), .CIN(C[38]), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__3_849 genblk1_39_fa (.A(A[39]), .B(B[39]), .CIN(C[39]), .SUM(result[39]), 
      .COUT(carry[40]));
   FA__3_845 genblk1_40_fa (.A(A[40]), .B(B[40]), .CIN(C[40]), .SUM(result[40]), 
      .COUT(carry[41]));
   FA__3_841 genblk1_41_fa (.A(), .B(B[41]), .CIN(C[41]), .SUM(result[41]), 
      .COUT(carry[42]));
endmodule

module FA__3_1222(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__3_1218(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__3_1214(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__3_1210(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1206(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1202(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1198(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1194(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1190(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1186(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1182(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1178(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1174(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1170(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1166(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1162(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1158(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1154(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1150(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1146(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1142(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1138(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1134(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1130(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_1126(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__3_1122(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__3_1118(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__3_1259(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__3_1222 genblk1_9_fa (.A(A[9]), .B(B[9]), .CIN(), .SUM(result[9]), 
      .COUT(carry[10]));
   FA__3_1218 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__3_1214 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__3_1210 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(C[12]), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__3_1206 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(C[13]), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__3_1202 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(C[14]), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__3_1198 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__3_1194 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__3_1190 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__3_1186 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__3_1182 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__3_1178 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__3_1174 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__3_1170 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__3_1166 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__3_1162 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__3_1158 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__3_1154 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__3_1150 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__3_1146 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__3_1142 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__3_1138 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__3_1134 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__3_1130 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__3_1126 genblk1_33_fa (.A(), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__3_1122 genblk1_34_fa (.A(), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__3_1118 genblk1_35_fa (.A(), .B(B[35]), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
endmodule

module FA__3_15(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__3_19(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__3_23(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_27(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_31(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_35(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_39(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_43(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_47(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_51(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_55(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_59(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_63(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_67(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_71(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_75(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_79(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_83(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_87(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_91(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_95(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_99(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_103(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_107(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__3_111(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__3_115(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module CSAlike__0_118(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__3_15 genblk1_3_fa (.A(A[3]), .B(B[3]), .CIN(), .SUM(), .COUT(carry[4]));
   FA__3_19 genblk1_4_fa (.A(A[4]), .B(B[4]), .CIN(), .SUM(result[4]), .COUT(
      carry[5]));
   FA__3_23 genblk1_5_fa (.A(A[5]), .B(B[5]), .CIN(C[5]), .SUM(result[5]), 
      .COUT(carry[6]));
   FA__3_27 genblk1_6_fa (.A(A[6]), .B(B[6]), .CIN(C[6]), .SUM(result[6]), 
      .COUT(carry[7]));
   FA__3_31 genblk1_7_fa (.A(A[7]), .B(B[7]), .CIN(C[7]), .SUM(result[7]), 
      .COUT(carry[8]));
   FA__3_35 genblk1_8_fa (.A(A[8]), .B(B[8]), .CIN(C[8]), .SUM(result[8]), 
      .COUT(carry[9]));
   FA__3_39 genblk1_9_fa (.A(A[9]), .B(B[9]), .CIN(C[9]), .SUM(result[9]), 
      .COUT(carry[10]));
   FA__3_43 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(C[10]), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__3_47 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(C[11]), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__3_51 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(C[12]), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__3_55 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(C[13]), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__3_59 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(C[14]), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__3_63 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__3_67 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__3_71 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__3_75 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__3_79 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__3_83 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__3_87 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__3_91 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__3_95 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__3_99 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__3_103 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__3_107 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__3_111 genblk1_27_fa (.A(A[27]), .B(), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__3_115 genblk1_28_fa (.A(A[28]), .B(), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
endmodule

module FA__4_403(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_399(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_395(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_391(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_387(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_383(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_379(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_375(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_371(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_367(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_363(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_359(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_355(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_351(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_347(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_343(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_339(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_335(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_331(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_327(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_323(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_319(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module CSAlike__4_500(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__4_403 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__4_399 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__4_395 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__4_391 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__4_387 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__4_383 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__4_379 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__4_375 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__4_371 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__4_367 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__4_363 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__4_359 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__4_355 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__4_351 genblk1_37_fa (.A(A[37]), .B(B[37]), .CIN(), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__4_347 genblk1_38_fa (.A(A[38]), .B(B[38]), .CIN(), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__4_343 genblk1_39_fa (.A(A[39]), .B(B[39]), .CIN(), .SUM(result[39]), 
      .COUT(carry[40]));
   FA__4_339 genblk1_40_fa (.A(A[40]), .B(B[40]), .CIN(), .SUM(result[40]), 
      .COUT(carry[41]));
   FA__4_335 genblk1_41_fa (.A(A[41]), .B(B[41]), .CIN(), .SUM(result[41]), 
      .COUT(carry[42]));
   FA__4_331 genblk1_42_fa (.A(A[42]), .B(B[42]), .CIN(), .SUM(result[42]), 
      .COUT(carry[43]));
   FA__4_327 genblk1_43_fa (.A(A[43]), .B(B[43]), .CIN(), .SUM(result[43]), 
      .COUT(carry[44]));
   FA__4_323 genblk1_44_fa (.A(A[44]), .B(B[44]), .CIN(), .SUM(result[44]), 
      .COUT(carry[45]));
   FA__4_319 genblk1_45_fa (.A(A[45]), .B(B[45]), .CIN(), .SUM(result[45]), 
      .COUT(carry[46]));
endmodule

module FA__4_696(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_692(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_688(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_684(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_680(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_676(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_672(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_668(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_664(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_660(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_656(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_652(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_648(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_644(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_640(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_636(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_632(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_628(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_624(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_620(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_616(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_612(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_608(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_604(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__4_600(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__4_596(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__4_592(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__4_588(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__4_584(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__4_753(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__4_696 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__4_692 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__4_688 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__4_684 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__4_680 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__4_676 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__4_672 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__4_668 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__4_664 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__4_660 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__4_656 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__4_652 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__4_648 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__4_644 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__4_640 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__4_636 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__4_632 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__4_628 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__4_624 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__4_620 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__4_616 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__4_612 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__4_608 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(C[36]), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__4_604 genblk1_37_fa (.A(), .B(B[37]), .CIN(C[37]), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__4_600 genblk1_38_fa (.A(), .B(B[38]), .CIN(C[38]), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__4_596 genblk1_39_fa (.A(), .B(B[39]), .CIN(C[39]), .SUM(result[39]), 
      .COUT(carry[40]));
   FA__4_592 genblk1_40_fa (.A(), .B(B[40]), .CIN(C[40]), .SUM(result[40]), 
      .COUT(carry[41]));
   FA__4_588 genblk1_41_fa (.A(), .B(B[41]), .CIN(C[41]), .SUM(result[41]), 
      .COUT(carry[42]));
   FA__4_584 genblk1_42_fa (.A(), .B(B[42]), .CIN(C[42]), .SUM(result[42]), 
      .COUT(carry[43]));
endmodule

module FA__4_989(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_985(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_981(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_977(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_973(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_969(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_965(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_961(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_957(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_953(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_949(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_945(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_941(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_937(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_933(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_929(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_925(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_921(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_917(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_913(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_909(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_905(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_901(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_897(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_893(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_889(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_885(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__4_881(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module CSAlike__4_1006(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__4_989 genblk1_4_fa (.A(A[4]), .B(B[4]), .CIN(), .SUM(), .COUT(carry[5]));
   FA__4_985 genblk1_5_fa (.A(A[5]), .B(B[5]), .CIN(), .SUM(result[5]), .COUT(
      carry[6]));
   FA__4_981 genblk1_6_fa (.A(A[6]), .B(B[6]), .CIN(), .SUM(result[6]), .COUT(
      carry[7]));
   FA__4_977 genblk1_7_fa (.A(A[7]), .B(B[7]), .CIN(C[7]), .SUM(result[7]), 
      .COUT(carry[8]));
   FA__4_973 genblk1_8_fa (.A(A[8]), .B(B[8]), .CIN(C[8]), .SUM(result[8]), 
      .COUT(carry[9]));
   FA__4_969 genblk1_9_fa (.A(A[9]), .B(B[9]), .CIN(C[9]), .SUM(result[9]), 
      .COUT(carry[10]));
   FA__4_965 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(C[10]), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__4_961 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(C[11]), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__4_957 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(C[12]), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__4_953 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(C[13]), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__4_949 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(C[14]), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__4_945 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__4_941 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__4_937 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__4_933 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__4_929 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__4_925 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__4_921 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__4_917 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__4_913 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__4_909 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__4_905 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__4_901 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__4_897 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__4_893 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__4_889 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__4_885 genblk1_30_fa (.A(A[30]), .B(), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__4_881 genblk1_31_fa (.A(A[31]), .B(), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
endmodule

module FA__4_1174(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1170(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1166(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1162(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1158(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1154(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1150(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1146(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1142(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1138(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1134(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1130(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1126(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1122(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1118(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1114(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1110(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1106(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1102(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1098(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1094(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1090(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1086(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1082(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__4_1078(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module FA__4_1074(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__4_1259(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__4_1174 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__4_1170 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__4_1166 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__4_1162 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__4_1158 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__4_1154 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__4_1150 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__4_1146 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__4_1142 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__4_1138 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__4_1134 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__4_1130 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__4_1126 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__4_1122 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__4_1118 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__4_1114 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(C[36]), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__4_1110 genblk1_37_fa (.A(A[37]), .B(B[37]), .CIN(C[37]), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__4_1106 genblk1_38_fa (.A(A[38]), .B(B[38]), .CIN(C[38]), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__4_1102 genblk1_39_fa (.A(A[39]), .B(B[39]), .CIN(C[39]), .SUM(result[39]), 
      .COUT(carry[40]));
   FA__4_1098 genblk1_40_fa (.A(A[40]), .B(B[40]), .CIN(C[40]), .SUM(result[40]), 
      .COUT(carry[41]));
   FA__4_1094 genblk1_41_fa (.A(A[41]), .B(B[41]), .CIN(C[41]), .SUM(result[41]), 
      .COUT(carry[42]));
   FA__4_1090 genblk1_42_fa (.A(A[42]), .B(B[42]), .CIN(C[42]), .SUM(result[42]), 
      .COUT(carry[43]));
   FA__4_1086 genblk1_43_fa (.A(A[43]), .B(B[43]), .CIN(C[43]), .SUM(result[43]), 
      .COUT(carry[44]));
   FA__4_1082 genblk1_44_fa (.A(), .B(B[44]), .CIN(C[44]), .SUM(result[44]), 
      .COUT(carry[45]));
   FA__4_1078 genblk1_45_fa (.A(), .B(B[45]), .CIN(C[45]), .SUM(result[45]), 
      .COUT(carry[46]));
   FA__4_1074 genblk1_46_fa (.A(), .B(B[46]), .CIN(C[46]), .SUM(result[46]), 
      .COUT(carry[47]));
endmodule

module FA__4_1491(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1487(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1483(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1479(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1475(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1471(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1467(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1463(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1459(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1455(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1451(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1447(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1443(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1439(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1435(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1431(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1427(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1423(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1419(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1415(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1411(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1407(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1403(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1399(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1395(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1391(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1387(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1383(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1379(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__4_1375(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__4_1371(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__4_1367(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__4_1363(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module CSAlike__4_1512(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__4_1491 genblk1_5_fa (.A(A[5]), .B(B[5]), .CIN(), .SUM(), .COUT(carry[6]));
   FA__4_1487 genblk1_6_fa (.A(A[6]), .B(B[6]), .CIN(), .SUM(result[6]), 
      .COUT(carry[7]));
   FA__4_1483 genblk1_7_fa (.A(A[7]), .B(B[7]), .CIN(), .SUM(result[7]), 
      .COUT(carry[8]));
   FA__4_1479 genblk1_8_fa (.A(A[8]), .B(B[8]), .CIN(), .SUM(result[8]), 
      .COUT(carry[9]));
   FA__4_1475 genblk1_9_fa (.A(A[9]), .B(B[9]), .CIN(), .SUM(result[9]), 
      .COUT(carry[10]));
   FA__4_1471 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(C[10]), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__4_1467 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(C[11]), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__4_1463 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(C[12]), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__4_1459 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(C[13]), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__4_1455 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(C[14]), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__4_1451 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__4_1447 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__4_1443 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__4_1439 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__4_1435 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__4_1431 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__4_1427 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__4_1423 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__4_1419 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__4_1415 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__4_1411 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__4_1407 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__4_1403 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__4_1399 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__4_1395 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__4_1391 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__4_1387 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__4_1383 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__4_1379 genblk1_33_fa (.A(A[33]), .B(), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__4_1375 genblk1_34_fa (.A(A[34]), .B(), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__4_1371 genblk1_35_fa (.A(A[35]), .B(), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__4_1367 genblk1_36_fa (.A(A[36]), .B(), .CIN(C[36]), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__4_1363 genblk1_37_fa (.A(A[37]), .B(), .CIN(C[37]), .SUM(result[37]), 
      .COUT(carry[38]));
endmodule

module FA__4_1740(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1736(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1732(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1728(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1724(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1720(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1716(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1712(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1708(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1704(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1700(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1696(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1692(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1688(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1684(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1680(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1676(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1672(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1668(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1664(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1660(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1656(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1652(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1648(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1644(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1640(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1636(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1632(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1628(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1624(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1620(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1616(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1612(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1608(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__4_1604(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__4_1600(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__4_1596(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__4_1592(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__4_1588(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__4_1584(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(A), .A2(CIN), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(A), .B(CIN), .Z(SUM));
endmodule

module FA__4_1580(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(CIN), .Z(SUM));
   AND2_X1 i_0_1 (.A1(CIN), .A2(A), .ZN(COUT));
endmodule

module CSAlike__4_1765(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__4_1740 genblk1_6_fa (.A(A[6]), .B(B[6]), .CIN(), .SUM(), .COUT(carry[7]));
   FA__4_1736 genblk1_7_fa (.A(A[7]), .B(B[7]), .CIN(), .SUM(result[7]), 
      .COUT(carry[8]));
   FA__4_1732 genblk1_8_fa (.A(A[8]), .B(B[8]), .CIN(), .SUM(result[8]), 
      .COUT(carry[9]));
   FA__4_1728 genblk1_9_fa (.A(A[9]), .B(B[9]), .CIN(), .SUM(result[9]), 
      .COUT(carry[10]));
   FA__4_1724 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__4_1720 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__4_1716 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__4_1712 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__4_1708 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__4_1704 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(C[15]), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__4_1700 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(C[16]), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__4_1696 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(C[17]), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__4_1692 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(C[18]), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__4_1688 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(C[19]), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__4_1684 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(C[20]), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__4_1680 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(C[21]), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__4_1676 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__4_1672 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__4_1668 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__4_1664 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__4_1660 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__4_1656 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__4_1652 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__4_1648 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__4_1644 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__4_1640 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__4_1636 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__4_1632 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__4_1628 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__4_1624 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__4_1620 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(C[36]), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__4_1616 genblk1_37_fa (.A(A[37]), .B(B[37]), .CIN(C[37]), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__4_1612 genblk1_38_fa (.A(A[38]), .B(B[38]), .CIN(C[38]), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__4_1608 genblk1_39_fa (.A(A[39]), .B(), .CIN(C[39]), .SUM(result[39]), 
      .COUT(carry[40]));
   FA__4_1604 genblk1_40_fa (.A(A[40]), .B(), .CIN(C[40]), .SUM(result[40]), 
      .COUT(carry[41]));
   FA__4_1600 genblk1_41_fa (.A(A[41]), .B(), .CIN(C[41]), .SUM(result[41]), 
      .COUT(carry[42]));
   FA__4_1596 genblk1_42_fa (.A(A[42]), .B(), .CIN(C[42]), .SUM(result[42]), 
      .COUT(carry[43]));
   FA__4_1592 genblk1_43_fa (.A(A[43]), .B(), .CIN(C[43]), .SUM(result[43]), 
      .COUT(carry[44]));
   FA__4_1588 genblk1_44_fa (.A(A[44]), .B(), .CIN(C[44]), .SUM(result[44]), 
      .COUT(carry[45]));
   FA__4_1584 genblk1_45_fa (.A(A[45]), .B(), .CIN(C[45]), .SUM(result[45]), 
      .COUT(carry[46]));
   FA__4_1580 genblk1_46_fa (.A(A[46]), .B(), .CIN(C[46]), .SUM(result[46]), 
      .COUT(carry[47]));
endmodule

module FA__4_1989(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1985(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1981(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1977(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1973(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1969(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1965(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1961(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1957(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1953(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1949(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1945(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1941(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1937(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1933(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_1929(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1925(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1921(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1917(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1913(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1909(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1905(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1901(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1897(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1893(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1889(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1885(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1881(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1877(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1873(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1869(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1865(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1861(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1857(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1853(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1849(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1845(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1841(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1837(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1833(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   wire temp;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(temp));
   XOR2_X1 i_0_1 (.A(temp), .B(CIN), .Z(SUM));
   AOI22_X1 i_0_2 (.A1(A), .A2(B), .B1(temp), .B2(CIN), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(COUT));
endmodule

module FA__4_1829(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_1 (.A(B), .B(CIN), .Z(SUM));
endmodule

module CSAlike__4_2018(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__4_1989 genblk1_7_fa (.A(A[7]), .B(B[7]), .CIN(), .SUM(), .COUT(carry[8]));
   FA__4_1985 genblk1_8_fa (.A(A[8]), .B(B[8]), .CIN(), .SUM(result[8]), 
      .COUT(carry[9]));
   FA__4_1981 genblk1_9_fa (.A(A[9]), .B(B[9]), .CIN(), .SUM(result[9]), 
      .COUT(carry[10]));
   FA__4_1977 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__4_1973 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__4_1969 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__4_1965 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__4_1961 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__4_1957 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__4_1953 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__4_1949 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__4_1945 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__4_1941 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__4_1937 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__4_1933 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__4_1929 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(C[22]), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__4_1925 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(C[23]), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__4_1921 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(C[24]), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__4_1917 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(C[25]), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__4_1913 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(C[26]), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__4_1909 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(C[27]), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__4_1905 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(C[28]), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__4_1901 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(C[29]), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__4_1897 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(C[30]), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__4_1893 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(C[31]), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__4_1889 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(C[32]), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__4_1885 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(C[33]), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__4_1881 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(C[34]), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__4_1877 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(C[35]), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__4_1873 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(C[36]), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__4_1869 genblk1_37_fa (.A(A[37]), .B(B[37]), .CIN(C[37]), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__4_1865 genblk1_38_fa (.A(A[38]), .B(B[38]), .CIN(C[38]), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__4_1861 genblk1_39_fa (.A(A[39]), .B(B[39]), .CIN(C[39]), .SUM(result[39]), 
      .COUT(carry[40]));
   FA__4_1857 genblk1_40_fa (.A(A[40]), .B(B[40]), .CIN(C[40]), .SUM(result[40]), 
      .COUT(carry[41]));
   FA__4_1853 genblk1_41_fa (.A(A[41]), .B(B[41]), .CIN(C[41]), .SUM(result[41]), 
      .COUT(carry[42]));
   FA__4_1849 genblk1_42_fa (.A(A[42]), .B(B[42]), .CIN(C[42]), .SUM(result[42]), 
      .COUT(carry[43]));
   FA__4_1845 genblk1_43_fa (.A(A[43]), .B(B[43]), .CIN(C[43]), .SUM(result[43]), 
      .COUT(carry[44]));
   FA__4_1841 genblk1_44_fa (.A(A[44]), .B(B[44]), .CIN(C[44]), .SUM(result[44]), 
      .COUT(carry[45]));
   FA__4_1837 genblk1_45_fa (.A(A[45]), .B(B[45]), .CIN(C[45]), .SUM(result[45]), 
      .COUT(carry[46]));
   FA__4_1833 genblk1_46_fa (.A(A[46]), .B(B[46]), .CIN(C[46]), .SUM(result[46]), 
      .COUT(carry[47]));
   FA__4_1829 genblk1_47_fa (.A(), .B(B[47]), .CIN(C[47]), .SUM(result[47]), 
      .COUT());
endmodule

module FA__4_35(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_39(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_43(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_47(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_51(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_55(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_59(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_63(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_67(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_71(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_75(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_79(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_83(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_87(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_91(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_95(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_99(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_103(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_107(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_111(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_115(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_119(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_123(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(COUT));
endmodule

module FA__4_127(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_131(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_135(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_139(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_143(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_147(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_151(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_155(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_159(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_163(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_167(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_171(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_175(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_179(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_183(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_187(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   AND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(COUT));
   XOR2_X1 i_0_1 (.A(B), .B(A), .Z(SUM));
endmodule

module FA__4_191(A, B, CIN, SUM, COUT);
   input A;
   input B;
   input CIN;
   output SUM;
   output COUT;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(SUM));
endmodule

module CSAlike(result, carry, A, B, C);
   output [63:0]result;
   output [63:0]carry;
   input [63:0]A;
   input [63:0]B;
   input [63:0]C;

   FA__4_35 genblk1_8_fa (.A(A[8]), .B(B[8]), .CIN(), .SUM(), .COUT(carry[9]));
   FA__4_39 genblk1_9_fa (.A(A[9]), .B(B[9]), .CIN(), .SUM(result[9]), .COUT(
      carry[10]));
   FA__4_43 genblk1_10_fa (.A(A[10]), .B(B[10]), .CIN(), .SUM(result[10]), 
      .COUT(carry[11]));
   FA__4_47 genblk1_11_fa (.A(A[11]), .B(B[11]), .CIN(), .SUM(result[11]), 
      .COUT(carry[12]));
   FA__4_51 genblk1_12_fa (.A(A[12]), .B(B[12]), .CIN(), .SUM(result[12]), 
      .COUT(carry[13]));
   FA__4_55 genblk1_13_fa (.A(A[13]), .B(B[13]), .CIN(), .SUM(result[13]), 
      .COUT(carry[14]));
   FA__4_59 genblk1_14_fa (.A(A[14]), .B(B[14]), .CIN(), .SUM(result[14]), 
      .COUT(carry[15]));
   FA__4_63 genblk1_15_fa (.A(A[15]), .B(B[15]), .CIN(), .SUM(result[15]), 
      .COUT(carry[16]));
   FA__4_67 genblk1_16_fa (.A(A[16]), .B(B[16]), .CIN(), .SUM(result[16]), 
      .COUT(carry[17]));
   FA__4_71 genblk1_17_fa (.A(A[17]), .B(B[17]), .CIN(), .SUM(result[17]), 
      .COUT(carry[18]));
   FA__4_75 genblk1_18_fa (.A(A[18]), .B(B[18]), .CIN(), .SUM(result[18]), 
      .COUT(carry[19]));
   FA__4_79 genblk1_19_fa (.A(A[19]), .B(B[19]), .CIN(), .SUM(result[19]), 
      .COUT(carry[20]));
   FA__4_83 genblk1_20_fa (.A(A[20]), .B(B[20]), .CIN(), .SUM(result[20]), 
      .COUT(carry[21]));
   FA__4_87 genblk1_21_fa (.A(A[21]), .B(B[21]), .CIN(), .SUM(result[21]), 
      .COUT(carry[22]));
   FA__4_91 genblk1_22_fa (.A(A[22]), .B(B[22]), .CIN(), .SUM(result[22]), 
      .COUT(carry[23]));
   FA__4_95 genblk1_23_fa (.A(A[23]), .B(B[23]), .CIN(), .SUM(result[23]), 
      .COUT(carry[24]));
   FA__4_99 genblk1_24_fa (.A(A[24]), .B(B[24]), .CIN(), .SUM(result[24]), 
      .COUT(carry[25]));
   FA__4_103 genblk1_25_fa (.A(A[25]), .B(B[25]), .CIN(), .SUM(result[25]), 
      .COUT(carry[26]));
   FA__4_107 genblk1_26_fa (.A(A[26]), .B(B[26]), .CIN(), .SUM(result[26]), 
      .COUT(carry[27]));
   FA__4_111 genblk1_27_fa (.A(A[27]), .B(B[27]), .CIN(), .SUM(result[27]), 
      .COUT(carry[28]));
   FA__4_115 genblk1_28_fa (.A(A[28]), .B(B[28]), .CIN(), .SUM(result[28]), 
      .COUT(carry[29]));
   FA__4_119 genblk1_29_fa (.A(A[29]), .B(B[29]), .CIN(), .SUM(result[29]), 
      .COUT(carry[30]));
   FA__4_123 genblk1_30_fa (.A(A[30]), .B(B[30]), .CIN(), .SUM(result[30]), 
      .COUT(carry[31]));
   FA__4_127 genblk1_31_fa (.A(A[31]), .B(B[31]), .CIN(), .SUM(result[31]), 
      .COUT(carry[32]));
   FA__4_131 genblk1_32_fa (.A(A[32]), .B(B[32]), .CIN(), .SUM(result[32]), 
      .COUT(carry[33]));
   FA__4_135 genblk1_33_fa (.A(A[33]), .B(B[33]), .CIN(), .SUM(result[33]), 
      .COUT(carry[34]));
   FA__4_139 genblk1_34_fa (.A(A[34]), .B(B[34]), .CIN(), .SUM(result[34]), 
      .COUT(carry[35]));
   FA__4_143 genblk1_35_fa (.A(A[35]), .B(B[35]), .CIN(), .SUM(result[35]), 
      .COUT(carry[36]));
   FA__4_147 genblk1_36_fa (.A(A[36]), .B(B[36]), .CIN(), .SUM(result[36]), 
      .COUT(carry[37]));
   FA__4_151 genblk1_37_fa (.A(A[37]), .B(B[37]), .CIN(), .SUM(result[37]), 
      .COUT(carry[38]));
   FA__4_155 genblk1_38_fa (.A(A[38]), .B(B[38]), .CIN(), .SUM(result[38]), 
      .COUT(carry[39]));
   FA__4_159 genblk1_39_fa (.A(A[39]), .B(B[39]), .CIN(), .SUM(result[39]), 
      .COUT(carry[40]));
   FA__4_163 genblk1_40_fa (.A(A[40]), .B(B[40]), .CIN(), .SUM(result[40]), 
      .COUT(carry[41]));
   FA__4_167 genblk1_41_fa (.A(A[41]), .B(B[41]), .CIN(), .SUM(result[41]), 
      .COUT(carry[42]));
   FA__4_171 genblk1_42_fa (.A(A[42]), .B(B[42]), .CIN(), .SUM(result[42]), 
      .COUT(carry[43]));
   FA__4_175 genblk1_43_fa (.A(A[43]), .B(B[43]), .CIN(), .SUM(result[43]), 
      .COUT(carry[44]));
   FA__4_179 genblk1_44_fa (.A(A[44]), .B(B[44]), .CIN(), .SUM(result[44]), 
      .COUT(carry[45]));
   FA__4_183 genblk1_45_fa (.A(A[45]), .B(B[45]), .CIN(), .SUM(result[45]), 
      .COUT(carry[46]));
   FA__4_187 genblk1_46_fa (.A(A[46]), .B(B[46]), .CIN(), .SUM(result[46]), 
      .COUT(carry[47]));
   FA__4_191 genblk1_47_fa (.A(A[47]), .B(B[47]), .CIN(), .SUM(result[47]), 
      .COUT());
endmodule

module addIntermedaiteWires(Res, carry, normalizedWires);
   output [63:0]Res;
   output [63:0]carry;
   input [2047:0]normalizedWires;

   wire [63:0]\intermediateWiresStage1[15] ;
   wire [63:0]\intermediateWiresStage1[14] ;
   wire [63:0]\intermediateWiresStage1[13] ;
   wire [63:0]\intermediateWiresStage1[12] ;
   wire [63:0]\intermediateWiresStage1[11] ;
   wire [63:0]\intermediateWiresStage1[10] ;
   wire [63:0]\intermediateWiresStage1[9] ;
   wire [63:0]\intermediateWiresStage1[8] ;
   wire [63:0]\intermediateWiresStage1[7] ;
   wire [63:0]\intermediateWiresStage1[6] ;
   wire [63:0]\intermediateWiresStage1[5] ;
   wire [63:0]\intermediateWiresStage1[4] ;
   wire [63:0]\intermediateWiresStage1[3] ;
   wire [63:0]\intermediateWiresStage1[2] ;
   wire [63:0]\intermediateWiresStage1[1] ;
   wire [63:0]\intermediateWiresStage1[0] ;
   wire [63:0]\intermediateWiresStage2[9] ;
   wire [63:0]\intermediateWiresStage2[8] ;
   wire [63:0]\intermediateWiresStage2[7] ;
   wire [63:0]\intermediateWiresStage2[6] ;
   wire [63:0]\intermediateWiresStage2[5] ;
   wire [63:0]\intermediateWiresStage2[4] ;
   wire [63:0]\intermediateWiresStage2[3] ;
   wire [63:0]\intermediateWiresStage2[2] ;
   wire [63:0]\intermediateWiresStage2[1] ;
   wire [63:0]\intermediateWiresStage2[0] ;
   wire [63:0]\intermediateWiresStage3[7] ;
   wire [63:0]\intermediateWiresStage3[6] ;
   wire [63:0]\intermediateWiresStage3[5] ;
   wire [63:0]\intermediateWiresStage3[4] ;
   wire [63:0]\intermediateWiresStage3[3] ;
   wire [63:0]\intermediateWiresStage3[2] ;
   wire [63:0]\intermediateWiresStage3[1] ;
   wire [63:0]\intermediateWiresStage3[0] ;
   wire [63:0]\intermediateWiresStage4[5] ;
   wire [63:0]\intermediateWiresStage4[4] ;
   wire [63:0]\intermediateWiresStage4[3] ;
   wire [63:0]\intermediateWiresStage4[2] ;
   wire [63:0]\intermediateWiresStage4[1] ;
   wire [63:0]\intermediateWiresStage4[0] ;
   wire [63:0]\intermediateWiresStage5[3] ;
   wire [63:0]\intermediateWiresStage5[2] ;
   wire [63:0]\intermediateWiresStage5[1] ;
   wire [63:0]\intermediateWiresStage5[0] ;
   wire [63:0]\intermediateWiresStage6[1] ;
   wire [63:0]\intermediateWiresStage6[0] ;
   wire [63:0]\intermediateWiresStage7[1] ;
   wire [63:0]\intermediateWiresStage7[0] ;

   CSAlike__1_1006 genblk2_7_parallelAdderStage1 (.result({uc_0, uc_1, uc_2, 
      uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, 
      uc_14, uc_15, uc_16, uc_17, \intermediateWiresStage1[14] [45], 
      \intermediateWiresStage1[14] [44], \intermediateWiresStage1[14] [43], 
      \intermediateWiresStage1[14] [42], \intermediateWiresStage1[14] [41], 
      \intermediateWiresStage1[14] [40], \intermediateWiresStage1[14] [39], 
      \intermediateWiresStage1[14] [38], \intermediateWiresStage1[14] [37], 
      \intermediateWiresStage1[14] [36], \intermediateWiresStage1[14] [35], 
      \intermediateWiresStage1[14] [34], \intermediateWiresStage1[14] [33], 
      \intermediateWiresStage1[14] [32], \intermediateWiresStage1[14] [31], 
      \intermediateWiresStage1[14] [30], \intermediateWiresStage1[14] [29], 
      \intermediateWiresStage1[14] [28], \intermediateWiresStage1[14] [27], 
      \intermediateWiresStage1[14] [26], \intermediateWiresStage1[14] [25], 
      \intermediateWiresStage1[14] [24], \intermediateWiresStage1[14] [23], 
      \intermediateWiresStage1[14] [22], uc_18, uc_19, uc_20, uc_21, uc_22, 
      uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, uc_32, 
      uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39}), .carry({uc_40, uc_41, 
      uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49, uc_50, uc_51, 
      uc_52, uc_53, uc_54, uc_55, uc_56, \intermediateWiresStage1[15] [46], 
      \intermediateWiresStage1[15] [45], \intermediateWiresStage1[15] [44], 
      \intermediateWiresStage1[15] [43], \intermediateWiresStage1[15] [42], 
      \intermediateWiresStage1[15] [41], \intermediateWiresStage1[15] [40], 
      \intermediateWiresStage1[15] [39], \intermediateWiresStage1[15] [38], 
      \intermediateWiresStage1[15] [37], \intermediateWiresStage1[15] [36], 
      \intermediateWiresStage1[15] [35], \intermediateWiresStage1[15] [34], 
      \intermediateWiresStage1[15] [33], \intermediateWiresStage1[15] [32], 
      \intermediateWiresStage1[15] [31], \intermediateWiresStage1[15] [30], 
      \intermediateWiresStage1[15] [29], \intermediateWiresStage1[15] [28], 
      \intermediateWiresStage1[15] [27], \intermediateWiresStage1[15] [26], 
      \intermediateWiresStage1[15] [25], \intermediateWiresStage1[15] [24], 
      \intermediateWiresStage1[15] [23], uc_57, uc_58, uc_59, uc_60, uc_61, 
      uc_62, uc_63, uc_64, uc_65, uc_66, uc_67, uc_68, uc_69, uc_70, uc_71, 
      uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, uc_79}), .A({1'b0, uc_80, 
      uc_81, uc_82, uc_83, uc_84, uc_85, uc_86, uc_87, uc_88, uc_89, uc_90, 
      uc_91, uc_92, uc_93, uc_94, uc_95, uc_96, uc_97, normalizedWires[1388], 
      normalizedWires[1387], normalizedWires[1386], normalizedWires[1385], 
      normalizedWires[1384], normalizedWires[1383], normalizedWires[1382], 
      normalizedWires[1381], normalizedWires[1380], normalizedWires[1379], 
      normalizedWires[1378], normalizedWires[1377], normalizedWires[1376], 
      normalizedWires[1375], normalizedWires[1374], normalizedWires[1373], 
      normalizedWires[1372], normalizedWires[1371], normalizedWires[1370], 
      normalizedWires[1369], normalizedWires[1368], normalizedWires[1367], 
      normalizedWires[1366], uc_98, uc_99, uc_100, uc_101, uc_102, uc_103, 
      uc_104, uc_105, uc_106, uc_107, uc_108, uc_109, uc_110, uc_111, uc_112, 
      uc_113, uc_114, uc_115, uc_116, uc_117, uc_118, uc_119}), .B({1'b0, uc_120, 
      uc_121, uc_122, uc_123, uc_124, uc_125, uc_126, uc_127, uc_128, uc_129, 
      uc_130, uc_131, uc_132, uc_133, uc_134, uc_135, uc_136, 
      normalizedWires[1453], normalizedWires[1452], normalizedWires[1451], 
      normalizedWires[1450], normalizedWires[1449], normalizedWires[1448], 
      normalizedWires[1447], normalizedWires[1446], normalizedWires[1445], 
      normalizedWires[1444], normalizedWires[1443], normalizedWires[1442], 
      normalizedWires[1441], normalizedWires[1440], normalizedWires[1439], 
      normalizedWires[1438], normalizedWires[1437], normalizedWires[1436], 
      normalizedWires[1435], normalizedWires[1434], normalizedWires[1433], 
      normalizedWires[1432], normalizedWires[1431], normalizedWires[1430], 
      uc_137, uc_138, uc_139, uc_140, uc_141, uc_142, uc_143, uc_144, uc_145, 
      uc_146, uc_147, uc_148, uc_149, uc_150, uc_151, uc_152, uc_153, uc_154, 
      uc_155, uc_156, uc_157, uc_158}), .C({1'b0, uc_159, uc_160, uc_161, uc_162, 
      uc_163, uc_164, uc_165, uc_166, uc_167, uc_168, uc_169, uc_170, uc_171, 
      uc_172, uc_173, uc_174, uc_175, normalizedWires[1517], 
      normalizedWires[1516], normalizedWires[1515], normalizedWires[1514], 
      normalizedWires[1513], normalizedWires[1512], normalizedWires[1511], 
      normalizedWires[1510], normalizedWires[1509], normalizedWires[1508], 
      normalizedWires[1507], normalizedWires[1506], normalizedWires[1505], 
      normalizedWires[1504], normalizedWires[1503], normalizedWires[1502], 
      normalizedWires[1501], normalizedWires[1500], normalizedWires[1499], 
      normalizedWires[1498], normalizedWires[1497], normalizedWires[1496], 
      normalizedWires[1495], uc_176, uc_177, uc_178, uc_179, uc_180, uc_181, 
      uc_182, uc_183, uc_184, uc_185, uc_186, uc_187, uc_188, uc_189, uc_190, 
      uc_191, uc_192, uc_193, uc_194, uc_195, uc_196, uc_197, uc_198}));
   CSAlike__1_1259 genblk2_6_parallelAdderStage1 (.result({uc_199, uc_200, 
      uc_201, uc_202, uc_203, uc_204, uc_205, uc_206, uc_207, uc_208, uc_209, 
      uc_210, uc_211, uc_212, uc_213, uc_214, uc_215, uc_216, uc_217, uc_218, 
      uc_219, \intermediateWiresStage1[12] [42], 
      \intermediateWiresStage1[12] [41], \intermediateWiresStage1[12] [40], 
      \intermediateWiresStage1[12] [39], \intermediateWiresStage1[12] [38], 
      \intermediateWiresStage1[12] [37], \intermediateWiresStage1[12] [36], 
      \intermediateWiresStage1[12] [35], \intermediateWiresStage1[12] [34], 
      \intermediateWiresStage1[12] [33], \intermediateWiresStage1[12] [32], 
      \intermediateWiresStage1[12] [31], \intermediateWiresStage1[12] [30], 
      \intermediateWiresStage1[12] [29], \intermediateWiresStage1[12] [28], 
      \intermediateWiresStage1[12] [27], \intermediateWiresStage1[12] [26], 
      \intermediateWiresStage1[12] [25], \intermediateWiresStage1[12] [24], 
      \intermediateWiresStage1[12] [23], \intermediateWiresStage1[12] [22], 
      \intermediateWiresStage1[12] [21], \intermediateWiresStage1[12] [20], 
      \intermediateWiresStage1[12] [19], uc_220, uc_221, uc_222, uc_223, uc_224, 
      uc_225, uc_226, uc_227, uc_228, uc_229, uc_230, uc_231, uc_232, uc_233, 
      uc_234, uc_235, uc_236, uc_237, uc_238}), .carry({uc_239, uc_240, uc_241, 
      uc_242, uc_243, uc_244, uc_245, uc_246, uc_247, uc_248, uc_249, uc_250, 
      uc_251, uc_252, uc_253, uc_254, uc_255, uc_256, uc_257, uc_258, 
      \intermediateWiresStage1[13] [43], \intermediateWiresStage1[13] [42], 
      \intermediateWiresStage1[13] [41], \intermediateWiresStage1[13] [40], 
      \intermediateWiresStage1[13] [39], \intermediateWiresStage1[13] [38], 
      \intermediateWiresStage1[13] [37], \intermediateWiresStage1[13] [36], 
      \intermediateWiresStage1[13] [35], \intermediateWiresStage1[13] [34], 
      \intermediateWiresStage1[13] [33], \intermediateWiresStage1[13] [32], 
      \intermediateWiresStage1[13] [31], \intermediateWiresStage1[13] [30], 
      \intermediateWiresStage1[13] [29], \intermediateWiresStage1[13] [28], 
      \intermediateWiresStage1[13] [27], \intermediateWiresStage1[13] [26], 
      \intermediateWiresStage1[13] [25], \intermediateWiresStage1[13] [24], 
      \intermediateWiresStage1[13] [23], \intermediateWiresStage1[13] [22], 
      \intermediateWiresStage1[13] [21], \intermediateWiresStage1[13] [20], 
      uc_259, uc_260, uc_261, uc_262, uc_263, uc_264, uc_265, uc_266, uc_267, 
      uc_268, uc_269, uc_270, uc_271, uc_272, uc_273, uc_274, uc_275, uc_276, 
      uc_277, uc_278}), .A({1'b0, uc_279, uc_280, uc_281, uc_282, uc_283, uc_284, 
      uc_285, uc_286, uc_287, uc_288, uc_289, uc_290, uc_291, uc_292, uc_293, 
      uc_294, uc_295, uc_296, uc_297, uc_298, uc_299, normalizedWires[1193], 
      normalizedWires[1192], normalizedWires[1191], normalizedWires[1190], 
      normalizedWires[1189], normalizedWires[1188], normalizedWires[1187], 
      normalizedWires[1186], normalizedWires[1185], normalizedWires[1184], 
      normalizedWires[1183], normalizedWires[1182], normalizedWires[1181], 
      normalizedWires[1180], normalizedWires[1179], normalizedWires[1178], 
      normalizedWires[1177], normalizedWires[1176], normalizedWires[1175], 
      normalizedWires[1174], normalizedWires[1173], normalizedWires[1172], 
      normalizedWires[1171], uc_300, uc_301, uc_302, uc_303, uc_304, uc_305, 
      uc_306, uc_307, uc_308, uc_309, uc_310, uc_311, uc_312, uc_313, uc_314, 
      uc_315, uc_316, uc_317, uc_318}), .B({1'b0, uc_319, uc_320, uc_321, uc_322, 
      uc_323, uc_324, uc_325, uc_326, uc_327, uc_328, uc_329, uc_330, uc_331, 
      uc_332, uc_333, uc_334, uc_335, uc_336, uc_337, uc_338, 
      normalizedWires[1258], normalizedWires[1257], normalizedWires[1256], 
      normalizedWires[1255], normalizedWires[1254], normalizedWires[1253], 
      normalizedWires[1252], normalizedWires[1251], normalizedWires[1250], 
      normalizedWires[1249], normalizedWires[1248], normalizedWires[1247], 
      normalizedWires[1246], normalizedWires[1245], normalizedWires[1244], 
      normalizedWires[1243], normalizedWires[1242], normalizedWires[1241], 
      normalizedWires[1240], normalizedWires[1239], normalizedWires[1238], 
      normalizedWires[1237], normalizedWires[1236], normalizedWires[1235], 
      uc_339, uc_340, uc_341, uc_342, uc_343, uc_344, uc_345, uc_346, uc_347, 
      uc_348, uc_349, uc_350, uc_351, uc_352, uc_353, uc_354, uc_355, uc_356, 
      uc_357}), .C({1'b0, uc_358, uc_359, uc_360, uc_361, uc_362, uc_363, uc_364, 
      uc_365, uc_366, uc_367, uc_368, uc_369, uc_370, uc_371, uc_372, uc_373, 
      uc_374, uc_375, uc_376, uc_377, normalizedWires[1322], 
      normalizedWires[1321], normalizedWires[1320], normalizedWires[1319], 
      normalizedWires[1318], normalizedWires[1317], normalizedWires[1316], 
      normalizedWires[1315], normalizedWires[1314], normalizedWires[1313], 
      normalizedWires[1312], normalizedWires[1311], normalizedWires[1310], 
      normalizedWires[1309], normalizedWires[1308], normalizedWires[1307], 
      normalizedWires[1306], normalizedWires[1305], normalizedWires[1304], 
      normalizedWires[1303], normalizedWires[1302], normalizedWires[1301], 
      normalizedWires[1300], uc_378, uc_379, uc_380, uc_381, uc_382, uc_383, 
      uc_384, uc_385, uc_386, uc_387, uc_388, uc_389, uc_390, uc_391, uc_392, 
      uc_393, uc_394, uc_395, uc_396, uc_397}));
   CSAlike__1_1512 genblk2_5_parallelAdderStage1 (.result({uc_398, uc_399, 
      uc_400, uc_401, uc_402, uc_403, uc_404, uc_405, uc_406, uc_407, uc_408, 
      uc_409, uc_410, uc_411, uc_412, uc_413, uc_414, uc_415, uc_416, uc_417, 
      uc_418, uc_419, uc_420, uc_421, \intermediateWiresStage1[10] [39], 
      \intermediateWiresStage1[10] [38], \intermediateWiresStage1[10] [37], 
      \intermediateWiresStage1[10] [36], \intermediateWiresStage1[10] [35], 
      \intermediateWiresStage1[10] [34], \intermediateWiresStage1[10] [33], 
      \intermediateWiresStage1[10] [32], \intermediateWiresStage1[10] [31], 
      \intermediateWiresStage1[10] [30], \intermediateWiresStage1[10] [29], 
      \intermediateWiresStage1[10] [28], \intermediateWiresStage1[10] [27], 
      \intermediateWiresStage1[10] [26], \intermediateWiresStage1[10] [25], 
      \intermediateWiresStage1[10] [24], \intermediateWiresStage1[10] [23], 
      \intermediateWiresStage1[10] [22], \intermediateWiresStage1[10] [21], 
      \intermediateWiresStage1[10] [20], \intermediateWiresStage1[10] [19], 
      \intermediateWiresStage1[10] [18], \intermediateWiresStage1[10] [17], 
      \intermediateWiresStage1[10] [16], uc_422, uc_423, uc_424, uc_425, uc_426, 
      uc_427, uc_428, uc_429, uc_430, uc_431, uc_432, uc_433, uc_434, uc_435, 
      uc_436, uc_437}), .carry({uc_438, uc_439, uc_440, uc_441, uc_442, uc_443, 
      uc_444, uc_445, uc_446, uc_447, uc_448, uc_449, uc_450, uc_451, uc_452, 
      uc_453, uc_454, uc_455, uc_456, uc_457, uc_458, uc_459, uc_460, 
      \intermediateWiresStage1[11] [40], \intermediateWiresStage1[11] [39], 
      \intermediateWiresStage1[11] [38], \intermediateWiresStage1[11] [37], 
      \intermediateWiresStage1[11] [36], \intermediateWiresStage1[11] [35], 
      \intermediateWiresStage1[11] [34], \intermediateWiresStage1[11] [33], 
      \intermediateWiresStage1[11] [32], \intermediateWiresStage1[11] [31], 
      \intermediateWiresStage1[11] [30], \intermediateWiresStage1[11] [29], 
      \intermediateWiresStage1[11] [28], \intermediateWiresStage1[11] [27], 
      \intermediateWiresStage1[11] [26], \intermediateWiresStage1[11] [25], 
      \intermediateWiresStage1[11] [24], \intermediateWiresStage1[11] [23], 
      \intermediateWiresStage1[11] [22], \intermediateWiresStage1[11] [21], 
      \intermediateWiresStage1[11] [20], \intermediateWiresStage1[11] [19], 
      \intermediateWiresStage1[11] [18], \intermediateWiresStage1[11] [17], 
      uc_461, uc_462, uc_463, uc_464, uc_465, uc_466, uc_467, uc_468, uc_469, 
      uc_470, uc_471, uc_472, uc_473, uc_474, uc_475, uc_476, uc_477}), .A({1'b0, 
      uc_478, uc_479, uc_480, uc_481, uc_482, uc_483, uc_484, uc_485, uc_486, 
      uc_487, uc_488, uc_489, uc_490, uc_491, uc_492, uc_493, uc_494, uc_495, 
      uc_496, uc_497, uc_498, uc_499, uc_500, uc_501, normalizedWires[998], 
      normalizedWires[997], normalizedWires[996], normalizedWires[995], 
      normalizedWires[994], normalizedWires[993], normalizedWires[992], 
      normalizedWires[991], normalizedWires[990], normalizedWires[989], 
      normalizedWires[988], normalizedWires[987], normalizedWires[986], 
      normalizedWires[985], normalizedWires[984], normalizedWires[983], 
      normalizedWires[982], normalizedWires[981], normalizedWires[980], 
      normalizedWires[979], normalizedWires[978], normalizedWires[977], 
      normalizedWires[976], uc_502, uc_503, uc_504, uc_505, uc_506, uc_507, 
      uc_508, uc_509, uc_510, uc_511, uc_512, uc_513, uc_514, uc_515, uc_516, 
      uc_517}), .B({1'b0, uc_518, uc_519, uc_520, uc_521, uc_522, uc_523, uc_524, 
      uc_525, uc_526, uc_527, uc_528, uc_529, uc_530, uc_531, uc_532, uc_533, 
      uc_534, uc_535, uc_536, uc_537, uc_538, uc_539, uc_540, 
      normalizedWires[1063], normalizedWires[1062], normalizedWires[1061], 
      normalizedWires[1060], normalizedWires[1059], normalizedWires[1058], 
      normalizedWires[1057], normalizedWires[1056], normalizedWires[1055], 
      normalizedWires[1054], normalizedWires[1053], normalizedWires[1052], 
      normalizedWires[1051], normalizedWires[1050], normalizedWires[1049], 
      normalizedWires[1048], normalizedWires[1047], normalizedWires[1046], 
      normalizedWires[1045], normalizedWires[1044], normalizedWires[1043], 
      normalizedWires[1042], normalizedWires[1041], normalizedWires[1040], 
      uc_541, uc_542, uc_543, uc_544, uc_545, uc_546, uc_547, uc_548, uc_549, 
      uc_550, uc_551, uc_552, uc_553, uc_554, uc_555, uc_556}), .C({1'b0, uc_557, 
      uc_558, uc_559, uc_560, uc_561, uc_562, uc_563, uc_564, uc_565, uc_566, 
      uc_567, uc_568, uc_569, uc_570, uc_571, uc_572, uc_573, uc_574, uc_575, 
      uc_576, uc_577, uc_578, uc_579, normalizedWires[1127], 
      normalizedWires[1126], normalizedWires[1125], normalizedWires[1124], 
      normalizedWires[1123], normalizedWires[1122], normalizedWires[1121], 
      normalizedWires[1120], normalizedWires[1119], normalizedWires[1118], 
      normalizedWires[1117], normalizedWires[1116], normalizedWires[1115], 
      normalizedWires[1114], normalizedWires[1113], normalizedWires[1112], 
      normalizedWires[1111], normalizedWires[1110], normalizedWires[1109], 
      normalizedWires[1108], normalizedWires[1107], normalizedWires[1106], 
      normalizedWires[1105], uc_580, uc_581, uc_582, uc_583, uc_584, uc_585, 
      uc_586, uc_587, uc_588, uc_589, uc_590, uc_591, uc_592, uc_593, uc_594, 
      uc_595, uc_596}));
   CSAlike__1_1765 genblk2_4_parallelAdderStage1 (.result({uc_597, uc_598, 
      uc_599, uc_600, uc_601, uc_602, uc_603, uc_604, uc_605, uc_606, uc_607, 
      uc_608, uc_609, uc_610, uc_611, uc_612, uc_613, uc_614, uc_615, uc_616, 
      uc_617, uc_618, uc_619, uc_620, uc_621, uc_622, uc_623, 
      \intermediateWiresStage1[8] [36], \intermediateWiresStage1[8] [35], 
      \intermediateWiresStage1[8] [34], \intermediateWiresStage1[8] [33], 
      \intermediateWiresStage1[8] [32], \intermediateWiresStage1[8] [31], 
      \intermediateWiresStage1[8] [30], \intermediateWiresStage1[8] [29], 
      \intermediateWiresStage1[8] [28], \intermediateWiresStage1[8] [27], 
      \intermediateWiresStage1[8] [26], \intermediateWiresStage1[8] [25], 
      \intermediateWiresStage1[8] [24], \intermediateWiresStage1[8] [23], 
      \intermediateWiresStage1[8] [22], \intermediateWiresStage1[8] [21], 
      \intermediateWiresStage1[8] [20], \intermediateWiresStage1[8] [19], 
      \intermediateWiresStage1[8] [18], \intermediateWiresStage1[8] [17], 
      \intermediateWiresStage1[8] [16], \intermediateWiresStage1[8] [15], 
      \intermediateWiresStage1[8] [14], \intermediateWiresStage1[8] [13], uc_624, 
      uc_625, uc_626, uc_627, uc_628, uc_629, uc_630, uc_631, uc_632, uc_633, 
      uc_634, uc_635, uc_636}), .carry({uc_637, uc_638, uc_639, uc_640, uc_641, 
      uc_642, uc_643, uc_644, uc_645, uc_646, uc_647, uc_648, uc_649, uc_650, 
      uc_651, uc_652, uc_653, uc_654, uc_655, uc_656, uc_657, uc_658, uc_659, 
      uc_660, uc_661, uc_662, \intermediateWiresStage1[9] [37], 
      \intermediateWiresStage1[9] [36], \intermediateWiresStage1[9] [35], 
      \intermediateWiresStage1[9] [34], \intermediateWiresStage1[9] [33], 
      \intermediateWiresStage1[9] [32], \intermediateWiresStage1[9] [31], 
      \intermediateWiresStage1[9] [30], \intermediateWiresStage1[9] [29], 
      \intermediateWiresStage1[9] [28], \intermediateWiresStage1[9] [27], 
      \intermediateWiresStage1[9] [26], \intermediateWiresStage1[9] [25], 
      \intermediateWiresStage1[9] [24], \intermediateWiresStage1[9] [23], 
      \intermediateWiresStage1[9] [22], \intermediateWiresStage1[9] [21], 
      \intermediateWiresStage1[9] [20], \intermediateWiresStage1[9] [19], 
      \intermediateWiresStage1[9] [18], \intermediateWiresStage1[9] [17], 
      \intermediateWiresStage1[9] [16], \intermediateWiresStage1[9] [15], 
      \intermediateWiresStage1[9] [14], uc_663, uc_664, uc_665, uc_666, uc_667, 
      uc_668, uc_669, uc_670, uc_671, uc_672, uc_673, uc_674, uc_675, uc_676}), 
      .A({1'b0, uc_677, uc_678, uc_679, uc_680, uc_681, uc_682, uc_683, uc_684, 
      uc_685, uc_686, uc_687, uc_688, uc_689, uc_690, uc_691, uc_692, uc_693, 
      uc_694, uc_695, uc_696, uc_697, uc_698, uc_699, uc_700, uc_701, uc_702, 
      uc_703, normalizedWires[803], normalizedWires[802], normalizedWires[801], 
      normalizedWires[800], normalizedWires[799], normalizedWires[798], 
      normalizedWires[797], normalizedWires[796], normalizedWires[795], 
      normalizedWires[794], normalizedWires[793], normalizedWires[792], 
      normalizedWires[791], normalizedWires[790], normalizedWires[789], 
      normalizedWires[788], normalizedWires[787], normalizedWires[786], 
      normalizedWires[785], normalizedWires[784], normalizedWires[783], 
      normalizedWires[782], normalizedWires[781], uc_704, uc_705, uc_706, uc_707, 
      uc_708, uc_709, uc_710, uc_711, uc_712, uc_713, uc_714, uc_715, uc_716}), 
      .B({1'b0, uc_717, uc_718, uc_719, uc_720, uc_721, uc_722, uc_723, uc_724, 
      uc_725, uc_726, uc_727, uc_728, uc_729, uc_730, uc_731, uc_732, uc_733, 
      uc_734, uc_735, uc_736, uc_737, uc_738, uc_739, uc_740, uc_741, uc_742, 
      normalizedWires[868], normalizedWires[867], normalizedWires[866], 
      normalizedWires[865], normalizedWires[864], normalizedWires[863], 
      normalizedWires[862], normalizedWires[861], normalizedWires[860], 
      normalizedWires[859], normalizedWires[858], normalizedWires[857], 
      normalizedWires[856], normalizedWires[855], normalizedWires[854], 
      normalizedWires[853], normalizedWires[852], normalizedWires[851], 
      normalizedWires[850], normalizedWires[849], normalizedWires[848], 
      normalizedWires[847], normalizedWires[846], normalizedWires[845], uc_743, 
      uc_744, uc_745, uc_746, uc_747, uc_748, uc_749, uc_750, uc_751, uc_752, 
      uc_753, uc_754, uc_755}), .C({1'b0, uc_756, uc_757, uc_758, uc_759, uc_760, 
      uc_761, uc_762, uc_763, uc_764, uc_765, uc_766, uc_767, uc_768, uc_769, 
      uc_770, uc_771, uc_772, uc_773, uc_774, uc_775, uc_776, uc_777, uc_778, 
      uc_779, uc_780, uc_781, normalizedWires[932], normalizedWires[931], 
      normalizedWires[930], normalizedWires[929], normalizedWires[928], 
      normalizedWires[927], normalizedWires[926], normalizedWires[925], 
      normalizedWires[924], normalizedWires[923], normalizedWires[922], 
      normalizedWires[921], normalizedWires[920], normalizedWires[919], 
      normalizedWires[918], normalizedWires[917], normalizedWires[916], 
      normalizedWires[915], normalizedWires[914], normalizedWires[913], 
      normalizedWires[912], normalizedWires[911], normalizedWires[910], uc_782, 
      uc_783, uc_784, uc_785, uc_786, uc_787, uc_788, uc_789, uc_790, uc_791, 
      uc_792, uc_793, uc_794, uc_795}));
   CSAlike__1_2018 genblk2_3_parallelAdderStage1 (.result({uc_796, uc_797, 
      uc_798, uc_799, uc_800, uc_801, uc_802, uc_803, uc_804, uc_805, uc_806, 
      uc_807, uc_808, uc_809, uc_810, uc_811, uc_812, uc_813, uc_814, uc_815, 
      uc_816, uc_817, uc_818, uc_819, uc_820, uc_821, uc_822, uc_823, uc_824, 
      uc_825, \intermediateWiresStage1[6] [33], \intermediateWiresStage1[6] [32], 
      \intermediateWiresStage1[6] [31], \intermediateWiresStage1[6] [30], 
      \intermediateWiresStage1[6] [29], \intermediateWiresStage1[6] [28], 
      \intermediateWiresStage1[6] [27], \intermediateWiresStage1[6] [26], 
      \intermediateWiresStage1[6] [25], \intermediateWiresStage1[6] [24], 
      \intermediateWiresStage1[6] [23], \intermediateWiresStage1[6] [22], 
      \intermediateWiresStage1[6] [21], \intermediateWiresStage1[6] [20], 
      \intermediateWiresStage1[6] [19], \intermediateWiresStage1[6] [18], 
      \intermediateWiresStage1[6] [17], \intermediateWiresStage1[6] [16], 
      \intermediateWiresStage1[6] [15], \intermediateWiresStage1[6] [14], 
      \intermediateWiresStage1[6] [13], \intermediateWiresStage1[6] [12], 
      \intermediateWiresStage1[6] [11], \intermediateWiresStage1[6] [10], uc_826, 
      uc_827, uc_828, uc_829, uc_830, uc_831, uc_832, uc_833, uc_834, uc_835}), 
      .carry({uc_836, uc_837, uc_838, uc_839, uc_840, uc_841, uc_842, uc_843, 
      uc_844, uc_845, uc_846, uc_847, uc_848, uc_849, uc_850, uc_851, uc_852, 
      uc_853, uc_854, uc_855, uc_856, uc_857, uc_858, uc_859, uc_860, uc_861, 
      uc_862, uc_863, uc_864, \intermediateWiresStage1[7] [34], 
      \intermediateWiresStage1[7] [33], \intermediateWiresStage1[7] [32], 
      \intermediateWiresStage1[7] [31], \intermediateWiresStage1[7] [30], 
      \intermediateWiresStage1[7] [29], \intermediateWiresStage1[7] [28], 
      \intermediateWiresStage1[7] [27], \intermediateWiresStage1[7] [26], 
      \intermediateWiresStage1[7] [25], \intermediateWiresStage1[7] [24], 
      \intermediateWiresStage1[7] [23], \intermediateWiresStage1[7] [22], 
      \intermediateWiresStage1[7] [21], \intermediateWiresStage1[7] [20], 
      \intermediateWiresStage1[7] [19], \intermediateWiresStage1[7] [18], 
      \intermediateWiresStage1[7] [17], \intermediateWiresStage1[7] [16], 
      \intermediateWiresStage1[7] [15], \intermediateWiresStage1[7] [14], 
      \intermediateWiresStage1[7] [13], \intermediateWiresStage1[7] [12], 
      \intermediateWiresStage1[7] [11], uc_865, uc_866, uc_867, uc_868, uc_869, 
      uc_870, uc_871, uc_872, uc_873, uc_874, uc_875}), .A({1'b0, uc_876, uc_877, 
      uc_878, uc_879, uc_880, uc_881, uc_882, uc_883, uc_884, uc_885, uc_886, 
      uc_887, uc_888, uc_889, uc_890, uc_891, uc_892, uc_893, uc_894, uc_895, 
      uc_896, uc_897, uc_898, uc_899, uc_900, uc_901, uc_902, uc_903, uc_904, 
      uc_905, normalizedWires[608], normalizedWires[607], normalizedWires[606], 
      normalizedWires[605], normalizedWires[604], normalizedWires[603], 
      normalizedWires[602], normalizedWires[601], normalizedWires[600], 
      normalizedWires[599], normalizedWires[598], normalizedWires[597], 
      normalizedWires[596], normalizedWires[595], normalizedWires[594], 
      normalizedWires[593], normalizedWires[592], normalizedWires[591], 
      normalizedWires[590], normalizedWires[589], normalizedWires[588], 
      normalizedWires[587], normalizedWires[586], uc_906, uc_907, uc_908, uc_909, 
      uc_910, uc_911, uc_912, uc_913, uc_914, uc_915}), .B({1'b0, uc_916, uc_917, 
      uc_918, uc_919, uc_920, uc_921, uc_922, uc_923, uc_924, uc_925, uc_926, 
      uc_927, uc_928, uc_929, uc_930, uc_931, uc_932, uc_933, uc_934, uc_935, 
      uc_936, uc_937, uc_938, uc_939, uc_940, uc_941, uc_942, uc_943, uc_944, 
      normalizedWires[673], normalizedWires[672], normalizedWires[671], 
      normalizedWires[670], normalizedWires[669], normalizedWires[668], 
      normalizedWires[667], normalizedWires[666], normalizedWires[665], 
      normalizedWires[664], normalizedWires[663], normalizedWires[662], 
      normalizedWires[661], normalizedWires[660], normalizedWires[659], 
      normalizedWires[658], normalizedWires[657], normalizedWires[656], 
      normalizedWires[655], normalizedWires[654], normalizedWires[653], 
      normalizedWires[652], normalizedWires[651], normalizedWires[650], uc_945, 
      uc_946, uc_947, uc_948, uc_949, uc_950, uc_951, uc_952, uc_953, uc_954}), 
      .C({1'b0, uc_955, uc_956, uc_957, uc_958, uc_959, uc_960, uc_961, uc_962, 
      uc_963, uc_964, uc_965, uc_966, uc_967, uc_968, uc_969, uc_970, uc_971, 
      uc_972, uc_973, uc_974, uc_975, uc_976, uc_977, uc_978, uc_979, uc_980, 
      uc_981, uc_982, uc_983, normalizedWires[737], normalizedWires[736], 
      normalizedWires[735], normalizedWires[734], normalizedWires[733], 
      normalizedWires[732], normalizedWires[731], normalizedWires[730], 
      normalizedWires[729], normalizedWires[728], normalizedWires[727], 
      normalizedWires[726], normalizedWires[725], normalizedWires[724], 
      normalizedWires[723], normalizedWires[722], normalizedWires[721], 
      normalizedWires[720], normalizedWires[719], normalizedWires[718], 
      normalizedWires[717], normalizedWires[716], normalizedWires[715], uc_984, 
      uc_985, uc_986, uc_987, uc_988, uc_989, uc_990, uc_991, uc_992, uc_993, 
      uc_994}));
   CSAlike__1_2271 genblk2_2_parallelAdderStage1 (.result({uc_995, uc_996, 
      uc_997, uc_998, uc_999, uc_1000, uc_1001, uc_1002, uc_1003, uc_1004, 
      uc_1005, uc_1006, uc_1007, uc_1008, uc_1009, uc_1010, uc_1011, uc_1012, 
      uc_1013, uc_1014, uc_1015, uc_1016, uc_1017, uc_1018, uc_1019, uc_1020, 
      uc_1021, uc_1022, uc_1023, uc_1024, uc_1025, uc_1026, uc_1027, 
      \intermediateWiresStage1[4] [30], \intermediateWiresStage1[4] [29], 
      \intermediateWiresStage1[4] [28], \intermediateWiresStage1[4] [27], 
      \intermediateWiresStage1[4] [26], \intermediateWiresStage1[4] [25], 
      \intermediateWiresStage1[4] [24], \intermediateWiresStage1[4] [23], 
      \intermediateWiresStage1[4] [22], \intermediateWiresStage1[4] [21], 
      \intermediateWiresStage1[4] [20], \intermediateWiresStage1[4] [19], 
      \intermediateWiresStage1[4] [18], \intermediateWiresStage1[4] [17], 
      \intermediateWiresStage1[4] [16], \intermediateWiresStage1[4] [15], 
      \intermediateWiresStage1[4] [14], \intermediateWiresStage1[4] [13], 
      \intermediateWiresStage1[4] [12], \intermediateWiresStage1[4] [11], 
      \intermediateWiresStage1[4] [10], \intermediateWiresStage1[4] [9], 
      \intermediateWiresStage1[4] [8], \intermediateWiresStage1[4] [7], uc_1028, 
      uc_1029, uc_1030, uc_1031, uc_1032, uc_1033, uc_1034}), .carry({uc_1035, 
      uc_1036, uc_1037, uc_1038, uc_1039, uc_1040, uc_1041, uc_1042, uc_1043, 
      uc_1044, uc_1045, uc_1046, uc_1047, uc_1048, uc_1049, uc_1050, uc_1051, 
      uc_1052, uc_1053, uc_1054, uc_1055, uc_1056, uc_1057, uc_1058, uc_1059, 
      uc_1060, uc_1061, uc_1062, uc_1063, uc_1064, uc_1065, uc_1066, 
      \intermediateWiresStage1[5] [31], \intermediateWiresStage1[5] [30], 
      \intermediateWiresStage1[5] [29], \intermediateWiresStage1[5] [28], 
      \intermediateWiresStage1[5] [27], \intermediateWiresStage1[5] [26], 
      \intermediateWiresStage1[5] [25], \intermediateWiresStage1[5] [24], 
      \intermediateWiresStage1[5] [23], \intermediateWiresStage1[5] [22], 
      \intermediateWiresStage1[5] [21], \intermediateWiresStage1[5] [20], 
      \intermediateWiresStage1[5] [19], \intermediateWiresStage1[5] [18], 
      \intermediateWiresStage1[5] [17], \intermediateWiresStage1[5] [16], 
      \intermediateWiresStage1[5] [15], \intermediateWiresStage1[5] [14], 
      \intermediateWiresStage1[5] [13], \intermediateWiresStage1[5] [12], 
      \intermediateWiresStage1[5] [11], \intermediateWiresStage1[5] [10], 
      \intermediateWiresStage1[5] [9], \intermediateWiresStage1[5] [8], uc_1067, 
      uc_1068, uc_1069, uc_1070, uc_1071, uc_1072, uc_1073, uc_1074}), .A({1'b0, 
      uc_1075, uc_1076, uc_1077, uc_1078, uc_1079, uc_1080, uc_1081, uc_1082, 
      uc_1083, uc_1084, uc_1085, uc_1086, uc_1087, uc_1088, uc_1089, uc_1090, 
      uc_1091, uc_1092, uc_1093, uc_1094, uc_1095, uc_1096, uc_1097, uc_1098, 
      uc_1099, uc_1100, uc_1101, uc_1102, uc_1103, uc_1104, uc_1105, uc_1106, 
      uc_1107, normalizedWires[413], normalizedWires[412], normalizedWires[411], 
      normalizedWires[410], normalizedWires[409], normalizedWires[408], 
      normalizedWires[407], normalizedWires[406], normalizedWires[405], 
      normalizedWires[404], normalizedWires[403], normalizedWires[402], 
      normalizedWires[401], normalizedWires[400], normalizedWires[399], 
      normalizedWires[398], normalizedWires[397], normalizedWires[396], 
      normalizedWires[395], normalizedWires[394], normalizedWires[393], 
      normalizedWires[392], normalizedWires[391], uc_1108, uc_1109, uc_1110, 
      uc_1111, uc_1112, uc_1113, uc_1114}), .B({1'b0, uc_1115, uc_1116, uc_1117, 
      uc_1118, uc_1119, uc_1120, uc_1121, uc_1122, uc_1123, uc_1124, uc_1125, 
      uc_1126, uc_1127, uc_1128, uc_1129, uc_1130, uc_1131, uc_1132, uc_1133, 
      uc_1134, uc_1135, uc_1136, uc_1137, uc_1138, uc_1139, uc_1140, uc_1141, 
      uc_1142, uc_1143, uc_1144, uc_1145, uc_1146, normalizedWires[478], 
      normalizedWires[477], normalizedWires[476], normalizedWires[475], 
      normalizedWires[474], normalizedWires[473], normalizedWires[472], 
      normalizedWires[471], normalizedWires[470], normalizedWires[469], 
      normalizedWires[468], normalizedWires[467], normalizedWires[466], 
      normalizedWires[465], normalizedWires[464], normalizedWires[463], 
      normalizedWires[462], normalizedWires[461], normalizedWires[460], 
      normalizedWires[459], normalizedWires[458], normalizedWires[457], 
      normalizedWires[456], normalizedWires[455], uc_1147, uc_1148, uc_1149, 
      uc_1150, uc_1151, uc_1152, uc_1153}), .C({1'b0, uc_1154, uc_1155, uc_1156, 
      uc_1157, uc_1158, uc_1159, uc_1160, uc_1161, uc_1162, uc_1163, uc_1164, 
      uc_1165, uc_1166, uc_1167, uc_1168, uc_1169, uc_1170, uc_1171, uc_1172, 
      uc_1173, uc_1174, uc_1175, uc_1176, uc_1177, uc_1178, uc_1179, uc_1180, 
      uc_1181, uc_1182, uc_1183, uc_1184, uc_1185, normalizedWires[542], 
      normalizedWires[541], normalizedWires[540], normalizedWires[539], 
      normalizedWires[538], normalizedWires[537], normalizedWires[536], 
      normalizedWires[535], normalizedWires[534], normalizedWires[533], 
      normalizedWires[532], normalizedWires[531], normalizedWires[530], 
      normalizedWires[529], normalizedWires[528], normalizedWires[527], 
      normalizedWires[526], normalizedWires[525], normalizedWires[524], 
      normalizedWires[523], normalizedWires[522], normalizedWires[521], 
      normalizedWires[520], uc_1186, uc_1187, uc_1188, uc_1189, uc_1190, uc_1191, 
      uc_1192, uc_1193}));
   CSAlike__1_2524 genblk2_1_parallelAdderStage1 (.result({uc_1194, uc_1195, 
      uc_1196, uc_1197, uc_1198, uc_1199, uc_1200, uc_1201, uc_1202, uc_1203, 
      uc_1204, uc_1205, uc_1206, uc_1207, uc_1208, uc_1209, uc_1210, uc_1211, 
      uc_1212, uc_1213, uc_1214, uc_1215, uc_1216, uc_1217, uc_1218, uc_1219, 
      uc_1220, uc_1221, uc_1222, uc_1223, uc_1224, uc_1225, uc_1226, uc_1227, 
      uc_1228, uc_1229, \intermediateWiresStage1[2] [27], 
      \intermediateWiresStage1[2] [26], \intermediateWiresStage1[2] [25], 
      \intermediateWiresStage1[2] [24], \intermediateWiresStage1[2] [23], 
      \intermediateWiresStage1[2] [22], \intermediateWiresStage1[2] [21], 
      \intermediateWiresStage1[2] [20], \intermediateWiresStage1[2] [19], 
      \intermediateWiresStage1[2] [18], \intermediateWiresStage1[2] [17], 
      \intermediateWiresStage1[2] [16], \intermediateWiresStage1[2] [15], 
      \intermediateWiresStage1[2] [14], \intermediateWiresStage1[2] [13], 
      \intermediateWiresStage1[2] [12], \intermediateWiresStage1[2] [11], 
      \intermediateWiresStage1[2] [10], \intermediateWiresStage1[2] [9], 
      \intermediateWiresStage1[2] [8], \intermediateWiresStage1[2] [7], 
      \intermediateWiresStage1[2] [6], \intermediateWiresStage1[2] [5], 
      \intermediateWiresStage1[2] [4], uc_1230, uc_1231, uc_1232, uc_1233}), 
      .carry({uc_1234, uc_1235, uc_1236, uc_1237, uc_1238, uc_1239, uc_1240, 
      uc_1241, uc_1242, uc_1243, uc_1244, uc_1245, uc_1246, uc_1247, uc_1248, 
      uc_1249, uc_1250, uc_1251, uc_1252, uc_1253, uc_1254, uc_1255, uc_1256, 
      uc_1257, uc_1258, uc_1259, uc_1260, uc_1261, uc_1262, uc_1263, uc_1264, 
      uc_1265, uc_1266, uc_1267, uc_1268, \intermediateWiresStage1[3] [28], 
      \intermediateWiresStage1[3] [27], \intermediateWiresStage1[3] [26], 
      \intermediateWiresStage1[3] [25], \intermediateWiresStage1[3] [24], 
      \intermediateWiresStage1[3] [23], \intermediateWiresStage1[3] [22], 
      \intermediateWiresStage1[3] [21], \intermediateWiresStage1[3] [20], 
      \intermediateWiresStage1[3] [19], \intermediateWiresStage1[3] [18], 
      \intermediateWiresStage1[3] [17], \intermediateWiresStage1[3] [16], 
      \intermediateWiresStage1[3] [15], \intermediateWiresStage1[3] [14], 
      \intermediateWiresStage1[3] [13], \intermediateWiresStage1[3] [12], 
      \intermediateWiresStage1[3] [11], \intermediateWiresStage1[3] [10], 
      \intermediateWiresStage1[3] [9], \intermediateWiresStage1[3] [8], 
      \intermediateWiresStage1[3] [7], \intermediateWiresStage1[3] [6], 
      \intermediateWiresStage1[3] [5], uc_1269, uc_1270, uc_1271, uc_1272, 
      uc_1273}), .A({1'b0, uc_1274, uc_1275, uc_1276, uc_1277, uc_1278, uc_1279, 
      uc_1280, uc_1281, uc_1282, uc_1283, uc_1284, uc_1285, uc_1286, uc_1287, 
      uc_1288, uc_1289, uc_1290, uc_1291, uc_1292, uc_1293, uc_1294, uc_1295, 
      uc_1296, uc_1297, uc_1298, uc_1299, uc_1300, uc_1301, uc_1302, uc_1303, 
      uc_1304, uc_1305, uc_1306, uc_1307, uc_1308, uc_1309, normalizedWires[218], 
      normalizedWires[217], normalizedWires[216], normalizedWires[215], 
      normalizedWires[214], normalizedWires[213], normalizedWires[212], 
      normalizedWires[211], normalizedWires[210], normalizedWires[209], 
      normalizedWires[208], normalizedWires[207], normalizedWires[206], 
      normalizedWires[205], normalizedWires[204], normalizedWires[203], 
      normalizedWires[202], normalizedWires[201], normalizedWires[200], 
      normalizedWires[199], normalizedWires[198], normalizedWires[197], 
      normalizedWires[196], uc_1310, uc_1311, uc_1312, uc_1313}), .B({1'b0, 
      uc_1314, uc_1315, uc_1316, uc_1317, uc_1318, uc_1319, uc_1320, uc_1321, 
      uc_1322, uc_1323, uc_1324, uc_1325, uc_1326, uc_1327, uc_1328, uc_1329, 
      uc_1330, uc_1331, uc_1332, uc_1333, uc_1334, uc_1335, uc_1336, uc_1337, 
      uc_1338, uc_1339, uc_1340, uc_1341, uc_1342, uc_1343, uc_1344, uc_1345, 
      uc_1346, uc_1347, uc_1348, normalizedWires[283], normalizedWires[282], 
      normalizedWires[281], normalizedWires[280], normalizedWires[279], 
      normalizedWires[278], normalizedWires[277], normalizedWires[276], 
      normalizedWires[275], normalizedWires[274], normalizedWires[273], 
      normalizedWires[272], normalizedWires[271], normalizedWires[270], 
      normalizedWires[269], normalizedWires[268], normalizedWires[267], 
      normalizedWires[266], normalizedWires[265], normalizedWires[264], 
      normalizedWires[263], normalizedWires[262], normalizedWires[261], 
      normalizedWires[260], uc_1349, uc_1350, uc_1351, uc_1352}), .C({1'b0, 
      uc_1353, uc_1354, uc_1355, uc_1356, uc_1357, uc_1358, uc_1359, uc_1360, 
      uc_1361, uc_1362, uc_1363, uc_1364, uc_1365, uc_1366, uc_1367, uc_1368, 
      uc_1369, uc_1370, uc_1371, uc_1372, uc_1373, uc_1374, uc_1375, uc_1376, 
      uc_1377, uc_1378, uc_1379, uc_1380, uc_1381, uc_1382, uc_1383, uc_1384, 
      uc_1385, uc_1386, uc_1387, normalizedWires[347], normalizedWires[346], 
      normalizedWires[345], normalizedWires[344], normalizedWires[343], 
      normalizedWires[342], normalizedWires[341], normalizedWires[340], 
      normalizedWires[339], normalizedWires[338], normalizedWires[337], 
      normalizedWires[336], normalizedWires[335], normalizedWires[334], 
      normalizedWires[333], normalizedWires[332], normalizedWires[331], 
      normalizedWires[330], normalizedWires[329], normalizedWires[328], 
      normalizedWires[327], normalizedWires[326], normalizedWires[325], uc_1388, 
      uc_1389, uc_1390, uc_1391, uc_1392}));
   CSAlike__0_108 genblk2_0_parallelAdderStage1 (.result({uc_1393, uc_1394, 
      uc_1395, uc_1396, uc_1397, uc_1398, uc_1399, uc_1400, uc_1401, uc_1402, 
      uc_1403, uc_1404, uc_1405, uc_1406, uc_1407, uc_1408, uc_1409, uc_1410, 
      uc_1411, uc_1412, uc_1413, uc_1414, uc_1415, uc_1416, uc_1417, uc_1418, 
      uc_1419, uc_1420, uc_1421, uc_1422, uc_1423, uc_1424, uc_1425, uc_1426, 
      uc_1427, uc_1428, uc_1429, uc_1430, uc_1431, 
      \intermediateWiresStage1[0] [24], \intermediateWiresStage1[0] [23], 
      \intermediateWiresStage1[0] [22], \intermediateWiresStage1[0] [21], 
      \intermediateWiresStage1[0] [20], \intermediateWiresStage1[0] [19], 
      \intermediateWiresStage1[0] [18], \intermediateWiresStage1[0] [17], 
      \intermediateWiresStage1[0] [16], \intermediateWiresStage1[0] [15], 
      \intermediateWiresStage1[0] [14], \intermediateWiresStage1[0] [13], 
      \intermediateWiresStage1[0] [12], \intermediateWiresStage1[0] [11], 
      \intermediateWiresStage1[0] [10], \intermediateWiresStage1[0] [9], 
      \intermediateWiresStage1[0] [8], \intermediateWiresStage1[0] [7], 
      \intermediateWiresStage1[0] [6], \intermediateWiresStage1[0] [5], 
      \intermediateWiresStage1[0] [4], \intermediateWiresStage1[0] [3], 
      \intermediateWiresStage1[0] [2], uc_1432, uc_1433}), .carry({uc_1434, 
      uc_1435, uc_1436, uc_1437, uc_1438, uc_1439, uc_1440, uc_1441, uc_1442, 
      uc_1443, uc_1444, uc_1445, uc_1446, uc_1447, uc_1448, uc_1449, uc_1450, 
      uc_1451, uc_1452, uc_1453, uc_1454, uc_1455, uc_1456, uc_1457, uc_1458, 
      uc_1459, uc_1460, uc_1461, uc_1462, uc_1463, uc_1464, uc_1465, uc_1466, 
      uc_1467, uc_1468, uc_1469, uc_1470, uc_1471, 
      \intermediateWiresStage1[1] [25], \intermediateWiresStage1[1] [24], 
      \intermediateWiresStage1[1] [23], \intermediateWiresStage1[1] [22], 
      \intermediateWiresStage1[1] [21], \intermediateWiresStage1[1] [20], 
      \intermediateWiresStage1[1] [19], \intermediateWiresStage1[1] [18], 
      \intermediateWiresStage1[1] [17], \intermediateWiresStage1[1] [16], 
      \intermediateWiresStage1[1] [15], \intermediateWiresStage1[1] [14], 
      \intermediateWiresStage1[1] [13], \intermediateWiresStage1[1] [12], 
      \intermediateWiresStage1[1] [11], \intermediateWiresStage1[1] [10], 
      \intermediateWiresStage1[1] [9], \intermediateWiresStage1[1] [8], 
      \intermediateWiresStage1[1] [7], \intermediateWiresStage1[1] [6], 
      \intermediateWiresStage1[1] [5], \intermediateWiresStage1[1] [4], 
      \intermediateWiresStage1[1] [3], \intermediateWiresStage1[1] [2], uc_1472, 
      uc_1473}), .A({1'b0, uc_1474, uc_1475, uc_1476, uc_1477, uc_1478, uc_1479, 
      uc_1480, uc_1481, uc_1482, uc_1483, uc_1484, uc_1485, uc_1486, uc_1487, 
      uc_1488, uc_1489, uc_1490, uc_1491, uc_1492, uc_1493, uc_1494, uc_1495, 
      uc_1496, uc_1497, uc_1498, uc_1499, uc_1500, uc_1501, uc_1502, uc_1503, 
      uc_1504, uc_1505, uc_1506, uc_1507, uc_1508, uc_1509, uc_1510, uc_1511, 
      uc_1512, normalizedWires[23], normalizedWires[22], normalizedWires[21], 
      normalizedWires[20], normalizedWires[19], normalizedWires[18], 
      normalizedWires[17], normalizedWires[16], normalizedWires[15], 
      normalizedWires[14], normalizedWires[13], normalizedWires[12], 
      normalizedWires[11], normalizedWires[10], normalizedWires[9], 
      normalizedWires[8], normalizedWires[7], normalizedWires[6], 
      normalizedWires[5], normalizedWires[4], normalizedWires[3], 
      normalizedWires[2], normalizedWires[1], uc_1513}), .B({1'b0, uc_1514, 
      uc_1515, uc_1516, uc_1517, uc_1518, uc_1519, uc_1520, uc_1521, uc_1522, 
      uc_1523, uc_1524, uc_1525, uc_1526, uc_1527, uc_1528, uc_1529, uc_1530, 
      uc_1531, uc_1532, uc_1533, uc_1534, uc_1535, uc_1536, uc_1537, uc_1538, 
      uc_1539, uc_1540, uc_1541, uc_1542, uc_1543, uc_1544, uc_1545, uc_1546, 
      uc_1547, uc_1548, uc_1549, uc_1550, uc_1551, normalizedWires[88], 
      normalizedWires[87], normalizedWires[86], normalizedWires[85], 
      normalizedWires[84], normalizedWires[83], normalizedWires[82], 
      normalizedWires[81], normalizedWires[80], normalizedWires[79], 
      normalizedWires[78], normalizedWires[77], normalizedWires[76], 
      normalizedWires[75], normalizedWires[74], normalizedWires[73], 
      normalizedWires[72], normalizedWires[71], normalizedWires[70], 
      normalizedWires[69], normalizedWires[68], normalizedWires[67], 
      normalizedWires[66], normalizedWires[65], uc_1552}), .C({1'b0, uc_1553, 
      uc_1554, uc_1555, uc_1556, uc_1557, uc_1558, uc_1559, uc_1560, uc_1561, 
      uc_1562, uc_1563, uc_1564, uc_1565, uc_1566, uc_1567, uc_1568, uc_1569, 
      uc_1570, uc_1571, uc_1572, uc_1573, uc_1574, uc_1575, uc_1576, uc_1577, 
      uc_1578, uc_1579, uc_1580, uc_1581, uc_1582, uc_1583, uc_1584, uc_1585, 
      uc_1586, uc_1587, uc_1588, uc_1589, uc_1590, normalizedWires[152], 
      normalizedWires[151], normalizedWires[150], normalizedWires[149], 
      normalizedWires[148], normalizedWires[147], normalizedWires[146], 
      normalizedWires[145], normalizedWires[144], normalizedWires[143], 
      normalizedWires[142], normalizedWires[141], normalizedWires[140], 
      normalizedWires[139], normalizedWires[138], normalizedWires[137], 
      normalizedWires[136], normalizedWires[135], normalizedWires[134], 
      normalizedWires[133], normalizedWires[132], normalizedWires[131], 
      normalizedWires[130], uc_1591, uc_1592}));
   CSAlike__2_1006 genblk3_4_parallelAdderStage2 (.result({uc_1593, uc_1594, 
      uc_1595, uc_1596, uc_1597, uc_1598, uc_1599, uc_1600, uc_1601, uc_1602, 
      uc_1603, uc_1604, uc_1605, uc_1606, uc_1607, uc_1608, uc_1609, uc_1610, 
      uc_1611, uc_1612, \intermediateWiresStage2[8] [43], 
      \intermediateWiresStage2[8] [42], \intermediateWiresStage2[8] [41], 
      \intermediateWiresStage2[8] [40], \intermediateWiresStage2[8] [39], 
      \intermediateWiresStage2[8] [38], \intermediateWiresStage2[8] [37], 
      \intermediateWiresStage2[8] [36], \intermediateWiresStage2[8] [35], 
      \intermediateWiresStage2[8] [34], \intermediateWiresStage2[8] [33], 
      \intermediateWiresStage2[8] [32], \intermediateWiresStage2[8] [31], 
      \intermediateWiresStage2[8] [30], \intermediateWiresStage2[8] [29], 
      \intermediateWiresStage2[8] [28], \intermediateWiresStage2[8] [27], 
      \intermediateWiresStage2[8] [26], \intermediateWiresStage2[8] [25], 
      \intermediateWiresStage2[8] [24], \intermediateWiresStage2[8] [23], 
      \intermediateWiresStage2[8] [22], \intermediateWiresStage2[8] [21], 
      \intermediateWiresStage2[8] [20], uc_1613, uc_1614, uc_1615, uc_1616, 
      uc_1617, uc_1618, uc_1619, uc_1620, uc_1621, uc_1622, uc_1623, uc_1624, 
      uc_1625, uc_1626, uc_1627, uc_1628, uc_1629, uc_1630, uc_1631, uc_1632}), 
      .carry({uc_1633, uc_1634, uc_1635, uc_1636, uc_1637, uc_1638, uc_1639, 
      uc_1640, uc_1641, uc_1642, uc_1643, uc_1644, uc_1645, uc_1646, uc_1647, 
      uc_1648, uc_1649, uc_1650, uc_1651, \intermediateWiresStage2[9] [44], 
      \intermediateWiresStage2[9] [43], \intermediateWiresStage2[9] [42], 
      \intermediateWiresStage2[9] [41], \intermediateWiresStage2[9] [40], 
      \intermediateWiresStage2[9] [39], \intermediateWiresStage2[9] [38], 
      \intermediateWiresStage2[9] [37], \intermediateWiresStage2[9] [36], 
      \intermediateWiresStage2[9] [35], \intermediateWiresStage2[9] [34], 
      \intermediateWiresStage2[9] [33], \intermediateWiresStage2[9] [32], 
      \intermediateWiresStage2[9] [31], \intermediateWiresStage2[9] [30], 
      \intermediateWiresStage2[9] [29], \intermediateWiresStage2[9] [28], 
      \intermediateWiresStage2[9] [27], \intermediateWiresStage2[9] [26], 
      \intermediateWiresStage2[9] [25], \intermediateWiresStage2[9] [24], 
      \intermediateWiresStage2[9] [23], \intermediateWiresStage2[9] [22], 
      \intermediateWiresStage2[9] [21], uc_1652, uc_1653, uc_1654, uc_1655, 
      uc_1656, uc_1657, uc_1658, uc_1659, uc_1660, uc_1661, uc_1662, uc_1663, 
      uc_1664, uc_1665, uc_1666, uc_1667, uc_1668, uc_1669, uc_1670, uc_1671, 
      uc_1672}), .A({1'b0, uc_1673, uc_1674, uc_1675, uc_1676, uc_1677, uc_1678, 
      uc_1679, uc_1680, uc_1681, uc_1682, uc_1683, uc_1684, uc_1685, 1'b0, 1'b0, 
      uc_1686, uc_1687, uc_1688, uc_1689, normalizedWires[1323], 
      \intermediateWiresStage1[12] [42], \intermediateWiresStage1[12] [41], 
      \intermediateWiresStage1[12] [40], \intermediateWiresStage1[12] [39], 
      \intermediateWiresStage1[12] [38], \intermediateWiresStage1[12] [37], 
      \intermediateWiresStage1[12] [36], \intermediateWiresStage1[12] [35], 
      \intermediateWiresStage1[12] [34], \intermediateWiresStage1[12] [33], 
      \intermediateWiresStage1[12] [32], \intermediateWiresStage1[12] [31], 
      \intermediateWiresStage1[12] [30], \intermediateWiresStage1[12] [29], 
      \intermediateWiresStage1[12] [28], \intermediateWiresStage1[12] [27], 
      \intermediateWiresStage1[12] [26], \intermediateWiresStage1[12] [25], 
      \intermediateWiresStage1[12] [24], \intermediateWiresStage1[12] [23], 
      \intermediateWiresStage1[12] [22], \intermediateWiresStage1[12] [21], 
      \intermediateWiresStage1[12] [20], uc_1690, uc_1691, uc_1692, uc_1693, 
      uc_1694, uc_1695, uc_1696, uc_1697, uc_1698, uc_1699, uc_1700, uc_1701, 
      uc_1702, uc_1703, uc_1704, uc_1705, uc_1706, uc_1707, uc_1708, uc_1709}), 
      .B({1'b0, uc_1710, uc_1711, uc_1712, uc_1713, uc_1714, uc_1715, uc_1716, 
      uc_1717, uc_1718, uc_1719, uc_1720, uc_1721, 1'b0, 1'b0, 1'b0, uc_1722, 
      uc_1723, uc_1724, uc_1725, \intermediateWiresStage1[13] [43], 
      \intermediateWiresStage1[13] [42], \intermediateWiresStage1[13] [41], 
      \intermediateWiresStage1[13] [40], \intermediateWiresStage1[13] [39], 
      \intermediateWiresStage1[13] [38], \intermediateWiresStage1[13] [37], 
      \intermediateWiresStage1[13] [36], \intermediateWiresStage1[13] [35], 
      \intermediateWiresStage1[13] [34], \intermediateWiresStage1[13] [33], 
      \intermediateWiresStage1[13] [32], \intermediateWiresStage1[13] [31], 
      \intermediateWiresStage1[13] [30], \intermediateWiresStage1[13] [29], 
      \intermediateWiresStage1[13] [28], \intermediateWiresStage1[13] [27], 
      \intermediateWiresStage1[13] [26], \intermediateWiresStage1[13] [25], 
      \intermediateWiresStage1[13] [24], \intermediateWiresStage1[13] [23], 
      \intermediateWiresStage1[13] [22], \intermediateWiresStage1[13] [21], 
      \intermediateWiresStage1[13] [20], uc_1726, uc_1727, uc_1728, uc_1729, 
      uc_1730, uc_1731, uc_1732, uc_1733, uc_1734, uc_1735, uc_1736, uc_1737, 
      uc_1738, uc_1739, uc_1740, uc_1741, uc_1742, uc_1743, uc_1744, uc_1745}), 
      .C({1'b0, uc_1746, uc_1747, uc_1748, uc_1749, uc_1750, uc_1751, uc_1752, 
      uc_1753, uc_1754, uc_1755, uc_1756, uc_1757, 1'b0, 1'b0, 1'b0, uc_1758, 
      uc_1759, uc_1760, uc_1761, \intermediateWiresStage1[14] [43], 
      \intermediateWiresStage1[14] [42], \intermediateWiresStage1[14] [41], 
      \intermediateWiresStage1[14] [40], \intermediateWiresStage1[14] [39], 
      \intermediateWiresStage1[14] [38], \intermediateWiresStage1[14] [37], 
      \intermediateWiresStage1[14] [36], \intermediateWiresStage1[14] [35], 
      \intermediateWiresStage1[14] [34], \intermediateWiresStage1[14] [33], 
      \intermediateWiresStage1[14] [32], \intermediateWiresStage1[14] [31], 
      \intermediateWiresStage1[14] [30], \intermediateWiresStage1[14] [29], 
      \intermediateWiresStage1[14] [28], \intermediateWiresStage1[14] [27], 
      \intermediateWiresStage1[14] [26], \intermediateWiresStage1[14] [25], 
      \intermediateWiresStage1[14] [24], \intermediateWiresStage1[14] [23], 
      \intermediateWiresStage1[14] [22], normalizedWires[1365], uc_1762, uc_1763, 
      uc_1764, uc_1765, uc_1766, uc_1767, uc_1768, uc_1769, uc_1770, uc_1771, 
      uc_1772, uc_1773, uc_1774, uc_1775, uc_1776, uc_1777, uc_1778, uc_1779, 
      uc_1780, uc_1781, uc_1782}));
   CSAlike__2_1259 genblk3_3_parallelAdderStage2 (.result({uc_1783, uc_1784, 
      uc_1785, uc_1786, uc_1787, uc_1788, uc_1789, uc_1790, uc_1791, uc_1792, 
      uc_1793, uc_1794, uc_1795, uc_1796, uc_1797, uc_1798, uc_1799, uc_1800, 
      uc_1801, uc_1802, uc_1803, uc_1804, uc_1805, 
      \intermediateWiresStage2[6] [40], \intermediateWiresStage2[6] [39], 
      \intermediateWiresStage2[6] [38], \intermediateWiresStage2[6] [37], 
      \intermediateWiresStage2[6] [36], \intermediateWiresStage2[6] [35], 
      \intermediateWiresStage2[6] [34], \intermediateWiresStage2[6] [33], 
      \intermediateWiresStage2[6] [32], \intermediateWiresStage2[6] [31], 
      \intermediateWiresStage2[6] [30], \intermediateWiresStage2[6] [29], 
      \intermediateWiresStage2[6] [28], \intermediateWiresStage2[6] [27], 
      \intermediateWiresStage2[6] [26], \intermediateWiresStage2[6] [25], 
      \intermediateWiresStage2[6] [24], \intermediateWiresStage2[6] [23], 
      \intermediateWiresStage2[6] [22], \intermediateWiresStage2[6] [21], 
      \intermediateWiresStage2[6] [20], \intermediateWiresStage2[6] [19], 
      \intermediateWiresStage2[6] [18], \intermediateWiresStage2[6] [17], 
      \intermediateWiresStage2[6] [16], \intermediateWiresStage2[6] [15], 
      uc_1806, uc_1807, uc_1808, uc_1809, uc_1810, uc_1811, uc_1812, uc_1813, 
      uc_1814, uc_1815, uc_1816, uc_1817, uc_1818, uc_1819, uc_1820}), .carry({
      uc_1821, uc_1822, uc_1823, uc_1824, uc_1825, uc_1826, uc_1827, uc_1828, 
      uc_1829, uc_1830, uc_1831, uc_1832, uc_1833, uc_1834, uc_1835, uc_1836, 
      uc_1837, uc_1838, uc_1839, uc_1840, uc_1841, uc_1842, 
      \intermediateWiresStage2[7] [41], \intermediateWiresStage2[7] [40], 
      \intermediateWiresStage2[7] [39], \intermediateWiresStage2[7] [38], 
      \intermediateWiresStage2[7] [37], \intermediateWiresStage2[7] [36], 
      \intermediateWiresStage2[7] [35], \intermediateWiresStage2[7] [34], 
      \intermediateWiresStage2[7] [33], \intermediateWiresStage2[7] [32], 
      \intermediateWiresStage2[7] [31], \intermediateWiresStage2[7] [30], 
      \intermediateWiresStage2[7] [29], \intermediateWiresStage2[7] [28], 
      \intermediateWiresStage2[7] [27], \intermediateWiresStage2[7] [26], 
      \intermediateWiresStage2[7] [25], \intermediateWiresStage2[7] [24], 
      \intermediateWiresStage2[7] [23], \intermediateWiresStage2[7] [22], 
      \intermediateWiresStage2[7] [21], \intermediateWiresStage2[7] [20], 
      \intermediateWiresStage2[7] [19], \intermediateWiresStage2[7] [18], 
      \intermediateWiresStage2[7] [17], \intermediateWiresStage2[7] [16], 
      uc_1843, uc_1844, uc_1845, uc_1846, uc_1847, uc_1848, uc_1849, uc_1850, 
      uc_1851, uc_1852, uc_1853, uc_1854, uc_1855, uc_1856, uc_1857, uc_1858}), 
      .A({1'b0, uc_1859, uc_1860, uc_1861, uc_1862, uc_1863, uc_1864, uc_1865, 
      uc_1866, uc_1867, uc_1868, uc_1869, uc_1870, uc_1871, uc_1872, uc_1873, 
      uc_1874, uc_1875, uc_1876, uc_1877, uc_1878, uc_1879, uc_1880, uc_1881, 
      uc_1882, uc_1883, \intermediateWiresStage1[9] [37], 
      \intermediateWiresStage1[9] [36], \intermediateWiresStage1[9] [35], 
      \intermediateWiresStage1[9] [34], \intermediateWiresStage1[9] [33], 
      \intermediateWiresStage1[9] [32], \intermediateWiresStage1[9] [31], 
      \intermediateWiresStage1[9] [30], \intermediateWiresStage1[9] [29], 
      \intermediateWiresStage1[9] [28], \intermediateWiresStage1[9] [27], 
      \intermediateWiresStage1[9] [26], \intermediateWiresStage1[9] [25], 
      \intermediateWiresStage1[9] [24], \intermediateWiresStage1[9] [23], 
      \intermediateWiresStage1[9] [22], \intermediateWiresStage1[9] [21], 
      \intermediateWiresStage1[9] [20], \intermediateWiresStage1[9] [19], 
      \intermediateWiresStage1[9] [18], \intermediateWiresStage1[9] [17], 
      \intermediateWiresStage1[9] [16], \intermediateWiresStage1[9] [15], 
      uc_1884, uc_1885, uc_1886, uc_1887, uc_1888, uc_1889, uc_1890, uc_1891, 
      uc_1892, uc_1893, uc_1894, uc_1895, uc_1896, uc_1897, uc_1898}), .B({1'b0, 
      uc_1899, uc_1900, uc_1901, uc_1902, uc_1903, uc_1904, uc_1905, uc_1906, 
      uc_1907, uc_1908, uc_1909, uc_1910, uc_1911, uc_1912, uc_1913, uc_1914, 
      uc_1915, uc_1916, uc_1917, uc_1918, uc_1919, uc_1920, 
      normalizedWires[1128], \intermediateWiresStage1[10] [39], 
      \intermediateWiresStage1[10] [38], \intermediateWiresStage1[10] [37], 
      \intermediateWiresStage1[10] [36], \intermediateWiresStage1[10] [35], 
      \intermediateWiresStage1[10] [34], \intermediateWiresStage1[10] [33], 
      \intermediateWiresStage1[10] [32], \intermediateWiresStage1[10] [31], 
      \intermediateWiresStage1[10] [30], \intermediateWiresStage1[10] [29], 
      \intermediateWiresStage1[10] [28], \intermediateWiresStage1[10] [27], 
      \intermediateWiresStage1[10] [26], \intermediateWiresStage1[10] [25], 
      \intermediateWiresStage1[10] [24], \intermediateWiresStage1[10] [23], 
      \intermediateWiresStage1[10] [22], \intermediateWiresStage1[10] [21], 
      \intermediateWiresStage1[10] [20], \intermediateWiresStage1[10] [19], 
      \intermediateWiresStage1[10] [18], \intermediateWiresStage1[10] [17], 
      \intermediateWiresStage1[10] [16], normalizedWires[975], uc_1921, uc_1922, 
      uc_1923, uc_1924, uc_1925, uc_1926, uc_1927, uc_1928, uc_1929, uc_1930, 
      uc_1931, uc_1932, uc_1933, uc_1934, uc_1935}), .C({1'b0, uc_1936, uc_1937, 
      uc_1938, uc_1939, uc_1940, uc_1941, uc_1942, uc_1943, uc_1944, uc_1945, 
      uc_1946, uc_1947, uc_1948, uc_1949, uc_1950, uc_1951, uc_1952, uc_1953, 
      uc_1954, uc_1955, uc_1956, uc_1957, \intermediateWiresStage1[11] [40], 
      \intermediateWiresStage1[11] [39], \intermediateWiresStage1[11] [38], 
      \intermediateWiresStage1[11] [37], \intermediateWiresStage1[11] [36], 
      \intermediateWiresStage1[11] [35], \intermediateWiresStage1[11] [34], 
      \intermediateWiresStage1[11] [33], \intermediateWiresStage1[11] [32], 
      \intermediateWiresStage1[11] [31], \intermediateWiresStage1[11] [30], 
      \intermediateWiresStage1[11] [29], \intermediateWiresStage1[11] [28], 
      \intermediateWiresStage1[11] [27], \intermediateWiresStage1[11] [26], 
      \intermediateWiresStage1[11] [25], \intermediateWiresStage1[11] [24], 
      \intermediateWiresStage1[11] [23], \intermediateWiresStage1[11] [22], 
      \intermediateWiresStage1[11] [21], \intermediateWiresStage1[11] [20], 
      \intermediateWiresStage1[11] [19], \intermediateWiresStage1[11] [18], 
      \intermediateWiresStage1[11] [17], uc_1958, uc_1959, uc_1960, uc_1961, 
      uc_1962, uc_1963, uc_1964, uc_1965, uc_1966, uc_1967, uc_1968, uc_1969, 
      uc_1970, uc_1971, uc_1972, uc_1973, uc_1974}));
   CSAlike__2_1512 genblk3_2_parallelAdderStage2 (.result({uc_1975, uc_1976, 
      uc_1977, uc_1978, uc_1979, uc_1980, uc_1981, uc_1982, uc_1983, uc_1984, 
      uc_1985, uc_1986, uc_1987, uc_1988, uc_1989, uc_1990, uc_1991, uc_1992, 
      uc_1993, uc_1994, uc_1995, uc_1996, uc_1997, uc_1998, uc_1999, uc_2000, 
      uc_2001, uc_2002, uc_2003, \intermediateWiresStage2[4] [34], 
      \intermediateWiresStage2[4] [33], \intermediateWiresStage2[4] [32], 
      \intermediateWiresStage2[4] [31], \intermediateWiresStage2[4] [30], 
      \intermediateWiresStage2[4] [29], \intermediateWiresStage2[4] [28], 
      \intermediateWiresStage2[4] [27], \intermediateWiresStage2[4] [26], 
      \intermediateWiresStage2[4] [25], \intermediateWiresStage2[4] [24], 
      \intermediateWiresStage2[4] [23], \intermediateWiresStage2[4] [22], 
      \intermediateWiresStage2[4] [21], \intermediateWiresStage2[4] [20], 
      \intermediateWiresStage2[4] [19], \intermediateWiresStage2[4] [18], 
      \intermediateWiresStage2[4] [17], \intermediateWiresStage2[4] [16], 
      \intermediateWiresStage2[4] [15], \intermediateWiresStage2[4] [14], 
      \intermediateWiresStage2[4] [13], \intermediateWiresStage2[4] [12], 
      \intermediateWiresStage2[4] [11], uc_2004, uc_2005, uc_2006, uc_2007, 
      uc_2008, uc_2009, uc_2010, uc_2011, uc_2012, uc_2013, uc_2014}), .carry({
      uc_2015, uc_2016, uc_2017, uc_2018, uc_2019, uc_2020, uc_2021, uc_2022, 
      uc_2023, uc_2024, uc_2025, uc_2026, uc_2027, uc_2028, uc_2029, uc_2030, 
      uc_2031, uc_2032, uc_2033, uc_2034, uc_2035, uc_2036, uc_2037, uc_2038, 
      uc_2039, uc_2040, uc_2041, uc_2042, \intermediateWiresStage2[5] [35], 
      \intermediateWiresStage2[5] [34], \intermediateWiresStage2[5] [33], 
      \intermediateWiresStage2[5] [32], \intermediateWiresStage2[5] [31], 
      \intermediateWiresStage2[5] [30], \intermediateWiresStage2[5] [29], 
      \intermediateWiresStage2[5] [28], \intermediateWiresStage2[5] [27], 
      \intermediateWiresStage2[5] [26], \intermediateWiresStage2[5] [25], 
      \intermediateWiresStage2[5] [24], \intermediateWiresStage2[5] [23], 
      \intermediateWiresStage2[5] [22], \intermediateWiresStage2[5] [21], 
      \intermediateWiresStage2[5] [20], \intermediateWiresStage2[5] [19], 
      \intermediateWiresStage2[5] [18], \intermediateWiresStage2[5] [17], 
      \intermediateWiresStage2[5] [16], \intermediateWiresStage2[5] [15], 
      \intermediateWiresStage2[5] [14], \intermediateWiresStage2[5] [13], 
      \intermediateWiresStage2[5] [12], uc_2043, uc_2044, uc_2045, uc_2046, 
      uc_2047, uc_2048, uc_2049, uc_2050, uc_2051, uc_2052, uc_2053, uc_2054}), 
      .A({1'b0, uc_2055, uc_2056, uc_2057, uc_2058, uc_2059, uc_2060, uc_2061, 
      uc_2062, uc_2063, uc_2064, uc_2065, uc_2066, uc_2067, uc_2068, uc_2069, 
      uc_2070, uc_2071, uc_2072, uc_2073, uc_2074, uc_2075, uc_2076, uc_2077, 
      uc_2078, uc_2079, uc_2080, uc_2081, uc_2082, normalizedWires[738], 
      \intermediateWiresStage1[6] [33], \intermediateWiresStage1[6] [32], 
      \intermediateWiresStage1[6] [31], \intermediateWiresStage1[6] [30], 
      \intermediateWiresStage1[6] [29], \intermediateWiresStage1[6] [28], 
      \intermediateWiresStage1[6] [27], \intermediateWiresStage1[6] [26], 
      \intermediateWiresStage1[6] [25], \intermediateWiresStage1[6] [24], 
      \intermediateWiresStage1[6] [23], \intermediateWiresStage1[6] [22], 
      \intermediateWiresStage1[6] [21], \intermediateWiresStage1[6] [20], 
      \intermediateWiresStage1[6] [19], \intermediateWiresStage1[6] [18], 
      \intermediateWiresStage1[6] [17], \intermediateWiresStage1[6] [16], 
      \intermediateWiresStage1[6] [15], \intermediateWiresStage1[6] [14], 
      \intermediateWiresStage1[6] [13], \intermediateWiresStage1[6] [12], 
      \intermediateWiresStage1[6] [11], uc_2083, uc_2084, uc_2085, uc_2086, 
      uc_2087, uc_2088, uc_2089, uc_2090, uc_2091, uc_2092, uc_2093}), .B({1'b0, 
      uc_2094, uc_2095, uc_2096, uc_2097, uc_2098, uc_2099, uc_2100, uc_2101, 
      uc_2102, uc_2103, uc_2104, uc_2105, uc_2106, uc_2107, uc_2108, uc_2109, 
      uc_2110, uc_2111, uc_2112, uc_2113, uc_2114, uc_2115, uc_2116, uc_2117, 
      uc_2118, uc_2119, uc_2120, uc_2121, \intermediateWiresStage1[7] [34], 
      \intermediateWiresStage1[7] [33], \intermediateWiresStage1[7] [32], 
      \intermediateWiresStage1[7] [31], \intermediateWiresStage1[7] [30], 
      \intermediateWiresStage1[7] [29], \intermediateWiresStage1[7] [28], 
      \intermediateWiresStage1[7] [27], \intermediateWiresStage1[7] [26], 
      \intermediateWiresStage1[7] [25], \intermediateWiresStage1[7] [24], 
      \intermediateWiresStage1[7] [23], \intermediateWiresStage1[7] [22], 
      \intermediateWiresStage1[7] [21], \intermediateWiresStage1[7] [20], 
      \intermediateWiresStage1[7] [19], \intermediateWiresStage1[7] [18], 
      \intermediateWiresStage1[7] [17], \intermediateWiresStage1[7] [16], 
      \intermediateWiresStage1[7] [15], \intermediateWiresStage1[7] [14], 
      \intermediateWiresStage1[7] [13], \intermediateWiresStage1[7] [12], 
      \intermediateWiresStage1[7] [11], uc_2122, uc_2123, uc_2124, uc_2125, 
      uc_2126, uc_2127, uc_2128, uc_2129, uc_2130, uc_2131, uc_2132}), .C({1'b0, 
      uc_2133, uc_2134, uc_2135, uc_2136, uc_2137, uc_2138, uc_2139, uc_2140, 
      uc_2141, uc_2142, uc_2143, uc_2144, uc_2145, uc_2146, uc_2147, uc_2148, 
      uc_2149, uc_2150, uc_2151, uc_2152, uc_2153, uc_2154, uc_2155, uc_2156, 
      uc_2157, uc_2158, uc_2159, uc_2160, \intermediateWiresStage1[8] [34], 
      \intermediateWiresStage1[8] [33], \intermediateWiresStage1[8] [32], 
      \intermediateWiresStage1[8] [31], \intermediateWiresStage1[8] [30], 
      \intermediateWiresStage1[8] [29], \intermediateWiresStage1[8] [28], 
      \intermediateWiresStage1[8] [27], \intermediateWiresStage1[8] [26], 
      \intermediateWiresStage1[8] [25], \intermediateWiresStage1[8] [24], 
      \intermediateWiresStage1[8] [23], \intermediateWiresStage1[8] [22], 
      \intermediateWiresStage1[8] [21], \intermediateWiresStage1[8] [20], 
      \intermediateWiresStage1[8] [19], \intermediateWiresStage1[8] [18], 
      \intermediateWiresStage1[8] [17], \intermediateWiresStage1[8] [16], 
      \intermediateWiresStage1[8] [15], \intermediateWiresStage1[8] [14], 
      \intermediateWiresStage1[8] [13], normalizedWires[780], uc_2161, uc_2162, 
      uc_2163, uc_2164, uc_2165, uc_2166, uc_2167, uc_2168, uc_2169, uc_2170, 
      uc_2171, uc_2172}));
   CSAlike__2_1765 genblk3_1_parallelAdderStage2 (.result({uc_2173, uc_2174, 
      uc_2175, uc_2176, uc_2177, uc_2178, uc_2179, uc_2180, uc_2181, uc_2182, 
      uc_2183, uc_2184, uc_2185, uc_2186, uc_2187, uc_2188, uc_2189, uc_2190, 
      uc_2191, uc_2192, uc_2193, uc_2194, uc_2195, uc_2196, uc_2197, uc_2198, 
      uc_2199, uc_2200, uc_2201, uc_2202, uc_2203, uc_2204, 
      \intermediateWiresStage2[2] [31], \intermediateWiresStage2[2] [30], 
      \intermediateWiresStage2[2] [29], \intermediateWiresStage2[2] [28], 
      \intermediateWiresStage2[2] [27], \intermediateWiresStage2[2] [26], 
      \intermediateWiresStage2[2] [25], \intermediateWiresStage2[2] [24], 
      \intermediateWiresStage2[2] [23], \intermediateWiresStage2[2] [22], 
      \intermediateWiresStage2[2] [21], \intermediateWiresStage2[2] [20], 
      \intermediateWiresStage2[2] [19], \intermediateWiresStage2[2] [18], 
      \intermediateWiresStage2[2] [17], \intermediateWiresStage2[2] [16], 
      \intermediateWiresStage2[2] [15], \intermediateWiresStage2[2] [14], 
      \intermediateWiresStage2[2] [13], \intermediateWiresStage2[2] [12], 
      \intermediateWiresStage2[2] [11], \intermediateWiresStage2[2] [10], 
      \intermediateWiresStage2[2] [9], \intermediateWiresStage2[2] [8], 
      \intermediateWiresStage2[2] [7], \intermediateWiresStage2[2] [6], uc_2205, 
      uc_2206, uc_2207, uc_2208, uc_2209, uc_2210}), .carry({uc_2211, uc_2212, 
      uc_2213, uc_2214, uc_2215, uc_2216, uc_2217, uc_2218, uc_2219, uc_2220, 
      uc_2221, uc_2222, uc_2223, uc_2224, uc_2225, uc_2226, uc_2227, uc_2228, 
      uc_2229, uc_2230, uc_2231, uc_2232, uc_2233, uc_2234, uc_2235, uc_2236, 
      uc_2237, uc_2238, uc_2239, uc_2240, uc_2241, 
      \intermediateWiresStage2[3] [32], \intermediateWiresStage2[3] [31], 
      \intermediateWiresStage2[3] [30], \intermediateWiresStage2[3] [29], 
      \intermediateWiresStage2[3] [28], \intermediateWiresStage2[3] [27], 
      \intermediateWiresStage2[3] [26], \intermediateWiresStage2[3] [25], 
      \intermediateWiresStage2[3] [24], \intermediateWiresStage2[3] [23], 
      \intermediateWiresStage2[3] [22], \intermediateWiresStage2[3] [21], 
      \intermediateWiresStage2[3] [20], \intermediateWiresStage2[3] [19], 
      \intermediateWiresStage2[3] [18], \intermediateWiresStage2[3] [17], 
      \intermediateWiresStage2[3] [16], \intermediateWiresStage2[3] [15], 
      \intermediateWiresStage2[3] [14], \intermediateWiresStage2[3] [13], 
      \intermediateWiresStage2[3] [12], \intermediateWiresStage2[3] [11], 
      \intermediateWiresStage2[3] [10], \intermediateWiresStage2[3] [9], 
      \intermediateWiresStage2[3] [8], \intermediateWiresStage2[3] [7], uc_2242, 
      uc_2243, uc_2244, uc_2245, uc_2246, uc_2247, uc_2248}), .A({1'b0, uc_2249, 
      uc_2250, uc_2251, uc_2252, uc_2253, uc_2254, uc_2255, uc_2256, uc_2257, 
      uc_2258, uc_2259, uc_2260, uc_2261, uc_2262, uc_2263, uc_2264, uc_2265, 
      uc_2266, uc_2267, uc_2268, uc_2269, uc_2270, uc_2271, uc_2272, uc_2273, 
      uc_2274, uc_2275, uc_2276, uc_2277, uc_2278, uc_2279, uc_2280, uc_2281, 
      uc_2282, \intermediateWiresStage1[3] [28], 
      \intermediateWiresStage1[3] [27], \intermediateWiresStage1[3] [26], 
      \intermediateWiresStage1[3] [25], \intermediateWiresStage1[3] [24], 
      \intermediateWiresStage1[3] [23], \intermediateWiresStage1[3] [22], 
      \intermediateWiresStage1[3] [21], \intermediateWiresStage1[3] [20], 
      \intermediateWiresStage1[3] [19], \intermediateWiresStage1[3] [18], 
      \intermediateWiresStage1[3] [17], \intermediateWiresStage1[3] [16], 
      \intermediateWiresStage1[3] [15], \intermediateWiresStage1[3] [14], 
      \intermediateWiresStage1[3] [13], \intermediateWiresStage1[3] [12], 
      \intermediateWiresStage1[3] [11], \intermediateWiresStage1[3] [10], 
      \intermediateWiresStage1[3] [9], \intermediateWiresStage1[3] [8], 
      \intermediateWiresStage1[3] [7], \intermediateWiresStage1[3] [6], uc_2283, 
      uc_2284, uc_2285, uc_2286, uc_2287, uc_2288}), .B({1'b0, uc_2289, uc_2290, 
      uc_2291, uc_2292, uc_2293, uc_2294, uc_2295, uc_2296, uc_2297, uc_2298, 
      uc_2299, uc_2300, uc_2301, uc_2302, uc_2303, uc_2304, uc_2305, uc_2306, 
      uc_2307, uc_2308, uc_2309, uc_2310, uc_2311, uc_2312, uc_2313, uc_2314, 
      uc_2315, uc_2316, uc_2317, uc_2318, uc_2319, normalizedWires[543], 
      \intermediateWiresStage1[4] [30], \intermediateWiresStage1[4] [29], 
      \intermediateWiresStage1[4] [28], \intermediateWiresStage1[4] [27], 
      \intermediateWiresStage1[4] [26], \intermediateWiresStage1[4] [25], 
      \intermediateWiresStage1[4] [24], \intermediateWiresStage1[4] [23], 
      \intermediateWiresStage1[4] [22], \intermediateWiresStage1[4] [21], 
      \intermediateWiresStage1[4] [20], \intermediateWiresStage1[4] [19], 
      \intermediateWiresStage1[4] [18], \intermediateWiresStage1[4] [17], 
      \intermediateWiresStage1[4] [16], \intermediateWiresStage1[4] [15], 
      \intermediateWiresStage1[4] [14], \intermediateWiresStage1[4] [13], 
      \intermediateWiresStage1[4] [12], \intermediateWiresStage1[4] [11], 
      \intermediateWiresStage1[4] [10], \intermediateWiresStage1[4] [9], 
      \intermediateWiresStage1[4] [8], \intermediateWiresStage1[4] [7], 
      normalizedWires[390], uc_2320, uc_2321, uc_2322, uc_2323, uc_2324, uc_2325}), 
      .C({1'b0, uc_2326, uc_2327, uc_2328, uc_2329, uc_2330, uc_2331, uc_2332, 
      uc_2333, uc_2334, uc_2335, uc_2336, uc_2337, uc_2338, uc_2339, uc_2340, 
      uc_2341, uc_2342, uc_2343, uc_2344, uc_2345, uc_2346, uc_2347, uc_2348, 
      uc_2349, uc_2350, uc_2351, uc_2352, uc_2353, uc_2354, uc_2355, uc_2356, 
      \intermediateWiresStage1[5] [31], \intermediateWiresStage1[5] [30], 
      \intermediateWiresStage1[5] [29], \intermediateWiresStage1[5] [28], 
      \intermediateWiresStage1[5] [27], \intermediateWiresStage1[5] [26], 
      \intermediateWiresStage1[5] [25], \intermediateWiresStage1[5] [24], 
      \intermediateWiresStage1[5] [23], \intermediateWiresStage1[5] [22], 
      \intermediateWiresStage1[5] [21], \intermediateWiresStage1[5] [20], 
      \intermediateWiresStage1[5] [19], \intermediateWiresStage1[5] [18], 
      \intermediateWiresStage1[5] [17], \intermediateWiresStage1[5] [16], 
      \intermediateWiresStage1[5] [15], \intermediateWiresStage1[5] [14], 
      \intermediateWiresStage1[5] [13], \intermediateWiresStage1[5] [12], 
      \intermediateWiresStage1[5] [11], \intermediateWiresStage1[5] [10], 
      \intermediateWiresStage1[5] [9], \intermediateWiresStage1[5] [8], uc_2357, 
      uc_2358, uc_2359, uc_2360, uc_2361, uc_2362, uc_2363, uc_2364}));
   CSAlike__0_113 genblk3_0_parallelAdderStage2 (.result({uc_2365, uc_2366, 
      uc_2367, uc_2368, uc_2369, uc_2370, uc_2371, uc_2372, uc_2373, uc_2374, 
      uc_2375, uc_2376, uc_2377, uc_2378, uc_2379, uc_2380, uc_2381, uc_2382, 
      uc_2383, uc_2384, uc_2385, uc_2386, uc_2387, uc_2388, uc_2389, uc_2390, 
      uc_2391, uc_2392, uc_2393, uc_2394, uc_2395, uc_2396, uc_2397, uc_2398, 
      uc_2399, uc_2400, uc_2401, uc_2402, \intermediateWiresStage2[0] [25], 
      \intermediateWiresStage2[0] [24], \intermediateWiresStage2[0] [23], 
      \intermediateWiresStage2[0] [22], \intermediateWiresStage2[0] [21], 
      \intermediateWiresStage2[0] [20], \intermediateWiresStage2[0] [19], 
      \intermediateWiresStage2[0] [18], \intermediateWiresStage2[0] [17], 
      \intermediateWiresStage2[0] [16], \intermediateWiresStage2[0] [15], 
      \intermediateWiresStage2[0] [14], \intermediateWiresStage2[0] [13], 
      \intermediateWiresStage2[0] [12], \intermediateWiresStage2[0] [11], 
      \intermediateWiresStage2[0] [10], \intermediateWiresStage2[0] [9], 
      \intermediateWiresStage2[0] [8], \intermediateWiresStage2[0] [7], 
      \intermediateWiresStage2[0] [6], \intermediateWiresStage2[0] [5], 
      \intermediateWiresStage2[0] [4], \intermediateWiresStage2[0] [3], uc_2403, 
      uc_2404, uc_2405}), .carry({uc_2406, uc_2407, uc_2408, uc_2409, uc_2410, 
      uc_2411, uc_2412, uc_2413, uc_2414, uc_2415, uc_2416, uc_2417, uc_2418, 
      uc_2419, uc_2420, uc_2421, uc_2422, uc_2423, uc_2424, uc_2425, uc_2426, 
      uc_2427, uc_2428, uc_2429, uc_2430, uc_2431, uc_2432, uc_2433, uc_2434, 
      uc_2435, uc_2436, uc_2437, uc_2438, uc_2439, uc_2440, uc_2441, uc_2442, 
      \intermediateWiresStage2[1] [26], \intermediateWiresStage2[1] [25], 
      \intermediateWiresStage2[1] [24], \intermediateWiresStage2[1] [23], 
      \intermediateWiresStage2[1] [22], \intermediateWiresStage2[1] [21], 
      \intermediateWiresStage2[1] [20], \intermediateWiresStage2[1] [19], 
      \intermediateWiresStage2[1] [18], \intermediateWiresStage2[1] [17], 
      \intermediateWiresStage2[1] [16], \intermediateWiresStage2[1] [15], 
      \intermediateWiresStage2[1] [14], \intermediateWiresStage2[1] [13], 
      \intermediateWiresStage2[1] [12], \intermediateWiresStage2[1] [11], 
      \intermediateWiresStage2[1] [10], \intermediateWiresStage2[1] [9], 
      \intermediateWiresStage2[1] [8], \intermediateWiresStage2[1] [7], 
      \intermediateWiresStage2[1] [6], \intermediateWiresStage2[1] [5], 
      \intermediateWiresStage2[1] [4], \intermediateWiresStage2[1] [3], uc_2443, 
      uc_2444, uc_2445}), .A({1'b0, uc_2446, uc_2447, uc_2448, uc_2449, uc_2450, 
      uc_2451, uc_2452, uc_2453, uc_2454, uc_2455, uc_2456, uc_2457, uc_2458, 
      uc_2459, uc_2460, uc_2461, uc_2462, uc_2463, uc_2464, uc_2465, uc_2466, 
      uc_2467, uc_2468, uc_2469, uc_2470, uc_2471, uc_2472, uc_2473, uc_2474, 
      uc_2475, uc_2476, uc_2477, uc_2478, uc_2479, uc_2480, uc_2481, uc_2482, 
      normalizedWires[153], \intermediateWiresStage1[0] [24], 
      \intermediateWiresStage1[0] [23], \intermediateWiresStage1[0] [22], 
      \intermediateWiresStage1[0] [21], \intermediateWiresStage1[0] [20], 
      \intermediateWiresStage1[0] [19], \intermediateWiresStage1[0] [18], 
      \intermediateWiresStage1[0] [17], \intermediateWiresStage1[0] [16], 
      \intermediateWiresStage1[0] [15], \intermediateWiresStage1[0] [14], 
      \intermediateWiresStage1[0] [13], \intermediateWiresStage1[0] [12], 
      \intermediateWiresStage1[0] [11], \intermediateWiresStage1[0] [10], 
      \intermediateWiresStage1[0] [9], \intermediateWiresStage1[0] [8], 
      \intermediateWiresStage1[0] [7], \intermediateWiresStage1[0] [6], 
      \intermediateWiresStage1[0] [5], \intermediateWiresStage1[0] [4], 
      \intermediateWiresStage1[0] [3], \intermediateWiresStage1[0] [2], uc_2483, 
      uc_2484}), .B({1'b0, uc_2485, uc_2486, uc_2487, uc_2488, uc_2489, uc_2490, 
      uc_2491, uc_2492, uc_2493, uc_2494, uc_2495, uc_2496, uc_2497, uc_2498, 
      uc_2499, uc_2500, uc_2501, uc_2502, uc_2503, uc_2504, uc_2505, uc_2506, 
      uc_2507, uc_2508, uc_2509, uc_2510, uc_2511, uc_2512, uc_2513, uc_2514, 
      uc_2515, uc_2516, uc_2517, uc_2518, uc_2519, uc_2520, uc_2521, 
      \intermediateWiresStage1[1] [25], \intermediateWiresStage1[1] [24], 
      \intermediateWiresStage1[1] [23], \intermediateWiresStage1[1] [22], 
      \intermediateWiresStage1[1] [21], \intermediateWiresStage1[1] [20], 
      \intermediateWiresStage1[1] [19], \intermediateWiresStage1[1] [18], 
      \intermediateWiresStage1[1] [17], \intermediateWiresStage1[1] [16], 
      \intermediateWiresStage1[1] [15], \intermediateWiresStage1[1] [14], 
      \intermediateWiresStage1[1] [13], \intermediateWiresStage1[1] [12], 
      \intermediateWiresStage1[1] [11], \intermediateWiresStage1[1] [10], 
      \intermediateWiresStage1[1] [9], \intermediateWiresStage1[1] [8], 
      \intermediateWiresStage1[1] [7], \intermediateWiresStage1[1] [6], 
      \intermediateWiresStage1[1] [5], \intermediateWiresStage1[1] [4], 
      \intermediateWiresStage1[1] [3], \intermediateWiresStage1[1] [2], uc_2522, 
      uc_2523}), .C({1'b0, uc_2524, uc_2525, uc_2526, uc_2527, uc_2528, uc_2529, 
      uc_2530, uc_2531, uc_2532, uc_2533, uc_2534, uc_2535, uc_2536, uc_2537, 
      uc_2538, uc_2539, uc_2540, uc_2541, uc_2542, uc_2543, uc_2544, uc_2545, 
      uc_2546, uc_2547, uc_2548, uc_2549, uc_2550, uc_2551, uc_2552, uc_2553, 
      uc_2554, uc_2555, uc_2556, uc_2557, uc_2558, uc_2559, uc_2560, 
      \intermediateWiresStage1[2] [25], \intermediateWiresStage1[2] [24], 
      \intermediateWiresStage1[2] [23], \intermediateWiresStage1[2] [22], 
      \intermediateWiresStage1[2] [21], \intermediateWiresStage1[2] [20], 
      \intermediateWiresStage1[2] [19], \intermediateWiresStage1[2] [18], 
      \intermediateWiresStage1[2] [17], \intermediateWiresStage1[2] [16], 
      \intermediateWiresStage1[2] [15], \intermediateWiresStage1[2] [14], 
      \intermediateWiresStage1[2] [13], \intermediateWiresStage1[2] [12], 
      \intermediateWiresStage1[2] [11], \intermediateWiresStage1[2] [10], 
      \intermediateWiresStage1[2] [9], \intermediateWiresStage1[2] [8], 
      \intermediateWiresStage1[2] [7], \intermediateWiresStage1[2] [6], 
      \intermediateWiresStage1[2] [5], \intermediateWiresStage1[2] [4], 
      normalizedWires[195], uc_2561, uc_2562, uc_2563}));
   CSAlike__3_753 genblk4_3_parallelAdderStage3 (.result({uc_2564, uc_2565, 
      uc_2566, uc_2567, uc_2568, uc_2569, uc_2570, uc_2571, uc_2572, uc_2573, 
      uc_2574, uc_2575, uc_2576, uc_2577, uc_2578, uc_2579, uc_2580, uc_2581, 
      uc_2582, \intermediateWiresStage3[6] [44], 
      \intermediateWiresStage3[6] [43], \intermediateWiresStage3[6] [42], 
      \intermediateWiresStage3[6] [41], \intermediateWiresStage3[6] [40], 
      \intermediateWiresStage3[6] [39], \intermediateWiresStage3[6] [38], 
      \intermediateWiresStage3[6] [37], \intermediateWiresStage3[6] [36], 
      \intermediateWiresStage3[6] [35], \intermediateWiresStage3[6] [34], 
      \intermediateWiresStage3[6] [33], \intermediateWiresStage3[6] [32], 
      \intermediateWiresStage3[6] [31], \intermediateWiresStage3[6] [30], 
      \intermediateWiresStage3[6] [29], \intermediateWiresStage3[6] [28], 
      \intermediateWiresStage3[6] [27], \intermediateWiresStage3[6] [26], 
      \intermediateWiresStage3[6] [25], \intermediateWiresStage3[6] [24], 
      \intermediateWiresStage3[6] [23], uc_2583, uc_2584, uc_2585, uc_2586, 
      uc_2587, uc_2588, uc_2589, uc_2590, uc_2591, uc_2592, uc_2593, uc_2594, 
      uc_2595, uc_2596, uc_2597, uc_2598, uc_2599, uc_2600, uc_2601, uc_2602, 
      uc_2603, uc_2604, uc_2605}), .carry({uc_2606, uc_2607, uc_2608, uc_2609, 
      uc_2610, uc_2611, uc_2612, uc_2613, uc_2614, uc_2615, uc_2616, uc_2617, 
      uc_2618, uc_2619, uc_2620, uc_2621, uc_2622, uc_2623, 
      \intermediateWiresStage3[7] [45], \intermediateWiresStage3[7] [44], 
      \intermediateWiresStage3[7] [43], \intermediateWiresStage3[7] [42], 
      \intermediateWiresStage3[7] [41], \intermediateWiresStage3[7] [40], 
      \intermediateWiresStage3[7] [39], \intermediateWiresStage3[7] [38], 
      \intermediateWiresStage3[7] [37], \intermediateWiresStage3[7] [36], 
      \intermediateWiresStage3[7] [35], \intermediateWiresStage3[7] [34], 
      \intermediateWiresStage3[7] [33], \intermediateWiresStage3[7] [32], 
      \intermediateWiresStage3[7] [31], \intermediateWiresStage3[7] [30], 
      \intermediateWiresStage3[7] [29], \intermediateWiresStage3[7] [28], 
      \intermediateWiresStage3[7] [27], \intermediateWiresStage3[7] [26], 
      \intermediateWiresStage3[7] [25], \intermediateWiresStage3[7] [24], 
      uc_2624, uc_2625, uc_2626, uc_2627, uc_2628, uc_2629, uc_2630, uc_2631, 
      uc_2632, uc_2633, uc_2634, uc_2635, uc_2636, uc_2637, uc_2638, uc_2639, 
      uc_2640, uc_2641, uc_2642, uc_2643, uc_2644, uc_2645, uc_2646, uc_2647}), 
      .A({1'b0, uc_2648, uc_2649, uc_2650, uc_2651, uc_2652, uc_2653, uc_2654, 
      uc_2655, uc_2656, uc_2657, uc_2658, uc_2659, uc_2660, uc_2661, uc_2662, 
      uc_2663, uc_2664, uc_2665, \intermediateWiresStage2[9] [44], 
      \intermediateWiresStage2[9] [43], \intermediateWiresStage2[9] [42], 
      \intermediateWiresStage2[9] [41], \intermediateWiresStage2[9] [40], 
      \intermediateWiresStage2[9] [39], \intermediateWiresStage2[9] [38], 
      \intermediateWiresStage2[9] [37], \intermediateWiresStage2[9] [36], 
      \intermediateWiresStage2[9] [35], \intermediateWiresStage2[9] [34], 
      \intermediateWiresStage2[9] [33], \intermediateWiresStage2[9] [32], 
      \intermediateWiresStage2[9] [31], \intermediateWiresStage2[9] [30], 
      \intermediateWiresStage2[9] [29], \intermediateWiresStage2[9] [28], 
      \intermediateWiresStage2[9] [27], \intermediateWiresStage2[9] [26], 
      \intermediateWiresStage2[9] [25], \intermediateWiresStage2[9] [24], 
      \intermediateWiresStage2[9] [23], uc_2666, uc_2667, uc_2668, uc_2669, 
      uc_2670, uc_2671, uc_2672, uc_2673, uc_2674, uc_2675, uc_2676, uc_2677, 
      uc_2678, uc_2679, uc_2680, uc_2681, uc_2682, uc_2683, uc_2684, uc_2685, 
      uc_2686, uc_2687, uc_2688}), .B({1'b0, uc_2689, uc_2690, uc_2691, uc_2692, 
      uc_2693, uc_2694, uc_2695, uc_2696, uc_2697, uc_2698, uc_2699, uc_2700, 
      uc_2701, uc_2702, uc_2703, uc_2704, uc_2705, uc_2706, 
      \intermediateWiresStage1[15] [44], \intermediateWiresStage1[15] [43], 
      \intermediateWiresStage1[15] [42], \intermediateWiresStage1[15] [41], 
      \intermediateWiresStage1[15] [40], \intermediateWiresStage1[15] [39], 
      \intermediateWiresStage1[15] [38], \intermediateWiresStage1[15] [37], 
      \intermediateWiresStage1[15] [36], \intermediateWiresStage1[15] [35], 
      \intermediateWiresStage1[15] [34], \intermediateWiresStage1[15] [33], 
      \intermediateWiresStage1[15] [32], \intermediateWiresStage1[15] [31], 
      \intermediateWiresStage1[15] [30], \intermediateWiresStage1[15] [29], 
      \intermediateWiresStage1[15] [28], \intermediateWiresStage1[15] [27], 
      \intermediateWiresStage1[15] [26], \intermediateWiresStage1[15] [25], 
      \intermediateWiresStage1[15] [24], \intermediateWiresStage1[15] [23], 
      uc_2707, uc_2708, uc_2709, uc_2710, uc_2711, uc_2712, uc_2713, uc_2714, 
      uc_2715, uc_2716, uc_2717, uc_2718, uc_2719, uc_2720, uc_2721, uc_2722, 
      uc_2723, uc_2724, uc_2725, uc_2726, uc_2727, uc_2728, uc_2729}), .C({1'b0, 
      uc_2730, uc_2731, uc_2732, uc_2733, uc_2734, uc_2735, uc_2736, uc_2737, 
      uc_2738, uc_2739, uc_2740, uc_2741, uc_2742, uc_2743, uc_2744, uc_2745, 
      uc_2746, uc_2747, uc_2748, uc_2749, uc_2750, uc_2751, uc_2752, uc_2753, 
      uc_2754, uc_2755, uc_2756, uc_2757, uc_2758, uc_2759, uc_2760, uc_2761, 
      uc_2762, uc_2763, uc_2764, uc_2765, uc_2766, uc_2767, uc_2768, uc_2769, 
      uc_2770, uc_2771, uc_2772, uc_2773, uc_2774, uc_2775, uc_2776, uc_2777, 
      uc_2778, uc_2779, uc_2780, uc_2781, uc_2782, uc_2783, uc_2784, uc_2785, 
      uc_2786, uc_2787, uc_2788, uc_2789, uc_2790, uc_2791, uc_2792}));
   CSAlike__3_1006 genblk4_2_parallelAdderStage3 (.result({uc_2793, uc_2794, 
      uc_2795, uc_2796, uc_2797, uc_2798, uc_2799, uc_2800, uc_2801, uc_2802, 
      uc_2803, uc_2804, uc_2805, uc_2806, uc_2807, uc_2808, uc_2809, uc_2810, 
      uc_2811, uc_2812, uc_2813, uc_2814, \intermediateWiresStage3[4] [41], 
      \intermediateWiresStage3[4] [40], \intermediateWiresStage3[4] [39], 
      \intermediateWiresStage3[4] [38], \intermediateWiresStage3[4] [37], 
      \intermediateWiresStage3[4] [36], \intermediateWiresStage3[4] [35], 
      \intermediateWiresStage3[4] [34], \intermediateWiresStage3[4] [33], 
      \intermediateWiresStage3[4] [32], \intermediateWiresStage3[4] [31], 
      \intermediateWiresStage3[4] [30], \intermediateWiresStage3[4] [29], 
      \intermediateWiresStage3[4] [28], \intermediateWiresStage3[4] [27], 
      \intermediateWiresStage3[4] [26], \intermediateWiresStage3[4] [25], 
      \intermediateWiresStage3[4] [24], \intermediateWiresStage3[4] [23], 
      \intermediateWiresStage3[4] [22], \intermediateWiresStage3[4] [21], 
      \intermediateWiresStage3[4] [20], \intermediateWiresStage3[4] [19], 
      \intermediateWiresStage3[4] [18], \intermediateWiresStage3[4] [17], 
      \intermediateWiresStage3[4] [16], uc_2815, uc_2816, uc_2817, uc_2818, 
      uc_2819, uc_2820, uc_2821, uc_2822, uc_2823, uc_2824, uc_2825, uc_2826, 
      uc_2827, uc_2828, uc_2829, uc_2830}), .carry({uc_2831, uc_2832, uc_2833, 
      uc_2834, uc_2835, uc_2836, uc_2837, uc_2838, uc_2839, uc_2840, uc_2841, 
      uc_2842, uc_2843, uc_2844, uc_2845, uc_2846, uc_2847, uc_2848, uc_2849, 
      uc_2850, uc_2851, \intermediateWiresStage3[5] [42], 
      \intermediateWiresStage3[5] [41], \intermediateWiresStage3[5] [40], 
      \intermediateWiresStage3[5] [39], \intermediateWiresStage3[5] [38], 
      \intermediateWiresStage3[5] [37], \intermediateWiresStage3[5] [36], 
      \intermediateWiresStage3[5] [35], \intermediateWiresStage3[5] [34], 
      \intermediateWiresStage3[5] [33], \intermediateWiresStage3[5] [32], 
      \intermediateWiresStage3[5] [31], \intermediateWiresStage3[5] [30], 
      \intermediateWiresStage3[5] [29], \intermediateWiresStage3[5] [28], 
      \intermediateWiresStage3[5] [27], \intermediateWiresStage3[5] [26], 
      \intermediateWiresStage3[5] [25], \intermediateWiresStage3[5] [24], 
      \intermediateWiresStage3[5] [23], \intermediateWiresStage3[5] [22], 
      \intermediateWiresStage3[5] [21], \intermediateWiresStage3[5] [20], 
      \intermediateWiresStage3[5] [19], \intermediateWiresStage3[5] [18], 
      \intermediateWiresStage3[5] [17], uc_2852, uc_2853, uc_2854, uc_2855, 
      uc_2856, uc_2857, uc_2858, uc_2859, uc_2860, uc_2861, uc_2862, uc_2863, 
      uc_2864, uc_2865, uc_2866, uc_2867, uc_2868}), .A({1'b0, uc_2869, uc_2870, 
      uc_2871, uc_2872, uc_2873, uc_2874, uc_2875, uc_2876, uc_2877, uc_2878, 
      uc_2879, uc_2880, uc_2881, uc_2882, uc_2883, uc_2884, uc_2885, uc_2886, 
      uc_2887, uc_2888, uc_2889, uc_2890, \intermediateWiresStage2[6] [40], 
      \intermediateWiresStage2[6] [39], \intermediateWiresStage2[6] [38], 
      \intermediateWiresStage2[6] [37], \intermediateWiresStage2[6] [36], 
      \intermediateWiresStage2[6] [35], \intermediateWiresStage2[6] [34], 
      \intermediateWiresStage2[6] [33], \intermediateWiresStage2[6] [32], 
      \intermediateWiresStage2[6] [31], \intermediateWiresStage2[6] [30], 
      \intermediateWiresStage2[6] [29], \intermediateWiresStage2[6] [28], 
      \intermediateWiresStage2[6] [27], \intermediateWiresStage2[6] [26], 
      \intermediateWiresStage2[6] [25], \intermediateWiresStage2[6] [24], 
      \intermediateWiresStage2[6] [23], \intermediateWiresStage2[6] [22], 
      \intermediateWiresStage2[6] [21], \intermediateWiresStage2[6] [20], 
      \intermediateWiresStage2[6] [19], \intermediateWiresStage2[6] [18], 
      \intermediateWiresStage2[6] [17], \intermediateWiresStage2[6] [16], 
      uc_2891, uc_2892, uc_2893, uc_2894, uc_2895, uc_2896, uc_2897, uc_2898, 
      uc_2899, uc_2900, uc_2901, uc_2902, uc_2903, uc_2904, uc_2905, uc_2906}), 
      .B({1'b0, uc_2907, uc_2908, uc_2909, uc_2910, uc_2911, uc_2912, uc_2913, 
      uc_2914, uc_2915, uc_2916, uc_2917, uc_2918, uc_2919, uc_2920, uc_2921, 
      uc_2922, uc_2923, uc_2924, uc_2925, uc_2926, uc_2927, 
      \intermediateWiresStage2[7] [41], \intermediateWiresStage2[7] [40], 
      \intermediateWiresStage2[7] [39], \intermediateWiresStage2[7] [38], 
      \intermediateWiresStage2[7] [37], \intermediateWiresStage2[7] [36], 
      \intermediateWiresStage2[7] [35], \intermediateWiresStage2[7] [34], 
      \intermediateWiresStage2[7] [33], \intermediateWiresStage2[7] [32], 
      \intermediateWiresStage2[7] [31], \intermediateWiresStage2[7] [30], 
      \intermediateWiresStage2[7] [29], \intermediateWiresStage2[7] [28], 
      \intermediateWiresStage2[7] [27], \intermediateWiresStage2[7] [26], 
      \intermediateWiresStage2[7] [25], \intermediateWiresStage2[7] [24], 
      \intermediateWiresStage2[7] [23], \intermediateWiresStage2[7] [22], 
      \intermediateWiresStage2[7] [21], \intermediateWiresStage2[7] [20], 
      \intermediateWiresStage2[7] [19], \intermediateWiresStage2[7] [18], 
      \intermediateWiresStage2[7] [17], \intermediateWiresStage2[7] [16], 
      uc_2928, uc_2929, uc_2930, uc_2931, uc_2932, uc_2933, uc_2934, uc_2935, 
      uc_2936, uc_2937, uc_2938, uc_2939, uc_2940, uc_2941, uc_2942, uc_2943}), 
      .C({1'b0, uc_2944, uc_2945, uc_2946, uc_2947, uc_2948, uc_2949, uc_2950, 
      uc_2951, uc_2952, uc_2953, uc_2954, uc_2955, uc_2956, uc_2957, uc_2958, 
      uc_2959, uc_2960, uc_2961, uc_2962, uc_2963, uc_2964, 
      \intermediateWiresStage2[8] [41], \intermediateWiresStage2[8] [40], 
      \intermediateWiresStage2[8] [39], \intermediateWiresStage2[8] [38], 
      \intermediateWiresStage2[8] [37], \intermediateWiresStage2[8] [36], 
      \intermediateWiresStage2[8] [35], \intermediateWiresStage2[8] [34], 
      \intermediateWiresStage2[8] [33], \intermediateWiresStage2[8] [32], 
      \intermediateWiresStage2[8] [31], \intermediateWiresStage2[8] [30], 
      \intermediateWiresStage2[8] [29], \intermediateWiresStage2[8] [28], 
      \intermediateWiresStage2[8] [27], \intermediateWiresStage2[8] [26], 
      \intermediateWiresStage2[8] [25], \intermediateWiresStage2[8] [24], 
      \intermediateWiresStage2[8] [23], \intermediateWiresStage2[8] [22], 
      \intermediateWiresStage2[8] [21], \intermediateWiresStage2[8] [20], 
      \intermediateWiresStage1[12] [19], normalizedWires[1170], uc_2965, uc_2966, 
      uc_2967, uc_2968, uc_2969, uc_2970, uc_2971, uc_2972, uc_2973, uc_2974, 
      uc_2975, uc_2976, uc_2977, uc_2978, uc_2979, uc_2980, uc_2981, uc_2982}));
   CSAlike__3_1259 genblk4_1_parallelAdderStage3 (.result({uc_2983, uc_2984, 
      uc_2985, uc_2986, uc_2987, uc_2988, uc_2989, uc_2990, uc_2991, uc_2992, 
      uc_2993, uc_2994, uc_2995, uc_2996, uc_2997, uc_2998, uc_2999, uc_3000, 
      uc_3001, uc_3002, uc_3003, uc_3004, uc_3005, uc_3006, uc_3007, uc_3008, 
      uc_3009, uc_3010, \intermediateWiresStage3[2] [35], 
      \intermediateWiresStage3[2] [34], \intermediateWiresStage3[2] [33], 
      \intermediateWiresStage3[2] [32], \intermediateWiresStage3[2] [31], 
      \intermediateWiresStage3[2] [30], \intermediateWiresStage3[2] [29], 
      \intermediateWiresStage3[2] [28], \intermediateWiresStage3[2] [27], 
      \intermediateWiresStage3[2] [26], \intermediateWiresStage3[2] [25], 
      \intermediateWiresStage3[2] [24], \intermediateWiresStage3[2] [23], 
      \intermediateWiresStage3[2] [22], \intermediateWiresStage3[2] [21], 
      \intermediateWiresStage3[2] [20], \intermediateWiresStage3[2] [19], 
      \intermediateWiresStage3[2] [18], \intermediateWiresStage3[2] [17], 
      \intermediateWiresStage3[2] [16], \intermediateWiresStage3[2] [15], 
      \intermediateWiresStage3[2] [14], \intermediateWiresStage3[2] [13], 
      \intermediateWiresStage3[2] [12], \intermediateWiresStage3[2] [11], 
      \intermediateWiresStage3[2] [10], \intermediateWiresStage3[2] [9], uc_3011, 
      uc_3012, uc_3013, uc_3014, uc_3015, uc_3016, uc_3017, uc_3018, uc_3019}), 
      .carry({uc_3020, uc_3021, uc_3022, uc_3023, uc_3024, uc_3025, uc_3026, 
      uc_3027, uc_3028, uc_3029, uc_3030, uc_3031, uc_3032, uc_3033, uc_3034, 
      uc_3035, uc_3036, uc_3037, uc_3038, uc_3039, uc_3040, uc_3041, uc_3042, 
      uc_3043, uc_3044, uc_3045, uc_3046, \intermediateWiresStage3[3] [36], 
      \intermediateWiresStage3[3] [35], \intermediateWiresStage3[3] [34], 
      \intermediateWiresStage3[3] [33], \intermediateWiresStage3[3] [32], 
      \intermediateWiresStage3[3] [31], \intermediateWiresStage3[3] [30], 
      \intermediateWiresStage3[3] [29], \intermediateWiresStage3[3] [28], 
      \intermediateWiresStage3[3] [27], \intermediateWiresStage3[3] [26], 
      \intermediateWiresStage3[3] [25], \intermediateWiresStage3[3] [24], 
      \intermediateWiresStage3[3] [23], \intermediateWiresStage3[3] [22], 
      \intermediateWiresStage3[3] [21], \intermediateWiresStage3[3] [20], 
      \intermediateWiresStage3[3] [19], \intermediateWiresStage3[3] [18], 
      \intermediateWiresStage3[3] [17], \intermediateWiresStage3[3] [16], 
      \intermediateWiresStage3[3] [15], \intermediateWiresStage3[3] [14], 
      \intermediateWiresStage3[3] [13], \intermediateWiresStage3[3] [12], 
      \intermediateWiresStage3[3] [11], \intermediateWiresStage3[3] [10], 
      uc_3047, uc_3048, uc_3049, uc_3050, uc_3051, uc_3052, uc_3053, uc_3054, 
      uc_3055, uc_3056}), .A({1'b0, uc_3057, uc_3058, uc_3059, uc_3060, uc_3061, 
      uc_3062, uc_3063, uc_3064, uc_3065, uc_3066, uc_3067, uc_3068, uc_3069, 
      uc_3070, uc_3071, uc_3072, uc_3073, uc_3074, uc_3075, uc_3076, uc_3077, 
      uc_3078, uc_3079, uc_3080, uc_3081, uc_3082, uc_3083, uc_3084, uc_3085, 
      uc_3086, \intermediateWiresStage2[3] [32], 
      \intermediateWiresStage2[3] [31], \intermediateWiresStage2[3] [30], 
      \intermediateWiresStage2[3] [29], \intermediateWiresStage2[3] [28], 
      \intermediateWiresStage2[3] [27], \intermediateWiresStage2[3] [26], 
      \intermediateWiresStage2[3] [25], \intermediateWiresStage2[3] [24], 
      \intermediateWiresStage2[3] [23], \intermediateWiresStage2[3] [22], 
      \intermediateWiresStage2[3] [21], \intermediateWiresStage2[3] [20], 
      \intermediateWiresStage2[3] [19], \intermediateWiresStage2[3] [18], 
      \intermediateWiresStage2[3] [17], \intermediateWiresStage2[3] [16], 
      \intermediateWiresStage2[3] [15], \intermediateWiresStage2[3] [14], 
      \intermediateWiresStage2[3] [13], \intermediateWiresStage2[3] [12], 
      \intermediateWiresStage2[3] [11], \intermediateWiresStage2[3] [10], 
      \intermediateWiresStage2[3] [9], uc_3087, uc_3088, uc_3089, uc_3090, 
      uc_3091, uc_3092, uc_3093, uc_3094, uc_3095}), .B({1'b0, uc_3096, uc_3097, 
      uc_3098, uc_3099, uc_3100, uc_3101, uc_3102, uc_3103, uc_3104, uc_3105, 
      uc_3106, uc_3107, uc_3108, uc_3109, uc_3110, uc_3111, uc_3112, uc_3113, 
      uc_3114, uc_3115, uc_3116, uc_3117, uc_3118, uc_3119, uc_3120, uc_3121, 
      uc_3122, \intermediateWiresStage1[8] [35], 
      \intermediateWiresStage2[4] [34], \intermediateWiresStage2[4] [33], 
      \intermediateWiresStage2[4] [32], \intermediateWiresStage2[4] [31], 
      \intermediateWiresStage2[4] [30], \intermediateWiresStage2[4] [29], 
      \intermediateWiresStage2[4] [28], \intermediateWiresStage2[4] [27], 
      \intermediateWiresStage2[4] [26], \intermediateWiresStage2[4] [25], 
      \intermediateWiresStage2[4] [24], \intermediateWiresStage2[4] [23], 
      \intermediateWiresStage2[4] [22], \intermediateWiresStage2[4] [21], 
      \intermediateWiresStage2[4] [20], \intermediateWiresStage2[4] [19], 
      \intermediateWiresStage2[4] [18], \intermediateWiresStage2[4] [17], 
      \intermediateWiresStage2[4] [16], \intermediateWiresStage2[4] [15], 
      \intermediateWiresStage2[4] [14], \intermediateWiresStage2[4] [13], 
      \intermediateWiresStage2[4] [12], \intermediateWiresStage2[4] [11], 
      \intermediateWiresStage1[6] [10], normalizedWires[585], uc_3123, uc_3124, 
      uc_3125, uc_3126, uc_3127, uc_3128, uc_3129, uc_3130, uc_3131}), .C({1'b0, 
      uc_3132, uc_3133, uc_3134, uc_3135, uc_3136, uc_3137, uc_3138, uc_3139, 
      uc_3140, uc_3141, uc_3142, uc_3143, uc_3144, uc_3145, uc_3146, uc_3147, 
      uc_3148, uc_3149, uc_3150, uc_3151, uc_3152, uc_3153, uc_3154, uc_3155, 
      uc_3156, uc_3157, uc_3158, \intermediateWiresStage2[5] [35], 
      \intermediateWiresStage2[5] [34], \intermediateWiresStage2[5] [33], 
      \intermediateWiresStage2[5] [32], \intermediateWiresStage2[5] [31], 
      \intermediateWiresStage2[5] [30], \intermediateWiresStage2[5] [29], 
      \intermediateWiresStage2[5] [28], \intermediateWiresStage2[5] [27], 
      \intermediateWiresStage2[5] [26], \intermediateWiresStage2[5] [25], 
      \intermediateWiresStage2[5] [24], \intermediateWiresStage2[5] [23], 
      \intermediateWiresStage2[5] [22], \intermediateWiresStage2[5] [21], 
      \intermediateWiresStage2[5] [20], \intermediateWiresStage2[5] [19], 
      \intermediateWiresStage2[5] [18], \intermediateWiresStage2[5] [17], 
      \intermediateWiresStage2[5] [16], \intermediateWiresStage2[5] [15], 
      \intermediateWiresStage2[5] [14], \intermediateWiresStage2[5] [13], 
      \intermediateWiresStage2[5] [12], uc_3159, uc_3160, uc_3161, uc_3162, 
      uc_3163, uc_3164, uc_3165, uc_3166, uc_3167, uc_3168, uc_3169, uc_3170}));
   CSAlike__0_118 genblk4_0_parallelAdderStage3 (.result({uc_3171, uc_3172, 
      uc_3173, uc_3174, uc_3175, uc_3176, uc_3177, uc_3178, uc_3179, uc_3180, 
      uc_3181, uc_3182, uc_3183, uc_3184, uc_3185, uc_3186, uc_3187, uc_3188, 
      uc_3189, uc_3190, uc_3191, uc_3192, uc_3193, uc_3194, uc_3195, uc_3196, 
      uc_3197, uc_3198, uc_3199, uc_3200, uc_3201, uc_3202, uc_3203, uc_3204, 
      uc_3205, \intermediateWiresStage3[0] [28], 
      \intermediateWiresStage3[0] [27], \intermediateWiresStage3[0] [26], 
      \intermediateWiresStage3[0] [25], \intermediateWiresStage3[0] [24], 
      \intermediateWiresStage3[0] [23], \intermediateWiresStage3[0] [22], 
      \intermediateWiresStage3[0] [21], \intermediateWiresStage3[0] [20], 
      \intermediateWiresStage3[0] [19], \intermediateWiresStage3[0] [18], 
      \intermediateWiresStage3[0] [17], \intermediateWiresStage3[0] [16], 
      \intermediateWiresStage3[0] [15], \intermediateWiresStage3[0] [14], 
      \intermediateWiresStage3[0] [13], \intermediateWiresStage3[0] [12], 
      \intermediateWiresStage3[0] [11], \intermediateWiresStage3[0] [10], 
      \intermediateWiresStage3[0] [9], \intermediateWiresStage3[0] [8], 
      \intermediateWiresStage3[0] [7], \intermediateWiresStage3[0] [6], 
      \intermediateWiresStage3[0] [5], \intermediateWiresStage3[0] [4], uc_3206, 
      uc_3207, uc_3208, uc_3209}), .carry({uc_3210, uc_3211, uc_3212, uc_3213, 
      uc_3214, uc_3215, uc_3216, uc_3217, uc_3218, uc_3219, uc_3220, uc_3221, 
      uc_3222, uc_3223, uc_3224, uc_3225, uc_3226, uc_3227, uc_3228, uc_3229, 
      uc_3230, uc_3231, uc_3232, uc_3233, uc_3234, uc_3235, uc_3236, uc_3237, 
      uc_3238, uc_3239, uc_3240, uc_3241, uc_3242, uc_3243, 
      \intermediateWiresStage3[1] [29], \intermediateWiresStage3[1] [28], 
      \intermediateWiresStage3[1] [27], \intermediateWiresStage3[1] [26], 
      \intermediateWiresStage3[1] [25], \intermediateWiresStage3[1] [24], 
      \intermediateWiresStage3[1] [23], \intermediateWiresStage3[1] [22], 
      \intermediateWiresStage3[1] [21], \intermediateWiresStage3[1] [20], 
      \intermediateWiresStage3[1] [19], \intermediateWiresStage3[1] [18], 
      \intermediateWiresStage3[1] [17], \intermediateWiresStage3[1] [16], 
      \intermediateWiresStage3[1] [15], \intermediateWiresStage3[1] [14], 
      \intermediateWiresStage3[1] [13], \intermediateWiresStage3[1] [12], 
      \intermediateWiresStage3[1] [11], \intermediateWiresStage3[1] [10], 
      \intermediateWiresStage3[1] [9], \intermediateWiresStage3[1] [8], 
      \intermediateWiresStage3[1] [7], \intermediateWiresStage3[1] [6], 
      \intermediateWiresStage3[1] [5], \intermediateWiresStage3[1] [4], uc_3244, 
      uc_3245, uc_3246, uc_3247}), .A({1'b0, uc_3248, uc_3249, uc_3250, uc_3251, 
      uc_3252, uc_3253, uc_3254, uc_3255, uc_3256, uc_3257, uc_3258, uc_3259, 
      uc_3260, uc_3261, uc_3262, uc_3263, uc_3264, uc_3265, uc_3266, uc_3267, 
      uc_3268, uc_3269, uc_3270, uc_3271, uc_3272, uc_3273, uc_3274, uc_3275, 
      uc_3276, uc_3277, uc_3278, uc_3279, uc_3280, uc_3281, normalizedWires[348], 
      \intermediateWiresStage1[2] [27], \intermediateWiresStage1[2] [26], 
      \intermediateWiresStage2[0] [25], \intermediateWiresStage2[0] [24], 
      \intermediateWiresStage2[0] [23], \intermediateWiresStage2[0] [22], 
      \intermediateWiresStage2[0] [21], \intermediateWiresStage2[0] [20], 
      \intermediateWiresStage2[0] [19], \intermediateWiresStage2[0] [18], 
      \intermediateWiresStage2[0] [17], \intermediateWiresStage2[0] [16], 
      \intermediateWiresStage2[0] [15], \intermediateWiresStage2[0] [14], 
      \intermediateWiresStage2[0] [13], \intermediateWiresStage2[0] [12], 
      \intermediateWiresStage2[0] [11], \intermediateWiresStage2[0] [10], 
      \intermediateWiresStage2[0] [9], \intermediateWiresStage2[0] [8], 
      \intermediateWiresStage2[0] [7], \intermediateWiresStage2[0] [6], 
      \intermediateWiresStage2[0] [5], \intermediateWiresStage2[0] [4], 
      \intermediateWiresStage2[0] [3], uc_3282, uc_3283, uc_3284}), .B({1'b0, 
      uc_3285, uc_3286, uc_3287, uc_3288, uc_3289, uc_3290, uc_3291, uc_3292, 
      uc_3293, uc_3294, uc_3295, uc_3296, uc_3297, uc_3298, uc_3299, uc_3300, 
      uc_3301, uc_3302, uc_3303, uc_3304, uc_3305, uc_3306, uc_3307, uc_3308, 
      uc_3309, uc_3310, uc_3311, uc_3312, uc_3313, uc_3314, uc_3315, uc_3316, 
      uc_3317, uc_3318, uc_3319, uc_3320, \intermediateWiresStage2[1] [26], 
      \intermediateWiresStage2[1] [25], \intermediateWiresStage2[1] [24], 
      \intermediateWiresStage2[1] [23], \intermediateWiresStage2[1] [22], 
      \intermediateWiresStage2[1] [21], \intermediateWiresStage2[1] [20], 
      \intermediateWiresStage2[1] [19], \intermediateWiresStage2[1] [18], 
      \intermediateWiresStage2[1] [17], \intermediateWiresStage2[1] [16], 
      \intermediateWiresStage2[1] [15], \intermediateWiresStage2[1] [14], 
      \intermediateWiresStage2[1] [13], \intermediateWiresStage2[1] [12], 
      \intermediateWiresStage2[1] [11], \intermediateWiresStage2[1] [10], 
      \intermediateWiresStage2[1] [9], \intermediateWiresStage2[1] [8], 
      \intermediateWiresStage2[1] [7], \intermediateWiresStage2[1] [6], 
      \intermediateWiresStage2[1] [5], \intermediateWiresStage2[1] [4], 
      \intermediateWiresStage2[1] [3], uc_3321, uc_3322, uc_3323}), .C({1'b0, 
      uc_3324, uc_3325, uc_3326, uc_3327, uc_3328, uc_3329, uc_3330, uc_3331, 
      uc_3332, uc_3333, uc_3334, uc_3335, uc_3336, uc_3337, uc_3338, uc_3339, 
      uc_3340, uc_3341, uc_3342, uc_3343, uc_3344, uc_3345, uc_3346, uc_3347, 
      uc_3348, uc_3349, uc_3350, uc_3351, uc_3352, uc_3353, uc_3354, uc_3355, 
      uc_3356, uc_3357, \intermediateWiresStage2[2] [28], 
      \intermediateWiresStage2[2] [27], \intermediateWiresStage2[2] [26], 
      \intermediateWiresStage2[2] [25], \intermediateWiresStage2[2] [24], 
      \intermediateWiresStage2[2] [23], \intermediateWiresStage2[2] [22], 
      \intermediateWiresStage2[2] [21], \intermediateWiresStage2[2] [20], 
      \intermediateWiresStage2[2] [19], \intermediateWiresStage2[2] [18], 
      \intermediateWiresStage2[2] [17], \intermediateWiresStage2[2] [16], 
      \intermediateWiresStage2[2] [15], \intermediateWiresStage2[2] [14], 
      \intermediateWiresStage2[2] [13], \intermediateWiresStage2[2] [12], 
      \intermediateWiresStage2[2] [11], \intermediateWiresStage2[2] [10], 
      \intermediateWiresStage2[2] [9], \intermediateWiresStage2[2] [8], 
      \intermediateWiresStage2[2] [7], \intermediateWiresStage2[2] [6], 
      \intermediateWiresStage1[3] [5], uc_3358, uc_3359, uc_3360, uc_3361, 
      uc_3362}));
   CSAlike__4_500 genblk5_2_parallelAdderStage4 (.result({uc_3363, uc_3364, 
      uc_3365, uc_3366, uc_3367, uc_3368, uc_3369, uc_3370, uc_3371, uc_3372, 
      uc_3373, uc_3374, uc_3375, uc_3376, uc_3377, uc_3378, uc_3379, uc_3380, 
      \intermediateWiresStage4[4] [45], \intermediateWiresStage4[4] [44], 
      \intermediateWiresStage4[4] [43], \intermediateWiresStage4[4] [42], 
      \intermediateWiresStage4[4] [41], \intermediateWiresStage4[4] [40], 
      \intermediateWiresStage4[4] [39], \intermediateWiresStage4[4] [38], 
      \intermediateWiresStage4[4] [37], \intermediateWiresStage4[4] [36], 
      \intermediateWiresStage4[4] [35], \intermediateWiresStage4[4] [34], 
      \intermediateWiresStage4[4] [33], \intermediateWiresStage4[4] [32], 
      \intermediateWiresStage4[4] [31], \intermediateWiresStage4[4] [30], 
      \intermediateWiresStage4[4] [29], \intermediateWiresStage4[4] [28], 
      \intermediateWiresStage4[4] [27], \intermediateWiresStage4[4] [26], 
      \intermediateWiresStage4[4] [25], \intermediateWiresStage4[4] [24], 
      uc_3381, uc_3382, uc_3383, uc_3384, uc_3385, uc_3386, uc_3387, uc_3388, 
      uc_3389, uc_3390, uc_3391, uc_3392, uc_3393, uc_3394, uc_3395, uc_3396, 
      uc_3397, uc_3398, uc_3399, uc_3400, uc_3401, uc_3402, uc_3403, uc_3404}), 
      .carry({uc_3405, uc_3406, uc_3407, uc_3408, uc_3409, uc_3410, uc_3411, 
      uc_3412, uc_3413, uc_3414, uc_3415, uc_3416, uc_3417, uc_3418, uc_3419, 
      uc_3420, uc_3421, \intermediateWiresStage4[5] [46], 
      \intermediateWiresStage4[5] [45], \intermediateWiresStage4[5] [44], 
      \intermediateWiresStage4[5] [43], \intermediateWiresStage4[5] [42], 
      \intermediateWiresStage4[5] [41], \intermediateWiresStage4[5] [40], 
      \intermediateWiresStage4[5] [39], \intermediateWiresStage4[5] [38], 
      \intermediateWiresStage4[5] [37], \intermediateWiresStage4[5] [36], 
      \intermediateWiresStage4[5] [35], \intermediateWiresStage4[5] [34], 
      \intermediateWiresStage4[5] [33], \intermediateWiresStage4[5] [32], 
      \intermediateWiresStage4[5] [31], \intermediateWiresStage4[5] [30], 
      \intermediateWiresStage4[5] [29], \intermediateWiresStage4[5] [28], 
      \intermediateWiresStage4[5] [27], \intermediateWiresStage4[5] [26], 
      \intermediateWiresStage4[5] [25], uc_3422, uc_3423, uc_3424, uc_3425, 
      uc_3426, uc_3427, uc_3428, uc_3429, uc_3430, uc_3431, uc_3432, uc_3433, 
      uc_3434, uc_3435, uc_3436, uc_3437, uc_3438, uc_3439, uc_3440, uc_3441, 
      uc_3442, uc_3443, uc_3444, uc_3445, uc_3446}), .A({1'b0, uc_3447, uc_3448, 
      uc_3449, uc_3450, uc_3451, uc_3452, uc_3453, uc_3454, uc_3455, uc_3456, 
      uc_3457, uc_3458, uc_3459, uc_3460, uc_3461, uc_3462, uc_3463, 
      \intermediateWiresStage1[15] [45], \intermediateWiresStage3[6] [44], 
      \intermediateWiresStage3[6] [43], \intermediateWiresStage3[6] [42], 
      \intermediateWiresStage3[6] [41], \intermediateWiresStage3[6] [40], 
      \intermediateWiresStage3[6] [39], \intermediateWiresStage3[6] [38], 
      \intermediateWiresStage3[6] [37], \intermediateWiresStage3[6] [36], 
      \intermediateWiresStage3[6] [35], \intermediateWiresStage3[6] [34], 
      \intermediateWiresStage3[6] [33], \intermediateWiresStage3[6] [32], 
      \intermediateWiresStage3[6] [31], \intermediateWiresStage3[6] [30], 
      \intermediateWiresStage3[6] [29], \intermediateWiresStage3[6] [28], 
      \intermediateWiresStage3[6] [27], \intermediateWiresStage3[6] [26], 
      \intermediateWiresStage3[6] [25], \intermediateWiresStage3[6] [24], 
      uc_3464, uc_3465, uc_3466, uc_3467, uc_3468, uc_3469, uc_3470, uc_3471, 
      uc_3472, uc_3473, uc_3474, uc_3475, uc_3476, uc_3477, uc_3478, uc_3479, 
      uc_3480, uc_3481, uc_3482, uc_3483, uc_3484, uc_3485, uc_3486, uc_3487}), 
      .B({1'b0, uc_3488, uc_3489, uc_3490, uc_3491, uc_3492, uc_3493, uc_3494, 
      uc_3495, uc_3496, uc_3497, uc_3498, uc_3499, uc_3500, uc_3501, uc_3502, 
      uc_3503, uc_3504, \intermediateWiresStage3[7] [45], 
      \intermediateWiresStage3[7] [44], \intermediateWiresStage3[7] [43], 
      \intermediateWiresStage3[7] [42], \intermediateWiresStage3[7] [41], 
      \intermediateWiresStage3[7] [40], \intermediateWiresStage3[7] [39], 
      \intermediateWiresStage3[7] [38], \intermediateWiresStage3[7] [37], 
      \intermediateWiresStage3[7] [36], \intermediateWiresStage3[7] [35], 
      \intermediateWiresStage3[7] [34], \intermediateWiresStage3[7] [33], 
      \intermediateWiresStage3[7] [32], \intermediateWiresStage3[7] [31], 
      \intermediateWiresStage3[7] [30], \intermediateWiresStage3[7] [29], 
      \intermediateWiresStage3[7] [28], \intermediateWiresStage3[7] [27], 
      \intermediateWiresStage3[7] [26], \intermediateWiresStage3[7] [25], 
      \intermediateWiresStage3[7] [24], uc_3505, uc_3506, uc_3507, uc_3508, 
      uc_3509, uc_3510, uc_3511, uc_3512, uc_3513, uc_3514, uc_3515, uc_3516, 
      uc_3517, uc_3518, uc_3519, uc_3520, uc_3521, uc_3522, uc_3523, uc_3524, 
      uc_3525, uc_3526, uc_3527, uc_3528}), .C({1'b0, uc_3529, uc_3530, uc_3531, 
      uc_3532, uc_3533, uc_3534, uc_3535, uc_3536, uc_3537, uc_3538, uc_3539, 
      uc_3540, uc_3541, uc_3542, uc_3543, uc_3544, uc_3545, uc_3546, uc_3547, 
      uc_3548, uc_3549, uc_3550, uc_3551, uc_3552, uc_3553, uc_3554, uc_3555, 
      uc_3556, uc_3557, uc_3558, uc_3559, uc_3560, uc_3561, uc_3562, uc_3563, 
      uc_3564, uc_3565, uc_3566, uc_3567, uc_3568, uc_3569, uc_3570, uc_3571, 
      uc_3572, uc_3573, uc_3574, uc_3575, uc_3576, uc_3577, uc_3578, uc_3579, 
      uc_3580, uc_3581, uc_3582, uc_3583, uc_3584, uc_3585, uc_3586, uc_3587, 
      uc_3588, uc_3589, uc_3590, uc_3591}));
   CSAlike__4_753 genblk5_1_parallelAdderStage4 (.result({uc_3592, uc_3593, 
      uc_3594, uc_3595, uc_3596, uc_3597, uc_3598, uc_3599, uc_3600, uc_3601, 
      uc_3602, uc_3603, uc_3604, uc_3605, uc_3606, uc_3607, uc_3608, uc_3609, 
      uc_3610, uc_3611, uc_3612, \intermediateWiresStage4[2] [42], 
      \intermediateWiresStage4[2] [41], \intermediateWiresStage4[2] [40], 
      \intermediateWiresStage4[2] [39], \intermediateWiresStage4[2] [38], 
      \intermediateWiresStage4[2] [37], \intermediateWiresStage4[2] [36], 
      \intermediateWiresStage4[2] [35], \intermediateWiresStage4[2] [34], 
      \intermediateWiresStage4[2] [33], \intermediateWiresStage4[2] [32], 
      \intermediateWiresStage4[2] [31], \intermediateWiresStage4[2] [30], 
      \intermediateWiresStage4[2] [29], \intermediateWiresStage4[2] [28], 
      \intermediateWiresStage4[2] [27], \intermediateWiresStage4[2] [26], 
      \intermediateWiresStage4[2] [25], \intermediateWiresStage4[2] [24], 
      \intermediateWiresStage4[2] [23], \intermediateWiresStage4[2] [22], 
      \intermediateWiresStage4[2] [21], \intermediateWiresStage4[2] [20], 
      \intermediateWiresStage4[2] [19], \intermediateWiresStage4[2] [18], 
      \intermediateWiresStage4[2] [17], \intermediateWiresStage4[2] [16], 
      \intermediateWiresStage4[2] [15], \intermediateWiresStage4[2] [14], 
      uc_3613, uc_3614, uc_3615, uc_3616, uc_3617, uc_3618, uc_3619, uc_3620, 
      uc_3621, uc_3622, uc_3623, uc_3624, uc_3625, uc_3626}), .carry({uc_3627, 
      uc_3628, uc_3629, uc_3630, uc_3631, uc_3632, uc_3633, uc_3634, uc_3635, 
      uc_3636, uc_3637, uc_3638, uc_3639, uc_3640, uc_3641, uc_3642, uc_3643, 
      uc_3644, uc_3645, uc_3646, \intermediateWiresStage4[3] [43], 
      \intermediateWiresStage4[3] [42], \intermediateWiresStage4[3] [41], 
      \intermediateWiresStage4[3] [40], \intermediateWiresStage4[3] [39], 
      \intermediateWiresStage4[3] [38], \intermediateWiresStage4[3] [37], 
      \intermediateWiresStage4[3] [36], \intermediateWiresStage4[3] [35], 
      \intermediateWiresStage4[3] [34], \intermediateWiresStage4[3] [33], 
      \intermediateWiresStage4[3] [32], \intermediateWiresStage4[3] [31], 
      \intermediateWiresStage4[3] [30], \intermediateWiresStage4[3] [29], 
      \intermediateWiresStage4[3] [28], \intermediateWiresStage4[3] [27], 
      \intermediateWiresStage4[3] [26], \intermediateWiresStage4[3] [25], 
      \intermediateWiresStage4[3] [24], \intermediateWiresStage4[3] [23], 
      \intermediateWiresStage4[3] [22], \intermediateWiresStage4[3] [21], 
      \intermediateWiresStage4[3] [20], \intermediateWiresStage4[3] [19], 
      \intermediateWiresStage4[3] [18], \intermediateWiresStage4[3] [17], 
      \intermediateWiresStage4[3] [16], \intermediateWiresStage4[3] [15], 
      uc_3647, uc_3648, uc_3649, uc_3650, uc_3651, uc_3652, uc_3653, uc_3654, 
      uc_3655, uc_3656, uc_3657, uc_3658, uc_3659, uc_3660, uc_3661}), .A({1'b0, 
      uc_3662, uc_3663, uc_3664, uc_3665, uc_3666, uc_3667, uc_3668, uc_3669, 
      uc_3670, uc_3671, uc_3672, uc_3673, uc_3674, uc_3675, uc_3676, uc_3677, 
      uc_3678, uc_3679, uc_3680, uc_3681, uc_3682, uc_3683, uc_3684, uc_3685, 
      uc_3686, uc_3687, \intermediateWiresStage3[3] [36], 
      \intermediateWiresStage3[3] [35], \intermediateWiresStage3[3] [34], 
      \intermediateWiresStage3[3] [33], \intermediateWiresStage3[3] [32], 
      \intermediateWiresStage3[3] [31], \intermediateWiresStage3[3] [30], 
      \intermediateWiresStage3[3] [29], \intermediateWiresStage3[3] [28], 
      \intermediateWiresStage3[3] [27], \intermediateWiresStage3[3] [26], 
      \intermediateWiresStage3[3] [25], \intermediateWiresStage3[3] [24], 
      \intermediateWiresStage3[3] [23], \intermediateWiresStage3[3] [22], 
      \intermediateWiresStage3[3] [21], \intermediateWiresStage3[3] [20], 
      \intermediateWiresStage3[3] [19], \intermediateWiresStage3[3] [18], 
      \intermediateWiresStage3[3] [17], \intermediateWiresStage3[3] [16], 
      \intermediateWiresStage3[3] [15], \intermediateWiresStage3[3] [14], 
      uc_3688, uc_3689, uc_3690, uc_3691, uc_3692, uc_3693, uc_3694, uc_3695, 
      uc_3696, uc_3697, uc_3698, uc_3699, uc_3700, uc_3701}), .B({1'b0, uc_3702, 
      uc_3703, uc_3704, uc_3705, uc_3706, uc_3707, uc_3708, uc_3709, uc_3710, 
      uc_3711, uc_3712, uc_3713, uc_3714, uc_3715, uc_3716, uc_3717, uc_3718, 
      uc_3719, uc_3720, uc_3721, \intermediateWiresStage2[8] [42], 
      \intermediateWiresStage3[4] [41], \intermediateWiresStage3[4] [40], 
      \intermediateWiresStage3[4] [39], \intermediateWiresStage3[4] [38], 
      \intermediateWiresStage3[4] [37], \intermediateWiresStage3[4] [36], 
      \intermediateWiresStage3[4] [35], \intermediateWiresStage3[4] [34], 
      \intermediateWiresStage3[4] [33], \intermediateWiresStage3[4] [32], 
      \intermediateWiresStage3[4] [31], \intermediateWiresStage3[4] [30], 
      \intermediateWiresStage3[4] [29], \intermediateWiresStage3[4] [28], 
      \intermediateWiresStage3[4] [27], \intermediateWiresStage3[4] [26], 
      \intermediateWiresStage3[4] [25], \intermediateWiresStage3[4] [24], 
      \intermediateWiresStage3[4] [23], \intermediateWiresStage3[4] [22], 
      \intermediateWiresStage3[4] [21], \intermediateWiresStage3[4] [20], 
      \intermediateWiresStage3[4] [19], \intermediateWiresStage3[4] [18], 
      \intermediateWiresStage3[4] [17], \intermediateWiresStage3[4] [16], 
      \intermediateWiresStage2[6] [15], \intermediateWiresStage1[9] [14], 
      uc_3722, uc_3723, uc_3724, uc_3725, uc_3726, uc_3727, uc_3728, uc_3729, 
      uc_3730, uc_3731, uc_3732, uc_3733, uc_3734, uc_3735}), .C({1'b0, uc_3736, 
      uc_3737, uc_3738, uc_3739, uc_3740, uc_3741, uc_3742, uc_3743, uc_3744, 
      uc_3745, uc_3746, uc_3747, uc_3748, uc_3749, uc_3750, uc_3751, uc_3752, 
      uc_3753, uc_3754, uc_3755, \intermediateWiresStage3[5] [42], 
      \intermediateWiresStage3[5] [41], \intermediateWiresStage3[5] [40], 
      \intermediateWiresStage3[5] [39], \intermediateWiresStage3[5] [38], 
      \intermediateWiresStage3[5] [37], \intermediateWiresStage3[5] [36], 
      \intermediateWiresStage3[5] [35], \intermediateWiresStage3[5] [34], 
      \intermediateWiresStage3[5] [33], \intermediateWiresStage3[5] [32], 
      \intermediateWiresStage3[5] [31], \intermediateWiresStage3[5] [30], 
      \intermediateWiresStage3[5] [29], \intermediateWiresStage3[5] [28], 
      \intermediateWiresStage3[5] [27], \intermediateWiresStage3[5] [26], 
      \intermediateWiresStage3[5] [25], \intermediateWiresStage3[5] [24], 
      \intermediateWiresStage3[5] [23], \intermediateWiresStage3[5] [22], 
      \intermediateWiresStage3[5] [21], \intermediateWiresStage3[5] [20], 
      \intermediateWiresStage3[5] [19], \intermediateWiresStage3[5] [18], 
      \intermediateWiresStage3[5] [17], uc_3756, uc_3757, uc_3758, uc_3759, 
      uc_3760, uc_3761, uc_3762, uc_3763, uc_3764, uc_3765, uc_3766, uc_3767, 
      uc_3768, uc_3769, uc_3770, uc_3771, uc_3772}));
   CSAlike__4_1006 genblk5_0_parallelAdderStage4 (.result({uc_3773, uc_3774, 
      uc_3775, uc_3776, uc_3777, uc_3778, uc_3779, uc_3780, uc_3781, uc_3782, 
      uc_3783, uc_3784, uc_3785, uc_3786, uc_3787, uc_3788, uc_3789, uc_3790, 
      uc_3791, uc_3792, uc_3793, uc_3794, uc_3795, uc_3796, uc_3797, uc_3798, 
      uc_3799, uc_3800, uc_3801, uc_3802, uc_3803, uc_3804, 
      \intermediateWiresStage4[0] [31], \intermediateWiresStage4[0] [30], 
      \intermediateWiresStage4[0] [29], \intermediateWiresStage4[0] [28], 
      \intermediateWiresStage4[0] [27], \intermediateWiresStage4[0] [26], 
      \intermediateWiresStage4[0] [25], \intermediateWiresStage4[0] [24], 
      \intermediateWiresStage4[0] [23], \intermediateWiresStage4[0] [22], 
      \intermediateWiresStage4[0] [21], \intermediateWiresStage4[0] [20], 
      \intermediateWiresStage4[0] [19], \intermediateWiresStage4[0] [18], 
      \intermediateWiresStage4[0] [17], \intermediateWiresStage4[0] [16], 
      \intermediateWiresStage4[0] [15], \intermediateWiresStage4[0] [14], 
      \intermediateWiresStage4[0] [13], \intermediateWiresStage4[0] [12], 
      \intermediateWiresStage4[0] [11], \intermediateWiresStage4[0] [10], 
      \intermediateWiresStage4[0] [9], \intermediateWiresStage4[0] [8], 
      \intermediateWiresStage4[0] [7], \intermediateWiresStage4[0] [6], 
      \intermediateWiresStage4[0] [5], uc_3805, uc_3806, uc_3807, uc_3808, 
      uc_3809}), .carry({uc_3810, uc_3811, uc_3812, uc_3813, uc_3814, uc_3815, 
      uc_3816, uc_3817, uc_3818, uc_3819, uc_3820, uc_3821, uc_3822, uc_3823, 
      uc_3824, uc_3825, uc_3826, uc_3827, uc_3828, uc_3829, uc_3830, uc_3831, 
      uc_3832, uc_3833, uc_3834, uc_3835, uc_3836, uc_3837, uc_3838, uc_3839, 
      uc_3840, \intermediateWiresStage4[1] [32], 
      \intermediateWiresStage4[1] [31], \intermediateWiresStage4[1] [30], 
      \intermediateWiresStage4[1] [29], \intermediateWiresStage4[1] [28], 
      \intermediateWiresStage4[1] [27], \intermediateWiresStage4[1] [26], 
      \intermediateWiresStage4[1] [25], \intermediateWiresStage4[1] [24], 
      \intermediateWiresStage4[1] [23], \intermediateWiresStage4[1] [22], 
      \intermediateWiresStage4[1] [21], \intermediateWiresStage4[1] [20], 
      \intermediateWiresStage4[1] [19], \intermediateWiresStage4[1] [18], 
      \intermediateWiresStage4[1] [17], \intermediateWiresStage4[1] [16], 
      \intermediateWiresStage4[1] [15], \intermediateWiresStage4[1] [14], 
      \intermediateWiresStage4[1] [13], \intermediateWiresStage4[1] [12], 
      \intermediateWiresStage4[1] [11], \intermediateWiresStage4[1] [10], 
      \intermediateWiresStage4[1] [9], \intermediateWiresStage4[1] [8], 
      \intermediateWiresStage4[1] [7], \intermediateWiresStage4[1] [6], 
      \intermediateWiresStage4[1] [5], uc_3841, uc_3842, uc_3843, uc_3844, 
      uc_3845}), .A({1'b0, uc_3846, uc_3847, uc_3848, uc_3849, uc_3850, uc_3851, 
      uc_3852, uc_3853, uc_3854, uc_3855, uc_3856, uc_3857, uc_3858, uc_3859, 
      uc_3860, uc_3861, uc_3862, uc_3863, uc_3864, uc_3865, uc_3866, uc_3867, 
      uc_3868, uc_3869, uc_3870, uc_3871, uc_3872, uc_3873, uc_3874, uc_3875, 
      uc_3876, \intermediateWiresStage2[2] [31], 
      \intermediateWiresStage2[2] [30], \intermediateWiresStage2[2] [29], 
      \intermediateWiresStage3[0] [28], \intermediateWiresStage3[0] [27], 
      \intermediateWiresStage3[0] [26], \intermediateWiresStage3[0] [25], 
      \intermediateWiresStage3[0] [24], \intermediateWiresStage3[0] [23], 
      \intermediateWiresStage3[0] [22], \intermediateWiresStage3[0] [21], 
      \intermediateWiresStage3[0] [20], \intermediateWiresStage3[0] [19], 
      \intermediateWiresStage3[0] [18], \intermediateWiresStage3[0] [17], 
      \intermediateWiresStage3[0] [16], \intermediateWiresStage3[0] [15], 
      \intermediateWiresStage3[0] [14], \intermediateWiresStage3[0] [13], 
      \intermediateWiresStage3[0] [12], \intermediateWiresStage3[0] [11], 
      \intermediateWiresStage3[0] [10], \intermediateWiresStage3[0] [9], 
      \intermediateWiresStage3[0] [8], \intermediateWiresStage3[0] [7], 
      \intermediateWiresStage3[0] [6], \intermediateWiresStage3[0] [5], 
      \intermediateWiresStage3[0] [4], uc_3877, uc_3878, uc_3879, uc_3880}), 
      .B({1'b0, uc_3881, uc_3882, uc_3883, uc_3884, uc_3885, uc_3886, uc_3887, 
      uc_3888, uc_3889, uc_3890, uc_3891, uc_3892, uc_3893, uc_3894, uc_3895, 
      uc_3896, uc_3897, uc_3898, uc_3899, uc_3900, uc_3901, uc_3902, uc_3903, 
      uc_3904, uc_3905, uc_3906, uc_3907, uc_3908, uc_3909, uc_3910, uc_3911, 
      uc_3912, uc_3913, \intermediateWiresStage3[1] [29], 
      \intermediateWiresStage3[1] [28], \intermediateWiresStage3[1] [27], 
      \intermediateWiresStage3[1] [26], \intermediateWiresStage3[1] [25], 
      \intermediateWiresStage3[1] [24], \intermediateWiresStage3[1] [23], 
      \intermediateWiresStage3[1] [22], \intermediateWiresStage3[1] [21], 
      \intermediateWiresStage3[1] [20], \intermediateWiresStage3[1] [19], 
      \intermediateWiresStage3[1] [18], \intermediateWiresStage3[1] [17], 
      \intermediateWiresStage3[1] [16], \intermediateWiresStage3[1] [15], 
      \intermediateWiresStage3[1] [14], \intermediateWiresStage3[1] [13], 
      \intermediateWiresStage3[1] [12], \intermediateWiresStage3[1] [11], 
      \intermediateWiresStage3[1] [10], \intermediateWiresStage3[1] [9], 
      \intermediateWiresStage3[1] [8], \intermediateWiresStage3[1] [7], 
      \intermediateWiresStage3[1] [6], \intermediateWiresStage3[1] [5], 
      \intermediateWiresStage3[1] [4], uc_3914, uc_3915, uc_3916, uc_3917}), 
      .C({1'b0, uc_3918, uc_3919, uc_3920, uc_3921, uc_3922, uc_3923, uc_3924, 
      uc_3925, uc_3926, uc_3927, uc_3928, uc_3929, uc_3930, uc_3931, uc_3932, 
      uc_3933, uc_3934, uc_3935, uc_3936, uc_3937, uc_3938, uc_3939, uc_3940, 
      uc_3941, uc_3942, uc_3943, uc_3944, uc_3945, uc_3946, uc_3947, uc_3948, 
      \intermediateWiresStage3[2] [31], \intermediateWiresStage3[2] [30], 
      \intermediateWiresStage3[2] [29], \intermediateWiresStage3[2] [28], 
      \intermediateWiresStage3[2] [27], \intermediateWiresStage3[2] [26], 
      \intermediateWiresStage3[2] [25], \intermediateWiresStage3[2] [24], 
      \intermediateWiresStage3[2] [23], \intermediateWiresStage3[2] [22], 
      \intermediateWiresStage3[2] [21], \intermediateWiresStage3[2] [20], 
      \intermediateWiresStage3[2] [19], \intermediateWiresStage3[2] [18], 
      \intermediateWiresStage3[2] [17], \intermediateWiresStage3[2] [16], 
      \intermediateWiresStage3[2] [15], \intermediateWiresStage3[2] [14], 
      \intermediateWiresStage3[2] [13], \intermediateWiresStage3[2] [12], 
      \intermediateWiresStage3[2] [11], \intermediateWiresStage3[2] [10], 
      \intermediateWiresStage3[2] [9], \intermediateWiresStage2[3] [8], 
      \intermediateWiresStage2[3] [7], uc_3949, uc_3950, uc_3951, uc_3952, 
      uc_3953, uc_3954, uc_3955}));
   CSAlike__4_1259 genblk6_1_parallelAdderStage5 (.result({uc_3956, uc_3957, 
      uc_3958, uc_3959, uc_3960, uc_3961, uc_3962, uc_3963, uc_3964, uc_3965, 
      uc_3966, uc_3967, uc_3968, uc_3969, uc_3970, uc_3971, uc_3972, 
      \intermediateWiresStage5[2] [46], \intermediateWiresStage5[2] [45], 
      \intermediateWiresStage5[2] [44], \intermediateWiresStage5[2] [43], 
      \intermediateWiresStage5[2] [42], \intermediateWiresStage5[2] [41], 
      \intermediateWiresStage5[2] [40], \intermediateWiresStage5[2] [39], 
      \intermediateWiresStage5[2] [38], \intermediateWiresStage5[2] [37], 
      \intermediateWiresStage5[2] [36], \intermediateWiresStage5[2] [35], 
      \intermediateWiresStage5[2] [34], \intermediateWiresStage5[2] [33], 
      \intermediateWiresStage5[2] [32], \intermediateWiresStage5[2] [31], 
      \intermediateWiresStage5[2] [30], \intermediateWiresStage5[2] [29], 
      \intermediateWiresStage5[2] [28], \intermediateWiresStage5[2] [27], 
      \intermediateWiresStage5[2] [26], \intermediateWiresStage5[2] [25], 
      \intermediateWiresStage5[2] [24], \intermediateWiresStage5[2] [23], 
      \intermediateWiresStage5[2] [22], \intermediateWiresStage5[2] [21], 
      uc_3973, uc_3974, uc_3975, uc_3976, uc_3977, uc_3978, uc_3979, uc_3980, 
      uc_3981, uc_3982, uc_3983, uc_3984, uc_3985, uc_3986, uc_3987, uc_3988, 
      uc_3989, uc_3990, uc_3991, uc_3992, uc_3993}), .carry({uc_3994, uc_3995, 
      uc_3996, uc_3997, uc_3998, uc_3999, uc_4000, uc_4001, uc_4002, uc_4003, 
      uc_4004, uc_4005, uc_4006, uc_4007, uc_4008, uc_4009, 
      \intermediateWiresStage5[3] [47], \intermediateWiresStage5[3] [46], 
      \intermediateWiresStage5[3] [45], \intermediateWiresStage5[3] [44], 
      \intermediateWiresStage5[3] [43], \intermediateWiresStage5[3] [42], 
      \intermediateWiresStage5[3] [41], \intermediateWiresStage5[3] [40], 
      \intermediateWiresStage5[3] [39], \intermediateWiresStage5[3] [38], 
      \intermediateWiresStage5[3] [37], \intermediateWiresStage5[3] [36], 
      \intermediateWiresStage5[3] [35], \intermediateWiresStage5[3] [34], 
      \intermediateWiresStage5[3] [33], \intermediateWiresStage5[3] [32], 
      \intermediateWiresStage5[3] [31], \intermediateWiresStage5[3] [30], 
      \intermediateWiresStage5[3] [29], \intermediateWiresStage5[3] [28], 
      \intermediateWiresStage5[3] [27], \intermediateWiresStage5[3] [26], 
      \intermediateWiresStage5[3] [25], \intermediateWiresStage5[3] [24], 
      \intermediateWiresStage5[3] [23], \intermediateWiresStage5[3] [22], 
      uc_4010, uc_4011, uc_4012, uc_4013, uc_4014, uc_4015, uc_4016, uc_4017, 
      uc_4018, uc_4019, uc_4020, uc_4021, uc_4022, uc_4023, uc_4024, uc_4025, 
      uc_4026, uc_4027, uc_4028, uc_4029, uc_4030, uc_4031}), .A({1'b0, uc_4032, 
      uc_4033, uc_4034, uc_4035, uc_4036, uc_4037, uc_4038, uc_4039, uc_4040, 
      uc_4041, uc_4042, uc_4043, uc_4044, uc_4045, uc_4046, uc_4047, uc_4048, 
      uc_4049, uc_4050, \intermediateWiresStage4[3] [43], 
      \intermediateWiresStage4[3] [42], \intermediateWiresStage4[3] [41], 
      \intermediateWiresStage4[3] [40], \intermediateWiresStage4[3] [39], 
      \intermediateWiresStage4[3] [38], \intermediateWiresStage4[3] [37], 
      \intermediateWiresStage4[3] [36], \intermediateWiresStage4[3] [35], 
      \intermediateWiresStage4[3] [34], \intermediateWiresStage4[3] [33], 
      \intermediateWiresStage4[3] [32], \intermediateWiresStage4[3] [31], 
      \intermediateWiresStage4[3] [30], \intermediateWiresStage4[3] [29], 
      \intermediateWiresStage4[3] [28], \intermediateWiresStage4[3] [27], 
      \intermediateWiresStage4[3] [26], \intermediateWiresStage4[3] [25], 
      \intermediateWiresStage4[3] [24], \intermediateWiresStage4[3] [23], 
      \intermediateWiresStage4[3] [22], \intermediateWiresStage4[3] [21], 
      uc_4051, uc_4052, uc_4053, uc_4054, uc_4055, uc_4056, uc_4057, uc_4058, 
      uc_4059, uc_4060, uc_4061, uc_4062, uc_4063, uc_4064, uc_4065, uc_4066, 
      uc_4067, uc_4068, uc_4069, uc_4070, uc_4071}), .B({1'b0, uc_4072, uc_4073, 
      uc_4074, uc_4075, uc_4076, uc_4077, uc_4078, uc_4079, uc_4080, uc_4081, 
      uc_4082, uc_4083, uc_4084, uc_4085, uc_4086, uc_4087, 
      \intermediateWiresStage1[15] [46], \intermediateWiresStage4[4] [45], 
      \intermediateWiresStage4[4] [44], \intermediateWiresStage4[4] [43], 
      \intermediateWiresStage4[4] [42], \intermediateWiresStage4[4] [41], 
      \intermediateWiresStage4[4] [40], \intermediateWiresStage4[4] [39], 
      \intermediateWiresStage4[4] [38], \intermediateWiresStage4[4] [37], 
      \intermediateWiresStage4[4] [36], \intermediateWiresStage4[4] [35], 
      \intermediateWiresStage4[4] [34], \intermediateWiresStage4[4] [33], 
      \intermediateWiresStage4[4] [32], \intermediateWiresStage4[4] [31], 
      \intermediateWiresStage4[4] [30], \intermediateWiresStage4[4] [29], 
      \intermediateWiresStage4[4] [28], \intermediateWiresStage4[4] [27], 
      \intermediateWiresStage4[4] [26], \intermediateWiresStage4[4] [25], 
      \intermediateWiresStage4[4] [24], \intermediateWiresStage3[6] [23], 
      \intermediateWiresStage2[9] [22], \intermediateWiresStage2[9] [21], 
      uc_4088, uc_4089, uc_4090, uc_4091, uc_4092, uc_4093, uc_4094, uc_4095, 
      uc_4096, uc_4097, uc_4098, uc_4099, uc_4100, uc_4101, uc_4102, uc_4103, 
      uc_4104, uc_4105, uc_4106, uc_4107, uc_4108}), .C({1'b0, uc_4109, uc_4110, 
      uc_4111, uc_4112, uc_4113, uc_4114, uc_4115, uc_4116, uc_4117, uc_4118, 
      uc_4119, uc_4120, uc_4121, uc_4122, uc_4123, uc_4124, 
      \intermediateWiresStage4[5] [46], \intermediateWiresStage4[5] [45], 
      \intermediateWiresStage4[5] [44], \intermediateWiresStage4[5] [43], 
      \intermediateWiresStage4[5] [42], \intermediateWiresStage4[5] [41], 
      \intermediateWiresStage4[5] [40], \intermediateWiresStage4[5] [39], 
      \intermediateWiresStage4[5] [38], \intermediateWiresStage4[5] [37], 
      \intermediateWiresStage4[5] [36], \intermediateWiresStage4[5] [35], 
      \intermediateWiresStage4[5] [34], \intermediateWiresStage4[5] [33], 
      \intermediateWiresStage4[5] [32], \intermediateWiresStage4[5] [31], 
      \intermediateWiresStage4[5] [30], \intermediateWiresStage4[5] [29], 
      \intermediateWiresStage4[5] [28], \intermediateWiresStage4[5] [27], 
      \intermediateWiresStage4[5] [26], \intermediateWiresStage4[5] [25], 
      uc_4125, uc_4126, uc_4127, uc_4128, uc_4129, uc_4130, uc_4131, uc_4132, 
      uc_4133, uc_4134, uc_4135, uc_4136, uc_4137, uc_4138, uc_4139, uc_4140, 
      uc_4141, uc_4142, uc_4143, uc_4144, uc_4145, uc_4146, uc_4147, uc_4148, 
      uc_4149}));
   CSAlike__4_1512 genblk6_0_parallelAdderStage5 (.result({uc_4150, uc_4151, 
      uc_4152, uc_4153, uc_4154, uc_4155, uc_4156, uc_4157, uc_4158, uc_4159, 
      uc_4160, uc_4161, uc_4162, uc_4163, uc_4164, uc_4165, uc_4166, uc_4167, 
      uc_4168, uc_4169, uc_4170, uc_4171, uc_4172, uc_4173, uc_4174, uc_4175, 
      \intermediateWiresStage5[0] [37], \intermediateWiresStage5[0] [36], 
      \intermediateWiresStage5[0] [35], \intermediateWiresStage5[0] [34], 
      \intermediateWiresStage5[0] [33], \intermediateWiresStage5[0] [32], 
      \intermediateWiresStage5[0] [31], \intermediateWiresStage5[0] [30], 
      \intermediateWiresStage5[0] [29], \intermediateWiresStage5[0] [28], 
      \intermediateWiresStage5[0] [27], \intermediateWiresStage5[0] [26], 
      \intermediateWiresStage5[0] [25], \intermediateWiresStage5[0] [24], 
      \intermediateWiresStage5[0] [23], \intermediateWiresStage5[0] [22], 
      \intermediateWiresStage5[0] [21], \intermediateWiresStage5[0] [20], 
      \intermediateWiresStage5[0] [19], \intermediateWiresStage5[0] [18], 
      \intermediateWiresStage5[0] [17], \intermediateWiresStage5[0] [16], 
      \intermediateWiresStage5[0] [15], \intermediateWiresStage5[0] [14], 
      \intermediateWiresStage5[0] [13], \intermediateWiresStage5[0] [12], 
      \intermediateWiresStage5[0] [11], \intermediateWiresStage5[0] [10], 
      \intermediateWiresStage5[0] [9], \intermediateWiresStage5[0] [8], 
      \intermediateWiresStage5[0] [7], \intermediateWiresStage5[0] [6], uc_4176, 
      uc_4177, uc_4178, uc_4179, uc_4180, uc_4181}), .carry({uc_4182, uc_4183, 
      uc_4184, uc_4185, uc_4186, uc_4187, uc_4188, uc_4189, uc_4190, uc_4191, 
      uc_4192, uc_4193, uc_4194, uc_4195, uc_4196, uc_4197, uc_4198, uc_4199, 
      uc_4200, uc_4201, uc_4202, uc_4203, uc_4204, uc_4205, uc_4206, 
      \intermediateWiresStage5[1] [38], \intermediateWiresStage5[1] [37], 
      \intermediateWiresStage5[1] [36], \intermediateWiresStage5[1] [35], 
      \intermediateWiresStage5[1] [34], \intermediateWiresStage5[1] [33], 
      \intermediateWiresStage5[1] [32], \intermediateWiresStage5[1] [31], 
      \intermediateWiresStage5[1] [30], \intermediateWiresStage5[1] [29], 
      \intermediateWiresStage5[1] [28], \intermediateWiresStage5[1] [27], 
      \intermediateWiresStage5[1] [26], \intermediateWiresStage5[1] [25], 
      \intermediateWiresStage5[1] [24], \intermediateWiresStage5[1] [23], 
      \intermediateWiresStage5[1] [22], \intermediateWiresStage5[1] [21], 
      \intermediateWiresStage5[1] [20], \intermediateWiresStage5[1] [19], 
      \intermediateWiresStage5[1] [18], \intermediateWiresStage5[1] [17], 
      \intermediateWiresStage5[1] [16], \intermediateWiresStage5[1] [15], 
      \intermediateWiresStage5[1] [14], \intermediateWiresStage5[1] [13], 
      \intermediateWiresStage5[1] [12], \intermediateWiresStage5[1] [11], 
      \intermediateWiresStage5[1] [10], \intermediateWiresStage5[1] [9], 
      \intermediateWiresStage5[1] [8], \intermediateWiresStage5[1] [7], 
      \intermediateWiresStage5[1] [6], uc_4207, uc_4208, uc_4209, uc_4210, 
      uc_4211, uc_4212}), .A({1'b0, uc_4213, uc_4214, uc_4215, uc_4216, uc_4217, 
      uc_4218, uc_4219, uc_4220, uc_4221, uc_4222, uc_4223, uc_4224, uc_4225, 
      uc_4226, uc_4227, uc_4228, uc_4229, uc_4230, uc_4231, uc_4232, uc_4233, 
      uc_4234, uc_4235, uc_4236, uc_4237, normalizedWires[933], 
      \intermediateWiresStage1[8] [36], \intermediateWiresStage3[2] [35], 
      \intermediateWiresStage3[2] [34], \intermediateWiresStage3[2] [33], 
      \intermediateWiresStage3[2] [32], \intermediateWiresStage4[0] [31], 
      \intermediateWiresStage4[0] [30], \intermediateWiresStage4[0] [29], 
      \intermediateWiresStage4[0] [28], \intermediateWiresStage4[0] [27], 
      \intermediateWiresStage4[0] [26], \intermediateWiresStage4[0] [25], 
      \intermediateWiresStage4[0] [24], \intermediateWiresStage4[0] [23], 
      \intermediateWiresStage4[0] [22], \intermediateWiresStage4[0] [21], 
      \intermediateWiresStage4[0] [20], \intermediateWiresStage4[0] [19], 
      \intermediateWiresStage4[0] [18], \intermediateWiresStage4[0] [17], 
      \intermediateWiresStage4[0] [16], \intermediateWiresStage4[0] [15], 
      \intermediateWiresStage4[0] [14], \intermediateWiresStage4[0] [13], 
      \intermediateWiresStage4[0] [12], \intermediateWiresStage4[0] [11], 
      \intermediateWiresStage4[0] [10], \intermediateWiresStage4[0] [9], 
      \intermediateWiresStage4[0] [8], \intermediateWiresStage4[0] [7], 
      \intermediateWiresStage4[0] [6], \intermediateWiresStage4[0] [5], uc_4238, 
      uc_4239, uc_4240, uc_4241, uc_4242}), .B({1'b0, uc_4243, uc_4244, uc_4245, 
      uc_4246, uc_4247, uc_4248, uc_4249, uc_4250, uc_4251, uc_4252, uc_4253, 
      uc_4254, uc_4255, uc_4256, uc_4257, uc_4258, uc_4259, uc_4260, uc_4261, 
      uc_4262, uc_4263, uc_4264, uc_4265, uc_4266, uc_4267, uc_4268, uc_4269, 
      uc_4270, uc_4271, uc_4272, \intermediateWiresStage4[1] [32], 
      \intermediateWiresStage4[1] [31], \intermediateWiresStage4[1] [30], 
      \intermediateWiresStage4[1] [29], \intermediateWiresStage4[1] [28], 
      \intermediateWiresStage4[1] [27], \intermediateWiresStage4[1] [26], 
      \intermediateWiresStage4[1] [25], \intermediateWiresStage4[1] [24], 
      \intermediateWiresStage4[1] [23], \intermediateWiresStage4[1] [22], 
      \intermediateWiresStage4[1] [21], \intermediateWiresStage4[1] [20], 
      \intermediateWiresStage4[1] [19], \intermediateWiresStage4[1] [18], 
      \intermediateWiresStage4[1] [17], \intermediateWiresStage4[1] [16], 
      \intermediateWiresStage4[1] [15], \intermediateWiresStage4[1] [14], 
      \intermediateWiresStage4[1] [13], \intermediateWiresStage4[1] [12], 
      \intermediateWiresStage4[1] [11], \intermediateWiresStage4[1] [10], 
      \intermediateWiresStage4[1] [9], \intermediateWiresStage4[1] [8], 
      \intermediateWiresStage4[1] [7], \intermediateWiresStage4[1] [6], 
      \intermediateWiresStage4[1] [5], uc_4273, uc_4274, uc_4275, uc_4276, 
      uc_4277}), .C({1'b0, uc_4278, uc_4279, uc_4280, uc_4281, uc_4282, uc_4283, 
      uc_4284, uc_4285, uc_4286, uc_4287, uc_4288, uc_4289, uc_4290, uc_4291, 
      uc_4292, uc_4293, uc_4294, uc_4295, uc_4296, uc_4297, uc_4298, uc_4299, 
      uc_4300, uc_4301, uc_4302, \intermediateWiresStage4[2] [37], 
      \intermediateWiresStage4[2] [36], \intermediateWiresStage4[2] [35], 
      \intermediateWiresStage4[2] [34], \intermediateWiresStage4[2] [33], 
      \intermediateWiresStage4[2] [32], \intermediateWiresStage4[2] [31], 
      \intermediateWiresStage4[2] [30], \intermediateWiresStage4[2] [29], 
      \intermediateWiresStage4[2] [28], \intermediateWiresStage4[2] [27], 
      \intermediateWiresStage4[2] [26], \intermediateWiresStage4[2] [25], 
      \intermediateWiresStage4[2] [24], \intermediateWiresStage4[2] [23], 
      \intermediateWiresStage4[2] [22], \intermediateWiresStage4[2] [21], 
      \intermediateWiresStage4[2] [20], \intermediateWiresStage4[2] [19], 
      \intermediateWiresStage4[2] [18], \intermediateWiresStage4[2] [17], 
      \intermediateWiresStage4[2] [16], \intermediateWiresStage4[2] [15], 
      \intermediateWiresStage4[2] [14], \intermediateWiresStage3[3] [13], 
      \intermediateWiresStage3[3] [12], \intermediateWiresStage3[3] [11], 
      \intermediateWiresStage3[3] [10], uc_4303, uc_4304, uc_4305, uc_4306, 
      uc_4307, uc_4308, uc_4309, uc_4310, uc_4311, uc_4312}));
   CSAlike__4_1765 genblk7_0_parallelAdderStage6 (.result({uc_4313, uc_4314, 
      uc_4315, uc_4316, uc_4317, uc_4318, uc_4319, uc_4320, uc_4321, uc_4322, 
      uc_4323, uc_4324, uc_4325, uc_4326, uc_4327, uc_4328, uc_4329, 
      \intermediateWiresStage6[0] [46], \intermediateWiresStage6[0] [45], 
      \intermediateWiresStage6[0] [44], \intermediateWiresStage6[0] [43], 
      \intermediateWiresStage6[0] [42], \intermediateWiresStage6[0] [41], 
      \intermediateWiresStage6[0] [40], \intermediateWiresStage6[0] [39], 
      \intermediateWiresStage6[0] [38], \intermediateWiresStage6[0] [37], 
      \intermediateWiresStage6[0] [36], \intermediateWiresStage6[0] [35], 
      \intermediateWiresStage6[0] [34], \intermediateWiresStage6[0] [33], 
      \intermediateWiresStage6[0] [32], \intermediateWiresStage6[0] [31], 
      \intermediateWiresStage6[0] [30], \intermediateWiresStage6[0] [29], 
      \intermediateWiresStage6[0] [28], \intermediateWiresStage6[0] [27], 
      \intermediateWiresStage6[0] [26], \intermediateWiresStage6[0] [25], 
      \intermediateWiresStage6[0] [24], \intermediateWiresStage6[0] [23], 
      \intermediateWiresStage6[0] [22], \intermediateWiresStage6[0] [21], 
      \intermediateWiresStage6[0] [20], \intermediateWiresStage6[0] [19], 
      \intermediateWiresStage6[0] [18], \intermediateWiresStage6[0] [17], 
      \intermediateWiresStage6[0] [16], \intermediateWiresStage6[0] [15], 
      \intermediateWiresStage6[0] [14], \intermediateWiresStage6[0] [13], 
      \intermediateWiresStage6[0] [12], \intermediateWiresStage6[0] [11], 
      \intermediateWiresStage6[0] [10], \intermediateWiresStage6[0] [9], 
      \intermediateWiresStage6[0] [8], \intermediateWiresStage6[0] [7], uc_4330, 
      uc_4331, uc_4332, uc_4333, uc_4334, uc_4335, uc_4336}), .carry({uc_4337, 
      uc_4338, uc_4339, uc_4340, uc_4341, uc_4342, uc_4343, uc_4344, uc_4345, 
      uc_4346, uc_4347, uc_4348, uc_4349, uc_4350, uc_4351, uc_4352, 
      \intermediateWiresStage6[1] [47], \intermediateWiresStage6[1] [46], 
      \intermediateWiresStage6[1] [45], \intermediateWiresStage6[1] [44], 
      \intermediateWiresStage6[1] [43], \intermediateWiresStage6[1] [42], 
      \intermediateWiresStage6[1] [41], \intermediateWiresStage6[1] [40], 
      \intermediateWiresStage6[1] [39], \intermediateWiresStage6[1] [38], 
      \intermediateWiresStage6[1] [37], \intermediateWiresStage6[1] [36], 
      \intermediateWiresStage6[1] [35], \intermediateWiresStage6[1] [34], 
      \intermediateWiresStage6[1] [33], \intermediateWiresStage6[1] [32], 
      \intermediateWiresStage6[1] [31], \intermediateWiresStage6[1] [30], 
      \intermediateWiresStage6[1] [29], \intermediateWiresStage6[1] [28], 
      \intermediateWiresStage6[1] [27], \intermediateWiresStage6[1] [26], 
      \intermediateWiresStage6[1] [25], \intermediateWiresStage6[1] [24], 
      \intermediateWiresStage6[1] [23], \intermediateWiresStage6[1] [22], 
      \intermediateWiresStage6[1] [21], \intermediateWiresStage6[1] [20], 
      \intermediateWiresStage6[1] [19], \intermediateWiresStage6[1] [18], 
      \intermediateWiresStage6[1] [17], \intermediateWiresStage6[1] [16], 
      \intermediateWiresStage6[1] [15], \intermediateWiresStage6[1] [14], 
      \intermediateWiresStage6[1] [13], \intermediateWiresStage6[1] [12], 
      \intermediateWiresStage6[1] [11], \intermediateWiresStage6[1] [10], 
      \intermediateWiresStage6[1] [9], \intermediateWiresStage6[1] [8], 
      \intermediateWiresStage6[1] [7], uc_4353, uc_4354, uc_4355, uc_4356, 
      uc_4357, uc_4358, uc_4359}), .A({1'b0, uc_4360, uc_4361, uc_4362, uc_4363, 
      uc_4364, uc_4365, uc_4366, uc_4367, uc_4368, uc_4369, uc_4370, uc_4371, 
      uc_4372, uc_4373, uc_4374, uc_4375, normalizedWires[1518], 
      \intermediateWiresStage1[14] [45], \intermediateWiresStage1[14] [44], 
      \intermediateWiresStage2[8] [43], \intermediateWiresStage4[2] [42], 
      \intermediateWiresStage4[2] [41], \intermediateWiresStage4[2] [40], 
      \intermediateWiresStage4[2] [39], \intermediateWiresStage4[2] [38], 
      \intermediateWiresStage5[0] [37], \intermediateWiresStage5[0] [36], 
      \intermediateWiresStage5[0] [35], \intermediateWiresStage5[0] [34], 
      \intermediateWiresStage5[0] [33], \intermediateWiresStage5[0] [32], 
      \intermediateWiresStage5[0] [31], \intermediateWiresStage5[0] [30], 
      \intermediateWiresStage5[0] [29], \intermediateWiresStage5[0] [28], 
      \intermediateWiresStage5[0] [27], \intermediateWiresStage5[0] [26], 
      \intermediateWiresStage5[0] [25], \intermediateWiresStage5[0] [24], 
      \intermediateWiresStage5[0] [23], \intermediateWiresStage5[0] [22], 
      \intermediateWiresStage5[0] [21], \intermediateWiresStage5[0] [20], 
      \intermediateWiresStage5[0] [19], \intermediateWiresStage5[0] [18], 
      \intermediateWiresStage5[0] [17], \intermediateWiresStage5[0] [16], 
      \intermediateWiresStage5[0] [15], \intermediateWiresStage5[0] [14], 
      \intermediateWiresStage5[0] [13], \intermediateWiresStage5[0] [12], 
      \intermediateWiresStage5[0] [11], \intermediateWiresStage5[0] [10], 
      \intermediateWiresStage5[0] [9], \intermediateWiresStage5[0] [8], 
      \intermediateWiresStage5[0] [7], \intermediateWiresStage5[0] [6], uc_4376, 
      uc_4377, uc_4378, uc_4379, uc_4380, uc_4381}), .B({1'b0, uc_4382, uc_4383, 
      uc_4384, uc_4385, uc_4386, uc_4387, uc_4388, uc_4389, uc_4390, uc_4391, 
      uc_4392, uc_4393, uc_4394, uc_4395, uc_4396, uc_4397, uc_4398, uc_4399, 
      uc_4400, uc_4401, uc_4402, uc_4403, uc_4404, uc_4405, 
      \intermediateWiresStage5[1] [38], \intermediateWiresStage5[1] [37], 
      \intermediateWiresStage5[1] [36], \intermediateWiresStage5[1] [35], 
      \intermediateWiresStage5[1] [34], \intermediateWiresStage5[1] [33], 
      \intermediateWiresStage5[1] [32], \intermediateWiresStage5[1] [31], 
      \intermediateWiresStage5[1] [30], \intermediateWiresStage5[1] [29], 
      \intermediateWiresStage5[1] [28], \intermediateWiresStage5[1] [27], 
      \intermediateWiresStage5[1] [26], \intermediateWiresStage5[1] [25], 
      \intermediateWiresStage5[1] [24], \intermediateWiresStage5[1] [23], 
      \intermediateWiresStage5[1] [22], \intermediateWiresStage5[1] [21], 
      \intermediateWiresStage5[1] [20], \intermediateWiresStage5[1] [19], 
      \intermediateWiresStage5[1] [18], \intermediateWiresStage5[1] [17], 
      \intermediateWiresStage5[1] [16], \intermediateWiresStage5[1] [15], 
      \intermediateWiresStage5[1] [14], \intermediateWiresStage5[1] [13], 
      \intermediateWiresStage5[1] [12], \intermediateWiresStage5[1] [11], 
      \intermediateWiresStage5[1] [10], \intermediateWiresStage5[1] [9], 
      \intermediateWiresStage5[1] [8], \intermediateWiresStage5[1] [7], 
      \intermediateWiresStage5[1] [6], uc_4406, uc_4407, uc_4408, uc_4409, 
      uc_4410, uc_4411}), .C({1'b0, uc_4412, uc_4413, uc_4414, uc_4415, uc_4416, 
      uc_4417, uc_4418, uc_4419, uc_4420, uc_4421, uc_4422, uc_4423, uc_4424, 
      uc_4425, uc_4426, uc_4427, \intermediateWiresStage5[2] [46], 
      \intermediateWiresStage5[2] [45], \intermediateWiresStage5[2] [44], 
      \intermediateWiresStage5[2] [43], \intermediateWiresStage5[2] [42], 
      \intermediateWiresStage5[2] [41], \intermediateWiresStage5[2] [40], 
      \intermediateWiresStage5[2] [39], \intermediateWiresStage5[2] [38], 
      \intermediateWiresStage5[2] [37], \intermediateWiresStage5[2] [36], 
      \intermediateWiresStage5[2] [35], \intermediateWiresStage5[2] [34], 
      \intermediateWiresStage5[2] [33], \intermediateWiresStage5[2] [32], 
      \intermediateWiresStage5[2] [31], \intermediateWiresStage5[2] [30], 
      \intermediateWiresStage5[2] [29], \intermediateWiresStage5[2] [28], 
      \intermediateWiresStage5[2] [27], \intermediateWiresStage5[2] [26], 
      \intermediateWiresStage5[2] [25], \intermediateWiresStage5[2] [24], 
      \intermediateWiresStage5[2] [23], \intermediateWiresStage5[2] [22], 
      \intermediateWiresStage5[2] [21], \intermediateWiresStage4[3] [20], 
      \intermediateWiresStage4[3] [19], \intermediateWiresStage4[3] [18], 
      \intermediateWiresStage4[3] [17], \intermediateWiresStage4[3] [16], 
      \intermediateWiresStage4[3] [15], uc_4428, uc_4429, uc_4430, uc_4431, 
      uc_4432, uc_4433, uc_4434, uc_4435, uc_4436, uc_4437, uc_4438, uc_4439, 
      uc_4440, uc_4441, uc_4442}));
   CSAlike__4_2018 genblk8_0_parallelAdderStage7 (.result({uc_4443, uc_4444, 
      uc_4445, uc_4446, uc_4447, uc_4448, uc_4449, uc_4450, uc_4451, uc_4452, 
      uc_4453, uc_4454, uc_4455, uc_4456, uc_4457, uc_4458, 
      \intermediateWiresStage7[0] [47], \intermediateWiresStage7[0] [46], 
      \intermediateWiresStage7[0] [45], \intermediateWiresStage7[0] [44], 
      \intermediateWiresStage7[0] [43], \intermediateWiresStage7[0] [42], 
      \intermediateWiresStage7[0] [41], \intermediateWiresStage7[0] [40], 
      \intermediateWiresStage7[0] [39], \intermediateWiresStage7[0] [38], 
      \intermediateWiresStage7[0] [37], \intermediateWiresStage7[0] [36], 
      \intermediateWiresStage7[0] [35], \intermediateWiresStage7[0] [34], 
      \intermediateWiresStage7[0] [33], \intermediateWiresStage7[0] [32], 
      \intermediateWiresStage7[0] [31], \intermediateWiresStage7[0] [30], 
      \intermediateWiresStage7[0] [29], \intermediateWiresStage7[0] [28], 
      \intermediateWiresStage7[0] [27], \intermediateWiresStage7[0] [26], 
      \intermediateWiresStage7[0] [25], \intermediateWiresStage7[0] [24], 
      \intermediateWiresStage7[0] [23], \intermediateWiresStage7[0] [22], 
      \intermediateWiresStage7[0] [21], \intermediateWiresStage7[0] [20], 
      \intermediateWiresStage7[0] [19], \intermediateWiresStage7[0] [18], 
      \intermediateWiresStage7[0] [17], \intermediateWiresStage7[0] [16], 
      \intermediateWiresStage7[0] [15], \intermediateWiresStage7[0] [14], 
      \intermediateWiresStage7[0] [13], \intermediateWiresStage7[0] [12], 
      \intermediateWiresStage7[0] [11], \intermediateWiresStage7[0] [10], 
      \intermediateWiresStage7[0] [9], \intermediateWiresStage7[0] [8], uc_4459, 
      uc_4460, uc_4461, uc_4462, uc_4463, uc_4464, uc_4465, uc_4466}), .carry({
      uc_4467, uc_4468, uc_4469, uc_4470, uc_4471, uc_4472, uc_4473, uc_4474, 
      uc_4475, uc_4476, uc_4477, uc_4478, uc_4479, uc_4480, uc_4481, uc_4482, 
      \intermediateWiresStage7[1] [47], \intermediateWiresStage7[1] [46], 
      \intermediateWiresStage7[1] [45], \intermediateWiresStage7[1] [44], 
      \intermediateWiresStage7[1] [43], \intermediateWiresStage7[1] [42], 
      \intermediateWiresStage7[1] [41], \intermediateWiresStage7[1] [40], 
      \intermediateWiresStage7[1] [39], \intermediateWiresStage7[1] [38], 
      \intermediateWiresStage7[1] [37], \intermediateWiresStage7[1] [36], 
      \intermediateWiresStage7[1] [35], \intermediateWiresStage7[1] [34], 
      \intermediateWiresStage7[1] [33], \intermediateWiresStage7[1] [32], 
      \intermediateWiresStage7[1] [31], \intermediateWiresStage7[1] [30], 
      \intermediateWiresStage7[1] [29], \intermediateWiresStage7[1] [28], 
      \intermediateWiresStage7[1] [27], \intermediateWiresStage7[1] [26], 
      \intermediateWiresStage7[1] [25], \intermediateWiresStage7[1] [24], 
      \intermediateWiresStage7[1] [23], \intermediateWiresStage7[1] [22], 
      \intermediateWiresStage7[1] [21], \intermediateWiresStage7[1] [20], 
      \intermediateWiresStage7[1] [19], \intermediateWiresStage7[1] [18], 
      \intermediateWiresStage7[1] [17], \intermediateWiresStage7[1] [16], 
      \intermediateWiresStage7[1] [15], \intermediateWiresStage7[1] [14], 
      \intermediateWiresStage7[1] [13], \intermediateWiresStage7[1] [12], 
      \intermediateWiresStage7[1] [11], \intermediateWiresStage7[1] [10], 
      \intermediateWiresStage7[1] [9], \intermediateWiresStage7[1] [8], uc_4483, 
      uc_4484, uc_4485, uc_4486, uc_4487, uc_4488, uc_4489, uc_4490}), .A({1'b0, 
      uc_4491, uc_4492, uc_4493, uc_4494, uc_4495, uc_4496, uc_4497, uc_4498, 
      uc_4499, uc_4500, uc_4501, uc_4502, uc_4503, uc_4504, uc_4505, uc_4506, 
      \intermediateWiresStage6[0] [46], \intermediateWiresStage6[0] [45], 
      \intermediateWiresStage6[0] [44], \intermediateWiresStage6[0] [43], 
      \intermediateWiresStage6[0] [42], \intermediateWiresStage6[0] [41], 
      \intermediateWiresStage6[0] [40], \intermediateWiresStage6[0] [39], 
      \intermediateWiresStage6[0] [38], \intermediateWiresStage6[0] [37], 
      \intermediateWiresStage6[0] [36], \intermediateWiresStage6[0] [35], 
      \intermediateWiresStage6[0] [34], \intermediateWiresStage6[0] [33], 
      \intermediateWiresStage6[0] [32], \intermediateWiresStage6[0] [31], 
      \intermediateWiresStage6[0] [30], \intermediateWiresStage6[0] [29], 
      \intermediateWiresStage6[0] [28], \intermediateWiresStage6[0] [27], 
      \intermediateWiresStage6[0] [26], \intermediateWiresStage6[0] [25], 
      \intermediateWiresStage6[0] [24], \intermediateWiresStage6[0] [23], 
      \intermediateWiresStage6[0] [22], \intermediateWiresStage6[0] [21], 
      \intermediateWiresStage6[0] [20], \intermediateWiresStage6[0] [19], 
      \intermediateWiresStage6[0] [18], \intermediateWiresStage6[0] [17], 
      \intermediateWiresStage6[0] [16], \intermediateWiresStage6[0] [15], 
      \intermediateWiresStage6[0] [14], \intermediateWiresStage6[0] [13], 
      \intermediateWiresStage6[0] [12], \intermediateWiresStage6[0] [11], 
      \intermediateWiresStage6[0] [10], \intermediateWiresStage6[0] [9], 
      \intermediateWiresStage6[0] [8], \intermediateWiresStage6[0] [7], uc_4507, 
      uc_4508, uc_4509, uc_4510, uc_4511, uc_4512, uc_4513}), .B({1'b0, uc_4514, 
      uc_4515, uc_4516, uc_4517, uc_4518, uc_4519, uc_4520, uc_4521, uc_4522, 
      uc_4523, uc_4524, uc_4525, uc_4526, uc_4527, uc_4528, 
      \intermediateWiresStage6[1] [47], \intermediateWiresStage6[1] [46], 
      \intermediateWiresStage6[1] [45], \intermediateWiresStage6[1] [44], 
      \intermediateWiresStage6[1] [43], \intermediateWiresStage6[1] [42], 
      \intermediateWiresStage6[1] [41], \intermediateWiresStage6[1] [40], 
      \intermediateWiresStage6[1] [39], \intermediateWiresStage6[1] [38], 
      \intermediateWiresStage6[1] [37], \intermediateWiresStage6[1] [36], 
      \intermediateWiresStage6[1] [35], \intermediateWiresStage6[1] [34], 
      \intermediateWiresStage6[1] [33], \intermediateWiresStage6[1] [32], 
      \intermediateWiresStage6[1] [31], \intermediateWiresStage6[1] [30], 
      \intermediateWiresStage6[1] [29], \intermediateWiresStage6[1] [28], 
      \intermediateWiresStage6[1] [27], \intermediateWiresStage6[1] [26], 
      \intermediateWiresStage6[1] [25], \intermediateWiresStage6[1] [24], 
      \intermediateWiresStage6[1] [23], \intermediateWiresStage6[1] [22], 
      \intermediateWiresStage6[1] [21], \intermediateWiresStage6[1] [20], 
      \intermediateWiresStage6[1] [19], \intermediateWiresStage6[1] [18], 
      \intermediateWiresStage6[1] [17], \intermediateWiresStage6[1] [16], 
      \intermediateWiresStage6[1] [15], \intermediateWiresStage6[1] [14], 
      \intermediateWiresStage6[1] [13], \intermediateWiresStage6[1] [12], 
      \intermediateWiresStage6[1] [11], \intermediateWiresStage6[1] [10], 
      \intermediateWiresStage6[1] [9], \intermediateWiresStage6[1] [8], 
      \intermediateWiresStage6[1] [7], uc_4529, uc_4530, uc_4531, uc_4532, 
      uc_4533, uc_4534, uc_4535}), .C({1'b0, uc_4536, uc_4537, uc_4538, uc_4539, 
      uc_4540, uc_4541, uc_4542, uc_4543, uc_4544, uc_4545, uc_4546, uc_4547, 
      uc_4548, uc_4549, uc_4550, \intermediateWiresStage5[3] [47], 
      \intermediateWiresStage5[3] [46], \intermediateWiresStage5[3] [45], 
      \intermediateWiresStage5[3] [44], \intermediateWiresStage5[3] [43], 
      \intermediateWiresStage5[3] [42], \intermediateWiresStage5[3] [41], 
      \intermediateWiresStage5[3] [40], \intermediateWiresStage5[3] [39], 
      \intermediateWiresStage5[3] [38], \intermediateWiresStage5[3] [37], 
      \intermediateWiresStage5[3] [36], \intermediateWiresStage5[3] [35], 
      \intermediateWiresStage5[3] [34], \intermediateWiresStage5[3] [33], 
      \intermediateWiresStage5[3] [32], \intermediateWiresStage5[3] [31], 
      \intermediateWiresStage5[3] [30], \intermediateWiresStage5[3] [29], 
      \intermediateWiresStage5[3] [28], \intermediateWiresStage5[3] [27], 
      \intermediateWiresStage5[3] [26], \intermediateWiresStage5[3] [25], 
      \intermediateWiresStage5[3] [24], \intermediateWiresStage5[3] [23], 
      \intermediateWiresStage5[3] [22], uc_4551, uc_4552, uc_4553, uc_4554, 
      uc_4555, uc_4556, uc_4557, uc_4558, uc_4559, uc_4560, uc_4561, uc_4562, 
      uc_4563, uc_4564, uc_4565, uc_4566, uc_4567, uc_4568, uc_4569, uc_4570, 
      uc_4571, uc_4572}));
   CSAlike genblk9_0_finalStage (.result({uc_4573, uc_4574, uc_4575, uc_4576, 
      uc_4577, uc_4578, uc_4579, uc_4580, uc_4581, uc_4582, uc_4583, uc_4584, 
      uc_4585, uc_4586, uc_4587, uc_4588, Res[47], Res[46], Res[45], Res[44], 
      Res[43], Res[42], Res[41], Res[40], Res[39], Res[38], Res[37], Res[36], 
      Res[35], Res[34], Res[33], Res[32], Res[31], Res[30], Res[29], Res[28], 
      Res[27], Res[26], Res[25], Res[24], Res[23], Res[22], Res[21], Res[20], 
      Res[19], Res[18], Res[17], Res[16], Res[15], Res[14], Res[13], Res[12], 
      Res[11], Res[10], Res[9], uc_4589, uc_4590, uc_4591, uc_4592, uc_4593, 
      uc_4594, uc_4595, uc_4596, uc_4597}), .carry({uc_4598, uc_4599, uc_4600, 
      uc_4601, uc_4602, uc_4603, uc_4604, uc_4605, uc_4606, uc_4607, uc_4608, 
      uc_4609, uc_4610, uc_4611, uc_4612, uc_4613, carry[47], carry[46], 
      carry[45], carry[44], carry[43], carry[42], carry[41], carry[40], 
      carry[39], carry[38], carry[37], carry[36], carry[35], carry[34], 
      carry[33], carry[32], carry[31], carry[30], carry[29], carry[28], 
      carry[27], carry[26], carry[25], carry[24], carry[23], carry[22], 
      carry[21], carry[20], carry[19], carry[18], carry[17], carry[16], 
      carry[15], carry[14], carry[13], carry[12], carry[11], carry[10], carry[9], 
      uc_4614, uc_4615, uc_4616, uc_4617, uc_4618, uc_4619, uc_4620, uc_4621, 
      uc_4622}), .A({1'b0, uc_4623, uc_4624, uc_4625, uc_4626, uc_4627, uc_4628, 
      uc_4629, uc_4630, uc_4631, uc_4632, uc_4633, uc_4634, uc_4635, uc_4636, 
      uc_4637, \intermediateWiresStage7[0] [47], 
      \intermediateWiresStage7[0] [46], \intermediateWiresStage7[0] [45], 
      \intermediateWiresStage7[0] [44], \intermediateWiresStage7[0] [43], 
      \intermediateWiresStage7[0] [42], \intermediateWiresStage7[0] [41], 
      \intermediateWiresStage7[0] [40], \intermediateWiresStage7[0] [39], 
      \intermediateWiresStage7[0] [38], \intermediateWiresStage7[0] [37], 
      \intermediateWiresStage7[0] [36], \intermediateWiresStage7[0] [35], 
      \intermediateWiresStage7[0] [34], \intermediateWiresStage7[0] [33], 
      \intermediateWiresStage7[0] [32], \intermediateWiresStage7[0] [31], 
      \intermediateWiresStage7[0] [30], \intermediateWiresStage7[0] [29], 
      \intermediateWiresStage7[0] [28], \intermediateWiresStage7[0] [27], 
      \intermediateWiresStage7[0] [26], \intermediateWiresStage7[0] [25], 
      \intermediateWiresStage7[0] [24], \intermediateWiresStage7[0] [23], 
      \intermediateWiresStage7[0] [22], \intermediateWiresStage7[0] [21], 
      \intermediateWiresStage7[0] [20], \intermediateWiresStage7[0] [19], 
      \intermediateWiresStage7[0] [18], \intermediateWiresStage7[0] [17], 
      \intermediateWiresStage7[0] [16], \intermediateWiresStage7[0] [15], 
      \intermediateWiresStage7[0] [14], \intermediateWiresStage7[0] [13], 
      \intermediateWiresStage7[0] [12], \intermediateWiresStage7[0] [11], 
      \intermediateWiresStage7[0] [10], \intermediateWiresStage7[0] [9], 
      \intermediateWiresStage7[0] [8], uc_4638, uc_4639, uc_4640, uc_4641, 
      uc_4642, uc_4643, uc_4644, uc_4645}), .B({1'b0, uc_4646, uc_4647, uc_4648, 
      uc_4649, uc_4650, uc_4651, uc_4652, uc_4653, uc_4654, uc_4655, uc_4656, 
      uc_4657, uc_4658, uc_4659, uc_4660, \intermediateWiresStage7[1] [47], 
      \intermediateWiresStage7[1] [46], \intermediateWiresStage7[1] [45], 
      \intermediateWiresStage7[1] [44], \intermediateWiresStage7[1] [43], 
      \intermediateWiresStage7[1] [42], \intermediateWiresStage7[1] [41], 
      \intermediateWiresStage7[1] [40], \intermediateWiresStage7[1] [39], 
      \intermediateWiresStage7[1] [38], \intermediateWiresStage7[1] [37], 
      \intermediateWiresStage7[1] [36], \intermediateWiresStage7[1] [35], 
      \intermediateWiresStage7[1] [34], \intermediateWiresStage7[1] [33], 
      \intermediateWiresStage7[1] [32], \intermediateWiresStage7[1] [31], 
      \intermediateWiresStage7[1] [30], \intermediateWiresStage7[1] [29], 
      \intermediateWiresStage7[1] [28], \intermediateWiresStage7[1] [27], 
      \intermediateWiresStage7[1] [26], \intermediateWiresStage7[1] [25], 
      \intermediateWiresStage7[1] [24], \intermediateWiresStage7[1] [23], 
      \intermediateWiresStage7[1] [22], \intermediateWiresStage7[1] [21], 
      \intermediateWiresStage7[1] [20], \intermediateWiresStage7[1] [19], 
      \intermediateWiresStage7[1] [18], \intermediateWiresStage7[1] [17], 
      \intermediateWiresStage7[1] [16], \intermediateWiresStage7[1] [15], 
      \intermediateWiresStage7[1] [14], \intermediateWiresStage7[1] [13], 
      \intermediateWiresStage7[1] [12], \intermediateWiresStage7[1] [11], 
      \intermediateWiresStage7[1] [10], \intermediateWiresStage7[1] [9], 
      \intermediateWiresStage7[1] [8], uc_4661, uc_4662, uc_4663, uc_4664, 
      uc_4665, uc_4666, uc_4667, uc_4668}), .C({1'b0, uc_4669, uc_4670, uc_4671, 
      uc_4672, uc_4673, uc_4674, uc_4675, uc_4676, uc_4677, uc_4678, uc_4679, 
      uc_4680, uc_4681, uc_4682, uc_4683, uc_4684, uc_4685, uc_4686, uc_4687, 
      uc_4688, uc_4689, uc_4690, uc_4691, uc_4692, uc_4693, uc_4694, uc_4695, 
      uc_4696, uc_4697, uc_4698, uc_4699, uc_4700, uc_4701, uc_4702, uc_4703, 
      uc_4704, uc_4705, uc_4706, uc_4707, uc_4708, uc_4709, uc_4710, uc_4711, 
      uc_4712, uc_4713, uc_4714, uc_4715, uc_4716, uc_4717, uc_4718, uc_4719, 
      uc_4720, uc_4721, uc_4722, uc_4723, uc_4724, uc_4725, uc_4726, uc_4727, 
      uc_4728, uc_4729, uc_4730, uc_4731}));
endmodule

module multiplyAllBits(normalizedWires, A, B);
   output [2047:0]normalizedWires;
   input [31:0]A;
   input [31:0]B;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;

   INV_X1 i_0_0 (.A(B[0]), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(A[0]), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(A[1]), .ZN(n_0_2));
   NOR2_X1 i_0_3 (.A1(n_0_0), .A2(n_0_2), .ZN(normalizedWires[1]));
   INV_X1 i_0_5 (.A(A[2]), .ZN(n_0_3));
   NOR2_X1 i_0_6 (.A1(n_0_0), .A2(n_0_3), .ZN(normalizedWires[2]));
   INV_X1 i_0_7 (.A(A[3]), .ZN(n_0_4));
   NOR2_X1 i_0_8 (.A1(n_0_0), .A2(n_0_4), .ZN(normalizedWires[3]));
   INV_X1 i_0_9 (.A(A[4]), .ZN(n_0_5));
   NOR2_X1 i_0_10 (.A1(n_0_0), .A2(n_0_5), .ZN(normalizedWires[4]));
   INV_X1 i_0_11 (.A(A[5]), .ZN(n_0_6));
   NOR2_X1 i_0_12 (.A1(n_0_0), .A2(n_0_6), .ZN(normalizedWires[5]));
   INV_X1 i_0_13 (.A(A[6]), .ZN(n_0_7));
   NOR2_X1 i_0_14 (.A1(n_0_0), .A2(n_0_7), .ZN(normalizedWires[6]));
   INV_X1 i_0_15 (.A(A[7]), .ZN(n_0_8));
   NOR2_X1 i_0_16 (.A1(n_0_0), .A2(n_0_8), .ZN(normalizedWires[7]));
   INV_X1 i_0_17 (.A(A[8]), .ZN(n_0_9));
   NOR2_X1 i_0_18 (.A1(n_0_0), .A2(n_0_9), .ZN(normalizedWires[8]));
   INV_X1 i_0_19 (.A(A[9]), .ZN(n_0_10));
   NOR2_X1 i_0_20 (.A1(n_0_0), .A2(n_0_10), .ZN(normalizedWires[9]));
   INV_X1 i_0_21 (.A(A[10]), .ZN(n_0_11));
   NOR2_X1 i_0_22 (.A1(n_0_0), .A2(n_0_11), .ZN(normalizedWires[10]));
   INV_X1 i_0_23 (.A(A[11]), .ZN(n_0_12));
   NOR2_X1 i_0_24 (.A1(n_0_0), .A2(n_0_12), .ZN(normalizedWires[11]));
   INV_X1 i_0_25 (.A(A[12]), .ZN(n_0_13));
   NOR2_X1 i_0_26 (.A1(n_0_0), .A2(n_0_13), .ZN(normalizedWires[12]));
   INV_X1 i_0_27 (.A(A[13]), .ZN(n_0_14));
   NOR2_X1 i_0_28 (.A1(n_0_0), .A2(n_0_14), .ZN(normalizedWires[13]));
   INV_X1 i_0_29 (.A(A[14]), .ZN(n_0_15));
   NOR2_X1 i_0_30 (.A1(n_0_0), .A2(n_0_15), .ZN(normalizedWires[14]));
   INV_X1 i_0_31 (.A(A[15]), .ZN(n_0_16));
   NOR2_X1 i_0_32 (.A1(n_0_0), .A2(n_0_16), .ZN(normalizedWires[15]));
   INV_X1 i_0_33 (.A(A[16]), .ZN(n_0_17));
   NOR2_X1 i_0_34 (.A1(n_0_0), .A2(n_0_17), .ZN(normalizedWires[16]));
   INV_X1 i_0_35 (.A(A[17]), .ZN(n_0_18));
   NOR2_X1 i_0_36 (.A1(n_0_0), .A2(n_0_18), .ZN(normalizedWires[17]));
   INV_X1 i_0_37 (.A(A[18]), .ZN(n_0_19));
   NOR2_X1 i_0_38 (.A1(n_0_0), .A2(n_0_19), .ZN(normalizedWires[18]));
   INV_X1 i_0_39 (.A(A[19]), .ZN(n_0_20));
   NOR2_X1 i_0_40 (.A1(n_0_0), .A2(n_0_20), .ZN(normalizedWires[19]));
   INV_X1 i_0_41 (.A(A[20]), .ZN(n_0_21));
   NOR2_X1 i_0_42 (.A1(n_0_0), .A2(n_0_21), .ZN(normalizedWires[20]));
   INV_X1 i_0_43 (.A(A[21]), .ZN(n_0_22));
   NOR2_X1 i_0_44 (.A1(n_0_0), .A2(n_0_22), .ZN(normalizedWires[21]));
   INV_X1 i_0_45 (.A(A[22]), .ZN(n_0_23));
   NOR2_X1 i_0_46 (.A1(n_0_0), .A2(n_0_23), .ZN(normalizedWires[22]));
   INV_X1 i_0_47 (.A(A[23]), .ZN(n_0_24));
   NOR2_X1 i_0_48 (.A1(n_0_0), .A2(n_0_24), .ZN(normalizedWires[23]));
   INV_X1 i_0_49 (.A(B[1]), .ZN(n_0_25));
   NOR2_X1 i_0_50 (.A1(n_0_25), .A2(n_0_1), .ZN(normalizedWires[65]));
   NOR2_X1 i_0_51 (.A1(n_0_25), .A2(n_0_2), .ZN(normalizedWires[66]));
   NOR2_X1 i_0_52 (.A1(n_0_25), .A2(n_0_3), .ZN(normalizedWires[67]));
   NOR2_X1 i_0_53 (.A1(n_0_25), .A2(n_0_4), .ZN(normalizedWires[68]));
   NOR2_X1 i_0_54 (.A1(n_0_25), .A2(n_0_5), .ZN(normalizedWires[69]));
   NOR2_X1 i_0_55 (.A1(n_0_25), .A2(n_0_6), .ZN(normalizedWires[70]));
   NOR2_X1 i_0_56 (.A1(n_0_25), .A2(n_0_7), .ZN(normalizedWires[71]));
   NOR2_X1 i_0_57 (.A1(n_0_25), .A2(n_0_8), .ZN(normalizedWires[72]));
   NOR2_X1 i_0_58 (.A1(n_0_25), .A2(n_0_9), .ZN(normalizedWires[73]));
   NOR2_X1 i_0_59 (.A1(n_0_25), .A2(n_0_10), .ZN(normalizedWires[74]));
   NOR2_X1 i_0_60 (.A1(n_0_25), .A2(n_0_11), .ZN(normalizedWires[75]));
   NOR2_X1 i_0_61 (.A1(n_0_25), .A2(n_0_12), .ZN(normalizedWires[76]));
   NOR2_X1 i_0_62 (.A1(n_0_25), .A2(n_0_13), .ZN(normalizedWires[77]));
   NOR2_X1 i_0_63 (.A1(n_0_25), .A2(n_0_14), .ZN(normalizedWires[78]));
   NOR2_X1 i_0_64 (.A1(n_0_25), .A2(n_0_15), .ZN(normalizedWires[79]));
   NOR2_X1 i_0_65 (.A1(n_0_25), .A2(n_0_16), .ZN(normalizedWires[80]));
   NOR2_X1 i_0_66 (.A1(n_0_25), .A2(n_0_17), .ZN(normalizedWires[81]));
   NOR2_X1 i_0_67 (.A1(n_0_25), .A2(n_0_18), .ZN(normalizedWires[82]));
   NOR2_X1 i_0_68 (.A1(n_0_25), .A2(n_0_19), .ZN(normalizedWires[83]));
   NOR2_X1 i_0_69 (.A1(n_0_25), .A2(n_0_20), .ZN(normalizedWires[84]));
   NOR2_X1 i_0_70 (.A1(n_0_25), .A2(n_0_21), .ZN(normalizedWires[85]));
   NOR2_X1 i_0_71 (.A1(n_0_25), .A2(n_0_22), .ZN(normalizedWires[86]));
   NOR2_X1 i_0_72 (.A1(n_0_25), .A2(n_0_23), .ZN(normalizedWires[87]));
   NOR2_X1 i_0_73 (.A1(n_0_25), .A2(n_0_24), .ZN(normalizedWires[88]));
   INV_X1 i_0_74 (.A(B[2]), .ZN(n_0_26));
   NOR2_X1 i_0_75 (.A1(n_0_26), .A2(n_0_1), .ZN(normalizedWires[130]));
   NOR2_X1 i_0_76 (.A1(n_0_26), .A2(n_0_2), .ZN(normalizedWires[131]));
   NOR2_X1 i_0_77 (.A1(n_0_26), .A2(n_0_3), .ZN(normalizedWires[132]));
   NOR2_X1 i_0_78 (.A1(n_0_26), .A2(n_0_4), .ZN(normalizedWires[133]));
   NOR2_X1 i_0_79 (.A1(n_0_26), .A2(n_0_5), .ZN(normalizedWires[134]));
   NOR2_X1 i_0_80 (.A1(n_0_26), .A2(n_0_6), .ZN(normalizedWires[135]));
   NOR2_X1 i_0_81 (.A1(n_0_26), .A2(n_0_7), .ZN(normalizedWires[136]));
   NOR2_X1 i_0_82 (.A1(n_0_26), .A2(n_0_8), .ZN(normalizedWires[137]));
   NOR2_X1 i_0_83 (.A1(n_0_26), .A2(n_0_9), .ZN(normalizedWires[138]));
   NOR2_X1 i_0_84 (.A1(n_0_26), .A2(n_0_10), .ZN(normalizedWires[139]));
   NOR2_X1 i_0_85 (.A1(n_0_26), .A2(n_0_11), .ZN(normalizedWires[140]));
   NOR2_X1 i_0_86 (.A1(n_0_26), .A2(n_0_12), .ZN(normalizedWires[141]));
   NOR2_X1 i_0_87 (.A1(n_0_26), .A2(n_0_13), .ZN(normalizedWires[142]));
   NOR2_X1 i_0_88 (.A1(n_0_26), .A2(n_0_14), .ZN(normalizedWires[143]));
   NOR2_X1 i_0_89 (.A1(n_0_26), .A2(n_0_15), .ZN(normalizedWires[144]));
   NOR2_X1 i_0_90 (.A1(n_0_26), .A2(n_0_16), .ZN(normalizedWires[145]));
   NOR2_X1 i_0_91 (.A1(n_0_26), .A2(n_0_17), .ZN(normalizedWires[146]));
   NOR2_X1 i_0_92 (.A1(n_0_26), .A2(n_0_18), .ZN(normalizedWires[147]));
   NOR2_X1 i_0_93 (.A1(n_0_26), .A2(n_0_19), .ZN(normalizedWires[148]));
   NOR2_X1 i_0_94 (.A1(n_0_26), .A2(n_0_20), .ZN(normalizedWires[149]));
   NOR2_X1 i_0_95 (.A1(n_0_26), .A2(n_0_21), .ZN(normalizedWires[150]));
   NOR2_X1 i_0_96 (.A1(n_0_26), .A2(n_0_22), .ZN(normalizedWires[151]));
   NOR2_X1 i_0_97 (.A1(n_0_26), .A2(n_0_23), .ZN(normalizedWires[152]));
   NOR2_X1 i_0_98 (.A1(n_0_26), .A2(n_0_24), .ZN(normalizedWires[153]));
   INV_X1 i_0_99 (.A(B[3]), .ZN(n_0_27));
   NOR2_X1 i_0_100 (.A1(n_0_27), .A2(n_0_1), .ZN(normalizedWires[195]));
   NOR2_X1 i_0_101 (.A1(n_0_27), .A2(n_0_2), .ZN(normalizedWires[196]));
   NOR2_X1 i_0_102 (.A1(n_0_27), .A2(n_0_3), .ZN(normalizedWires[197]));
   NOR2_X1 i_0_103 (.A1(n_0_27), .A2(n_0_4), .ZN(normalizedWires[198]));
   NOR2_X1 i_0_104 (.A1(n_0_27), .A2(n_0_5), .ZN(normalizedWires[199]));
   NOR2_X1 i_0_105 (.A1(n_0_27), .A2(n_0_6), .ZN(normalizedWires[200]));
   NOR2_X1 i_0_106 (.A1(n_0_27), .A2(n_0_7), .ZN(normalizedWires[201]));
   NOR2_X1 i_0_107 (.A1(n_0_27), .A2(n_0_8), .ZN(normalizedWires[202]));
   NOR2_X1 i_0_108 (.A1(n_0_27), .A2(n_0_9), .ZN(normalizedWires[203]));
   NOR2_X1 i_0_109 (.A1(n_0_27), .A2(n_0_10), .ZN(normalizedWires[204]));
   NOR2_X1 i_0_110 (.A1(n_0_27), .A2(n_0_11), .ZN(normalizedWires[205]));
   NOR2_X1 i_0_111 (.A1(n_0_27), .A2(n_0_12), .ZN(normalizedWires[206]));
   NOR2_X1 i_0_112 (.A1(n_0_27), .A2(n_0_13), .ZN(normalizedWires[207]));
   NOR2_X1 i_0_113 (.A1(n_0_27), .A2(n_0_14), .ZN(normalizedWires[208]));
   NOR2_X1 i_0_114 (.A1(n_0_27), .A2(n_0_15), .ZN(normalizedWires[209]));
   NOR2_X1 i_0_115 (.A1(n_0_27), .A2(n_0_16), .ZN(normalizedWires[210]));
   NOR2_X1 i_0_116 (.A1(n_0_27), .A2(n_0_17), .ZN(normalizedWires[211]));
   NOR2_X1 i_0_117 (.A1(n_0_27), .A2(n_0_18), .ZN(normalizedWires[212]));
   NOR2_X1 i_0_118 (.A1(n_0_27), .A2(n_0_19), .ZN(normalizedWires[213]));
   NOR2_X1 i_0_119 (.A1(n_0_27), .A2(n_0_20), .ZN(normalizedWires[214]));
   NOR2_X1 i_0_120 (.A1(n_0_27), .A2(n_0_21), .ZN(normalizedWires[215]));
   NOR2_X1 i_0_121 (.A1(n_0_27), .A2(n_0_22), .ZN(normalizedWires[216]));
   NOR2_X1 i_0_122 (.A1(n_0_27), .A2(n_0_23), .ZN(normalizedWires[217]));
   NOR2_X1 i_0_123 (.A1(n_0_27), .A2(n_0_24), .ZN(normalizedWires[218]));
   INV_X1 i_0_124 (.A(B[4]), .ZN(n_0_28));
   NOR2_X1 i_0_125 (.A1(n_0_28), .A2(n_0_1), .ZN(normalizedWires[260]));
   NOR2_X1 i_0_126 (.A1(n_0_28), .A2(n_0_2), .ZN(normalizedWires[261]));
   NOR2_X1 i_0_127 (.A1(n_0_28), .A2(n_0_3), .ZN(normalizedWires[262]));
   NOR2_X1 i_0_128 (.A1(n_0_28), .A2(n_0_4), .ZN(normalizedWires[263]));
   NOR2_X1 i_0_129 (.A1(n_0_28), .A2(n_0_5), .ZN(normalizedWires[264]));
   NOR2_X1 i_0_130 (.A1(n_0_28), .A2(n_0_6), .ZN(normalizedWires[265]));
   NOR2_X1 i_0_131 (.A1(n_0_28), .A2(n_0_7), .ZN(normalizedWires[266]));
   NOR2_X1 i_0_132 (.A1(n_0_28), .A2(n_0_8), .ZN(normalizedWires[267]));
   NOR2_X1 i_0_133 (.A1(n_0_28), .A2(n_0_9), .ZN(normalizedWires[268]));
   NOR2_X1 i_0_134 (.A1(n_0_28), .A2(n_0_10), .ZN(normalizedWires[269]));
   NOR2_X1 i_0_135 (.A1(n_0_28), .A2(n_0_11), .ZN(normalizedWires[270]));
   NOR2_X1 i_0_136 (.A1(n_0_28), .A2(n_0_12), .ZN(normalizedWires[271]));
   NOR2_X1 i_0_137 (.A1(n_0_28), .A2(n_0_13), .ZN(normalizedWires[272]));
   NOR2_X1 i_0_138 (.A1(n_0_28), .A2(n_0_14), .ZN(normalizedWires[273]));
   NOR2_X1 i_0_139 (.A1(n_0_28), .A2(n_0_15), .ZN(normalizedWires[274]));
   NOR2_X1 i_0_140 (.A1(n_0_28), .A2(n_0_16), .ZN(normalizedWires[275]));
   NOR2_X1 i_0_141 (.A1(n_0_28), .A2(n_0_17), .ZN(normalizedWires[276]));
   NOR2_X1 i_0_142 (.A1(n_0_28), .A2(n_0_18), .ZN(normalizedWires[277]));
   NOR2_X1 i_0_143 (.A1(n_0_28), .A2(n_0_19), .ZN(normalizedWires[278]));
   NOR2_X1 i_0_144 (.A1(n_0_28), .A2(n_0_20), .ZN(normalizedWires[279]));
   NOR2_X1 i_0_145 (.A1(n_0_28), .A2(n_0_21), .ZN(normalizedWires[280]));
   NOR2_X1 i_0_146 (.A1(n_0_28), .A2(n_0_22), .ZN(normalizedWires[281]));
   NOR2_X1 i_0_147 (.A1(n_0_28), .A2(n_0_23), .ZN(normalizedWires[282]));
   NOR2_X1 i_0_148 (.A1(n_0_28), .A2(n_0_24), .ZN(normalizedWires[283]));
   INV_X1 i_0_149 (.A(B[5]), .ZN(n_0_29));
   NOR2_X1 i_0_150 (.A1(n_0_29), .A2(n_0_1), .ZN(normalizedWires[325]));
   NOR2_X1 i_0_151 (.A1(n_0_29), .A2(n_0_2), .ZN(normalizedWires[326]));
   NOR2_X1 i_0_152 (.A1(n_0_29), .A2(n_0_3), .ZN(normalizedWires[327]));
   NOR2_X1 i_0_153 (.A1(n_0_29), .A2(n_0_4), .ZN(normalizedWires[328]));
   NOR2_X1 i_0_154 (.A1(n_0_29), .A2(n_0_5), .ZN(normalizedWires[329]));
   NOR2_X1 i_0_155 (.A1(n_0_29), .A2(n_0_6), .ZN(normalizedWires[330]));
   NOR2_X1 i_0_156 (.A1(n_0_29), .A2(n_0_7), .ZN(normalizedWires[331]));
   NOR2_X1 i_0_157 (.A1(n_0_29), .A2(n_0_8), .ZN(normalizedWires[332]));
   NOR2_X1 i_0_158 (.A1(n_0_29), .A2(n_0_9), .ZN(normalizedWires[333]));
   NOR2_X1 i_0_159 (.A1(n_0_29), .A2(n_0_10), .ZN(normalizedWires[334]));
   NOR2_X1 i_0_160 (.A1(n_0_29), .A2(n_0_11), .ZN(normalizedWires[335]));
   NOR2_X1 i_0_161 (.A1(n_0_29), .A2(n_0_12), .ZN(normalizedWires[336]));
   NOR2_X1 i_0_162 (.A1(n_0_29), .A2(n_0_13), .ZN(normalizedWires[337]));
   NOR2_X1 i_0_163 (.A1(n_0_29), .A2(n_0_14), .ZN(normalizedWires[338]));
   NOR2_X1 i_0_164 (.A1(n_0_29), .A2(n_0_15), .ZN(normalizedWires[339]));
   NOR2_X1 i_0_165 (.A1(n_0_29), .A2(n_0_16), .ZN(normalizedWires[340]));
   NOR2_X1 i_0_166 (.A1(n_0_29), .A2(n_0_17), .ZN(normalizedWires[341]));
   NOR2_X1 i_0_167 (.A1(n_0_29), .A2(n_0_18), .ZN(normalizedWires[342]));
   NOR2_X1 i_0_168 (.A1(n_0_29), .A2(n_0_19), .ZN(normalizedWires[343]));
   NOR2_X1 i_0_169 (.A1(n_0_29), .A2(n_0_20), .ZN(normalizedWires[344]));
   NOR2_X1 i_0_170 (.A1(n_0_29), .A2(n_0_21), .ZN(normalizedWires[345]));
   NOR2_X1 i_0_171 (.A1(n_0_29), .A2(n_0_22), .ZN(normalizedWires[346]));
   NOR2_X1 i_0_172 (.A1(n_0_29), .A2(n_0_23), .ZN(normalizedWires[347]));
   NOR2_X1 i_0_173 (.A1(n_0_29), .A2(n_0_24), .ZN(normalizedWires[348]));
   INV_X1 i_0_174 (.A(B[6]), .ZN(n_0_30));
   NOR2_X1 i_0_175 (.A1(n_0_30), .A2(n_0_1), .ZN(normalizedWires[390]));
   NOR2_X1 i_0_176 (.A1(n_0_30), .A2(n_0_2), .ZN(normalizedWires[391]));
   NOR2_X1 i_0_177 (.A1(n_0_30), .A2(n_0_3), .ZN(normalizedWires[392]));
   NOR2_X1 i_0_178 (.A1(n_0_30), .A2(n_0_4), .ZN(normalizedWires[393]));
   NOR2_X1 i_0_179 (.A1(n_0_30), .A2(n_0_5), .ZN(normalizedWires[394]));
   NOR2_X1 i_0_180 (.A1(n_0_30), .A2(n_0_6), .ZN(normalizedWires[395]));
   NOR2_X1 i_0_181 (.A1(n_0_30), .A2(n_0_7), .ZN(normalizedWires[396]));
   NOR2_X1 i_0_182 (.A1(n_0_30), .A2(n_0_8), .ZN(normalizedWires[397]));
   NOR2_X1 i_0_183 (.A1(n_0_30), .A2(n_0_9), .ZN(normalizedWires[398]));
   NOR2_X1 i_0_184 (.A1(n_0_30), .A2(n_0_10), .ZN(normalizedWires[399]));
   NOR2_X1 i_0_185 (.A1(n_0_30), .A2(n_0_11), .ZN(normalizedWires[400]));
   NOR2_X1 i_0_186 (.A1(n_0_30), .A2(n_0_12), .ZN(normalizedWires[401]));
   NOR2_X1 i_0_187 (.A1(n_0_30), .A2(n_0_13), .ZN(normalizedWires[402]));
   NOR2_X1 i_0_188 (.A1(n_0_30), .A2(n_0_14), .ZN(normalizedWires[403]));
   NOR2_X1 i_0_189 (.A1(n_0_30), .A2(n_0_15), .ZN(normalizedWires[404]));
   NOR2_X1 i_0_190 (.A1(n_0_30), .A2(n_0_16), .ZN(normalizedWires[405]));
   NOR2_X1 i_0_191 (.A1(n_0_30), .A2(n_0_17), .ZN(normalizedWires[406]));
   NOR2_X1 i_0_192 (.A1(n_0_30), .A2(n_0_18), .ZN(normalizedWires[407]));
   NOR2_X1 i_0_193 (.A1(n_0_30), .A2(n_0_19), .ZN(normalizedWires[408]));
   NOR2_X1 i_0_194 (.A1(n_0_30), .A2(n_0_20), .ZN(normalizedWires[409]));
   NOR2_X1 i_0_195 (.A1(n_0_30), .A2(n_0_21), .ZN(normalizedWires[410]));
   NOR2_X1 i_0_196 (.A1(n_0_30), .A2(n_0_22), .ZN(normalizedWires[411]));
   NOR2_X1 i_0_197 (.A1(n_0_30), .A2(n_0_23), .ZN(normalizedWires[412]));
   NOR2_X1 i_0_198 (.A1(n_0_30), .A2(n_0_24), .ZN(normalizedWires[413]));
   INV_X1 i_0_199 (.A(B[7]), .ZN(n_0_31));
   NOR2_X1 i_0_200 (.A1(n_0_31), .A2(n_0_1), .ZN(normalizedWires[455]));
   NOR2_X1 i_0_201 (.A1(n_0_31), .A2(n_0_2), .ZN(normalizedWires[456]));
   NOR2_X1 i_0_202 (.A1(n_0_31), .A2(n_0_3), .ZN(normalizedWires[457]));
   NOR2_X1 i_0_203 (.A1(n_0_31), .A2(n_0_4), .ZN(normalizedWires[458]));
   NOR2_X1 i_0_204 (.A1(n_0_31), .A2(n_0_5), .ZN(normalizedWires[459]));
   NOR2_X1 i_0_205 (.A1(n_0_31), .A2(n_0_6), .ZN(normalizedWires[460]));
   NOR2_X1 i_0_206 (.A1(n_0_31), .A2(n_0_7), .ZN(normalizedWires[461]));
   NOR2_X1 i_0_207 (.A1(n_0_31), .A2(n_0_8), .ZN(normalizedWires[462]));
   NOR2_X1 i_0_208 (.A1(n_0_31), .A2(n_0_9), .ZN(normalizedWires[463]));
   NOR2_X1 i_0_209 (.A1(n_0_31), .A2(n_0_10), .ZN(normalizedWires[464]));
   NOR2_X1 i_0_210 (.A1(n_0_31), .A2(n_0_11), .ZN(normalizedWires[465]));
   NOR2_X1 i_0_211 (.A1(n_0_31), .A2(n_0_12), .ZN(normalizedWires[466]));
   NOR2_X1 i_0_212 (.A1(n_0_31), .A2(n_0_13), .ZN(normalizedWires[467]));
   NOR2_X1 i_0_213 (.A1(n_0_31), .A2(n_0_14), .ZN(normalizedWires[468]));
   NOR2_X1 i_0_214 (.A1(n_0_31), .A2(n_0_15), .ZN(normalizedWires[469]));
   NOR2_X1 i_0_215 (.A1(n_0_31), .A2(n_0_16), .ZN(normalizedWires[470]));
   NOR2_X1 i_0_216 (.A1(n_0_31), .A2(n_0_17), .ZN(normalizedWires[471]));
   NOR2_X1 i_0_217 (.A1(n_0_31), .A2(n_0_18), .ZN(normalizedWires[472]));
   NOR2_X1 i_0_218 (.A1(n_0_31), .A2(n_0_19), .ZN(normalizedWires[473]));
   NOR2_X1 i_0_219 (.A1(n_0_31), .A2(n_0_20), .ZN(normalizedWires[474]));
   NOR2_X1 i_0_220 (.A1(n_0_31), .A2(n_0_21), .ZN(normalizedWires[475]));
   NOR2_X1 i_0_221 (.A1(n_0_31), .A2(n_0_22), .ZN(normalizedWires[476]));
   NOR2_X1 i_0_222 (.A1(n_0_31), .A2(n_0_23), .ZN(normalizedWires[477]));
   NOR2_X1 i_0_223 (.A1(n_0_31), .A2(n_0_24), .ZN(normalizedWires[478]));
   INV_X1 i_0_224 (.A(B[8]), .ZN(n_0_32));
   NOR2_X1 i_0_225 (.A1(n_0_32), .A2(n_0_1), .ZN(normalizedWires[520]));
   NOR2_X1 i_0_226 (.A1(n_0_32), .A2(n_0_2), .ZN(normalizedWires[521]));
   NOR2_X1 i_0_227 (.A1(n_0_32), .A2(n_0_3), .ZN(normalizedWires[522]));
   NOR2_X1 i_0_228 (.A1(n_0_32), .A2(n_0_4), .ZN(normalizedWires[523]));
   NOR2_X1 i_0_229 (.A1(n_0_32), .A2(n_0_5), .ZN(normalizedWires[524]));
   NOR2_X1 i_0_230 (.A1(n_0_32), .A2(n_0_6), .ZN(normalizedWires[525]));
   NOR2_X1 i_0_231 (.A1(n_0_32), .A2(n_0_7), .ZN(normalizedWires[526]));
   NOR2_X1 i_0_232 (.A1(n_0_32), .A2(n_0_8), .ZN(normalizedWires[527]));
   NOR2_X1 i_0_233 (.A1(n_0_32), .A2(n_0_9), .ZN(normalizedWires[528]));
   NOR2_X1 i_0_234 (.A1(n_0_32), .A2(n_0_10), .ZN(normalizedWires[529]));
   NOR2_X1 i_0_235 (.A1(n_0_32), .A2(n_0_11), .ZN(normalizedWires[530]));
   NOR2_X1 i_0_236 (.A1(n_0_32), .A2(n_0_12), .ZN(normalizedWires[531]));
   NOR2_X1 i_0_237 (.A1(n_0_32), .A2(n_0_13), .ZN(normalizedWires[532]));
   NOR2_X1 i_0_238 (.A1(n_0_32), .A2(n_0_14), .ZN(normalizedWires[533]));
   NOR2_X1 i_0_239 (.A1(n_0_32), .A2(n_0_15), .ZN(normalizedWires[534]));
   NOR2_X1 i_0_240 (.A1(n_0_32), .A2(n_0_16), .ZN(normalizedWires[535]));
   NOR2_X1 i_0_241 (.A1(n_0_32), .A2(n_0_17), .ZN(normalizedWires[536]));
   NOR2_X1 i_0_242 (.A1(n_0_32), .A2(n_0_18), .ZN(normalizedWires[537]));
   NOR2_X1 i_0_243 (.A1(n_0_32), .A2(n_0_19), .ZN(normalizedWires[538]));
   NOR2_X1 i_0_244 (.A1(n_0_32), .A2(n_0_20), .ZN(normalizedWires[539]));
   NOR2_X1 i_0_245 (.A1(n_0_32), .A2(n_0_21), .ZN(normalizedWires[540]));
   NOR2_X1 i_0_246 (.A1(n_0_32), .A2(n_0_22), .ZN(normalizedWires[541]));
   NOR2_X1 i_0_247 (.A1(n_0_32), .A2(n_0_23), .ZN(normalizedWires[542]));
   NOR2_X1 i_0_248 (.A1(n_0_32), .A2(n_0_24), .ZN(normalizedWires[543]));
   INV_X1 i_0_249 (.A(B[9]), .ZN(n_0_33));
   NOR2_X1 i_0_250 (.A1(n_0_33), .A2(n_0_1), .ZN(normalizedWires[585]));
   NOR2_X1 i_0_251 (.A1(n_0_33), .A2(n_0_2), .ZN(normalizedWires[586]));
   NOR2_X1 i_0_252 (.A1(n_0_33), .A2(n_0_3), .ZN(normalizedWires[587]));
   NOR2_X1 i_0_253 (.A1(n_0_33), .A2(n_0_4), .ZN(normalizedWires[588]));
   NOR2_X1 i_0_254 (.A1(n_0_33), .A2(n_0_5), .ZN(normalizedWires[589]));
   NOR2_X1 i_0_255 (.A1(n_0_33), .A2(n_0_6), .ZN(normalizedWires[590]));
   NOR2_X1 i_0_256 (.A1(n_0_33), .A2(n_0_7), .ZN(normalizedWires[591]));
   NOR2_X1 i_0_257 (.A1(n_0_33), .A2(n_0_8), .ZN(normalizedWires[592]));
   NOR2_X1 i_0_258 (.A1(n_0_33), .A2(n_0_9), .ZN(normalizedWires[593]));
   NOR2_X1 i_0_259 (.A1(n_0_33), .A2(n_0_10), .ZN(normalizedWires[594]));
   NOR2_X1 i_0_260 (.A1(n_0_33), .A2(n_0_11), .ZN(normalizedWires[595]));
   NOR2_X1 i_0_261 (.A1(n_0_33), .A2(n_0_12), .ZN(normalizedWires[596]));
   NOR2_X1 i_0_262 (.A1(n_0_33), .A2(n_0_13), .ZN(normalizedWires[597]));
   NOR2_X1 i_0_263 (.A1(n_0_33), .A2(n_0_14), .ZN(normalizedWires[598]));
   NOR2_X1 i_0_264 (.A1(n_0_33), .A2(n_0_15), .ZN(normalizedWires[599]));
   NOR2_X1 i_0_265 (.A1(n_0_33), .A2(n_0_16), .ZN(normalizedWires[600]));
   NOR2_X1 i_0_266 (.A1(n_0_33), .A2(n_0_17), .ZN(normalizedWires[601]));
   NOR2_X1 i_0_267 (.A1(n_0_33), .A2(n_0_18), .ZN(normalizedWires[602]));
   NOR2_X1 i_0_268 (.A1(n_0_33), .A2(n_0_19), .ZN(normalizedWires[603]));
   NOR2_X1 i_0_269 (.A1(n_0_33), .A2(n_0_20), .ZN(normalizedWires[604]));
   NOR2_X1 i_0_270 (.A1(n_0_33), .A2(n_0_21), .ZN(normalizedWires[605]));
   NOR2_X1 i_0_271 (.A1(n_0_33), .A2(n_0_22), .ZN(normalizedWires[606]));
   NOR2_X1 i_0_272 (.A1(n_0_33), .A2(n_0_23), .ZN(normalizedWires[607]));
   NOR2_X1 i_0_273 (.A1(n_0_33), .A2(n_0_24), .ZN(normalizedWires[608]));
   INV_X1 i_0_274 (.A(B[10]), .ZN(n_0_34));
   NOR2_X1 i_0_275 (.A1(n_0_34), .A2(n_0_1), .ZN(normalizedWires[650]));
   NOR2_X1 i_0_276 (.A1(n_0_34), .A2(n_0_2), .ZN(normalizedWires[651]));
   NOR2_X1 i_0_277 (.A1(n_0_34), .A2(n_0_3), .ZN(normalizedWires[652]));
   NOR2_X1 i_0_278 (.A1(n_0_34), .A2(n_0_4), .ZN(normalizedWires[653]));
   NOR2_X1 i_0_279 (.A1(n_0_34), .A2(n_0_5), .ZN(normalizedWires[654]));
   NOR2_X1 i_0_280 (.A1(n_0_34), .A2(n_0_6), .ZN(normalizedWires[655]));
   NOR2_X1 i_0_281 (.A1(n_0_34), .A2(n_0_7), .ZN(normalizedWires[656]));
   NOR2_X1 i_0_282 (.A1(n_0_34), .A2(n_0_8), .ZN(normalizedWires[657]));
   NOR2_X1 i_0_283 (.A1(n_0_34), .A2(n_0_9), .ZN(normalizedWires[658]));
   NOR2_X1 i_0_284 (.A1(n_0_34), .A2(n_0_10), .ZN(normalizedWires[659]));
   NOR2_X1 i_0_285 (.A1(n_0_34), .A2(n_0_11), .ZN(normalizedWires[660]));
   NOR2_X1 i_0_286 (.A1(n_0_34), .A2(n_0_12), .ZN(normalizedWires[661]));
   NOR2_X1 i_0_287 (.A1(n_0_34), .A2(n_0_13), .ZN(normalizedWires[662]));
   NOR2_X1 i_0_288 (.A1(n_0_34), .A2(n_0_14), .ZN(normalizedWires[663]));
   NOR2_X1 i_0_289 (.A1(n_0_34), .A2(n_0_15), .ZN(normalizedWires[664]));
   NOR2_X1 i_0_290 (.A1(n_0_34), .A2(n_0_16), .ZN(normalizedWires[665]));
   NOR2_X1 i_0_291 (.A1(n_0_34), .A2(n_0_17), .ZN(normalizedWires[666]));
   NOR2_X1 i_0_292 (.A1(n_0_34), .A2(n_0_18), .ZN(normalizedWires[667]));
   NOR2_X1 i_0_293 (.A1(n_0_34), .A2(n_0_19), .ZN(normalizedWires[668]));
   NOR2_X1 i_0_294 (.A1(n_0_34), .A2(n_0_20), .ZN(normalizedWires[669]));
   NOR2_X1 i_0_295 (.A1(n_0_34), .A2(n_0_21), .ZN(normalizedWires[670]));
   NOR2_X1 i_0_296 (.A1(n_0_34), .A2(n_0_22), .ZN(normalizedWires[671]));
   NOR2_X1 i_0_297 (.A1(n_0_34), .A2(n_0_23), .ZN(normalizedWires[672]));
   NOR2_X1 i_0_298 (.A1(n_0_34), .A2(n_0_24), .ZN(normalizedWires[673]));
   INV_X1 i_0_299 (.A(B[11]), .ZN(n_0_35));
   NOR2_X1 i_0_300 (.A1(n_0_35), .A2(n_0_1), .ZN(normalizedWires[715]));
   NOR2_X1 i_0_301 (.A1(n_0_35), .A2(n_0_2), .ZN(normalizedWires[716]));
   NOR2_X1 i_0_302 (.A1(n_0_35), .A2(n_0_3), .ZN(normalizedWires[717]));
   NOR2_X1 i_0_303 (.A1(n_0_35), .A2(n_0_4), .ZN(normalizedWires[718]));
   NOR2_X1 i_0_304 (.A1(n_0_35), .A2(n_0_5), .ZN(normalizedWires[719]));
   NOR2_X1 i_0_305 (.A1(n_0_35), .A2(n_0_6), .ZN(normalizedWires[720]));
   NOR2_X1 i_0_306 (.A1(n_0_35), .A2(n_0_7), .ZN(normalizedWires[721]));
   NOR2_X1 i_0_307 (.A1(n_0_35), .A2(n_0_8), .ZN(normalizedWires[722]));
   NOR2_X1 i_0_308 (.A1(n_0_35), .A2(n_0_9), .ZN(normalizedWires[723]));
   NOR2_X1 i_0_309 (.A1(n_0_35), .A2(n_0_10), .ZN(normalizedWires[724]));
   NOR2_X1 i_0_310 (.A1(n_0_35), .A2(n_0_11), .ZN(normalizedWires[725]));
   NOR2_X1 i_0_311 (.A1(n_0_35), .A2(n_0_12), .ZN(normalizedWires[726]));
   NOR2_X1 i_0_312 (.A1(n_0_35), .A2(n_0_13), .ZN(normalizedWires[727]));
   NOR2_X1 i_0_313 (.A1(n_0_35), .A2(n_0_14), .ZN(normalizedWires[728]));
   NOR2_X1 i_0_314 (.A1(n_0_35), .A2(n_0_15), .ZN(normalizedWires[729]));
   NOR2_X1 i_0_315 (.A1(n_0_35), .A2(n_0_16), .ZN(normalizedWires[730]));
   NOR2_X1 i_0_316 (.A1(n_0_35), .A2(n_0_17), .ZN(normalizedWires[731]));
   NOR2_X1 i_0_317 (.A1(n_0_35), .A2(n_0_18), .ZN(normalizedWires[732]));
   NOR2_X1 i_0_318 (.A1(n_0_35), .A2(n_0_19), .ZN(normalizedWires[733]));
   NOR2_X1 i_0_319 (.A1(n_0_35), .A2(n_0_20), .ZN(normalizedWires[734]));
   NOR2_X1 i_0_320 (.A1(n_0_35), .A2(n_0_21), .ZN(normalizedWires[735]));
   NOR2_X1 i_0_321 (.A1(n_0_35), .A2(n_0_22), .ZN(normalizedWires[736]));
   NOR2_X1 i_0_322 (.A1(n_0_35), .A2(n_0_23), .ZN(normalizedWires[737]));
   NOR2_X1 i_0_323 (.A1(n_0_35), .A2(n_0_24), .ZN(normalizedWires[738]));
   INV_X1 i_0_324 (.A(B[12]), .ZN(n_0_36));
   NOR2_X1 i_0_325 (.A1(n_0_36), .A2(n_0_1), .ZN(normalizedWires[780]));
   NOR2_X1 i_0_326 (.A1(n_0_36), .A2(n_0_2), .ZN(normalizedWires[781]));
   NOR2_X1 i_0_327 (.A1(n_0_36), .A2(n_0_3), .ZN(normalizedWires[782]));
   NOR2_X1 i_0_328 (.A1(n_0_36), .A2(n_0_4), .ZN(normalizedWires[783]));
   NOR2_X1 i_0_329 (.A1(n_0_36), .A2(n_0_5), .ZN(normalizedWires[784]));
   NOR2_X1 i_0_330 (.A1(n_0_36), .A2(n_0_6), .ZN(normalizedWires[785]));
   NOR2_X1 i_0_331 (.A1(n_0_36), .A2(n_0_7), .ZN(normalizedWires[786]));
   NOR2_X1 i_0_332 (.A1(n_0_36), .A2(n_0_8), .ZN(normalizedWires[787]));
   NOR2_X1 i_0_333 (.A1(n_0_36), .A2(n_0_9), .ZN(normalizedWires[788]));
   NOR2_X1 i_0_334 (.A1(n_0_36), .A2(n_0_10), .ZN(normalizedWires[789]));
   NOR2_X1 i_0_335 (.A1(n_0_36), .A2(n_0_11), .ZN(normalizedWires[790]));
   NOR2_X1 i_0_336 (.A1(n_0_36), .A2(n_0_12), .ZN(normalizedWires[791]));
   NOR2_X1 i_0_337 (.A1(n_0_36), .A2(n_0_13), .ZN(normalizedWires[792]));
   NOR2_X1 i_0_338 (.A1(n_0_36), .A2(n_0_14), .ZN(normalizedWires[793]));
   NOR2_X1 i_0_339 (.A1(n_0_36), .A2(n_0_15), .ZN(normalizedWires[794]));
   NOR2_X1 i_0_340 (.A1(n_0_36), .A2(n_0_16), .ZN(normalizedWires[795]));
   NOR2_X1 i_0_341 (.A1(n_0_36), .A2(n_0_17), .ZN(normalizedWires[796]));
   NOR2_X1 i_0_342 (.A1(n_0_36), .A2(n_0_18), .ZN(normalizedWires[797]));
   NOR2_X1 i_0_343 (.A1(n_0_36), .A2(n_0_19), .ZN(normalizedWires[798]));
   NOR2_X1 i_0_344 (.A1(n_0_36), .A2(n_0_20), .ZN(normalizedWires[799]));
   NOR2_X1 i_0_345 (.A1(n_0_36), .A2(n_0_21), .ZN(normalizedWires[800]));
   NOR2_X1 i_0_346 (.A1(n_0_36), .A2(n_0_22), .ZN(normalizedWires[801]));
   NOR2_X1 i_0_347 (.A1(n_0_36), .A2(n_0_23), .ZN(normalizedWires[802]));
   NOR2_X1 i_0_348 (.A1(n_0_36), .A2(n_0_24), .ZN(normalizedWires[803]));
   INV_X1 i_0_349 (.A(B[13]), .ZN(n_0_37));
   NOR2_X1 i_0_350 (.A1(n_0_37), .A2(n_0_1), .ZN(normalizedWires[845]));
   NOR2_X1 i_0_351 (.A1(n_0_37), .A2(n_0_2), .ZN(normalizedWires[846]));
   NOR2_X1 i_0_352 (.A1(n_0_37), .A2(n_0_3), .ZN(normalizedWires[847]));
   NOR2_X1 i_0_353 (.A1(n_0_37), .A2(n_0_4), .ZN(normalizedWires[848]));
   NOR2_X1 i_0_354 (.A1(n_0_37), .A2(n_0_5), .ZN(normalizedWires[849]));
   NOR2_X1 i_0_355 (.A1(n_0_37), .A2(n_0_6), .ZN(normalizedWires[850]));
   NOR2_X1 i_0_356 (.A1(n_0_37), .A2(n_0_7), .ZN(normalizedWires[851]));
   NOR2_X1 i_0_357 (.A1(n_0_37), .A2(n_0_8), .ZN(normalizedWires[852]));
   NOR2_X1 i_0_358 (.A1(n_0_37), .A2(n_0_9), .ZN(normalizedWires[853]));
   NOR2_X1 i_0_359 (.A1(n_0_37), .A2(n_0_10), .ZN(normalizedWires[854]));
   NOR2_X1 i_0_360 (.A1(n_0_37), .A2(n_0_11), .ZN(normalizedWires[855]));
   NOR2_X1 i_0_361 (.A1(n_0_37), .A2(n_0_12), .ZN(normalizedWires[856]));
   NOR2_X1 i_0_362 (.A1(n_0_37), .A2(n_0_13), .ZN(normalizedWires[857]));
   NOR2_X1 i_0_363 (.A1(n_0_37), .A2(n_0_14), .ZN(normalizedWires[858]));
   NOR2_X1 i_0_364 (.A1(n_0_37), .A2(n_0_15), .ZN(normalizedWires[859]));
   NOR2_X1 i_0_365 (.A1(n_0_37), .A2(n_0_16), .ZN(normalizedWires[860]));
   NOR2_X1 i_0_366 (.A1(n_0_37), .A2(n_0_17), .ZN(normalizedWires[861]));
   NOR2_X1 i_0_367 (.A1(n_0_37), .A2(n_0_18), .ZN(normalizedWires[862]));
   NOR2_X1 i_0_368 (.A1(n_0_37), .A2(n_0_19), .ZN(normalizedWires[863]));
   NOR2_X1 i_0_369 (.A1(n_0_37), .A2(n_0_20), .ZN(normalizedWires[864]));
   NOR2_X1 i_0_370 (.A1(n_0_37), .A2(n_0_21), .ZN(normalizedWires[865]));
   NOR2_X1 i_0_371 (.A1(n_0_37), .A2(n_0_22), .ZN(normalizedWires[866]));
   NOR2_X1 i_0_372 (.A1(n_0_37), .A2(n_0_23), .ZN(normalizedWires[867]));
   NOR2_X1 i_0_373 (.A1(n_0_37), .A2(n_0_24), .ZN(normalizedWires[868]));
   INV_X1 i_0_374 (.A(B[14]), .ZN(n_0_38));
   NOR2_X1 i_0_375 (.A1(n_0_38), .A2(n_0_1), .ZN(normalizedWires[910]));
   NOR2_X1 i_0_376 (.A1(n_0_38), .A2(n_0_2), .ZN(normalizedWires[911]));
   NOR2_X1 i_0_377 (.A1(n_0_38), .A2(n_0_3), .ZN(normalizedWires[912]));
   NOR2_X1 i_0_378 (.A1(n_0_38), .A2(n_0_4), .ZN(normalizedWires[913]));
   NOR2_X1 i_0_379 (.A1(n_0_38), .A2(n_0_5), .ZN(normalizedWires[914]));
   NOR2_X1 i_0_380 (.A1(n_0_38), .A2(n_0_6), .ZN(normalizedWires[915]));
   NOR2_X1 i_0_381 (.A1(n_0_38), .A2(n_0_7), .ZN(normalizedWires[916]));
   NOR2_X1 i_0_382 (.A1(n_0_38), .A2(n_0_8), .ZN(normalizedWires[917]));
   NOR2_X1 i_0_383 (.A1(n_0_38), .A2(n_0_9), .ZN(normalizedWires[918]));
   NOR2_X1 i_0_384 (.A1(n_0_38), .A2(n_0_10), .ZN(normalizedWires[919]));
   NOR2_X1 i_0_385 (.A1(n_0_38), .A2(n_0_11), .ZN(normalizedWires[920]));
   NOR2_X1 i_0_386 (.A1(n_0_38), .A2(n_0_12), .ZN(normalizedWires[921]));
   NOR2_X1 i_0_387 (.A1(n_0_38), .A2(n_0_13), .ZN(normalizedWires[922]));
   NOR2_X1 i_0_388 (.A1(n_0_38), .A2(n_0_14), .ZN(normalizedWires[923]));
   NOR2_X1 i_0_389 (.A1(n_0_38), .A2(n_0_15), .ZN(normalizedWires[924]));
   NOR2_X1 i_0_390 (.A1(n_0_38), .A2(n_0_16), .ZN(normalizedWires[925]));
   NOR2_X1 i_0_391 (.A1(n_0_38), .A2(n_0_17), .ZN(normalizedWires[926]));
   NOR2_X1 i_0_392 (.A1(n_0_38), .A2(n_0_18), .ZN(normalizedWires[927]));
   NOR2_X1 i_0_393 (.A1(n_0_38), .A2(n_0_19), .ZN(normalizedWires[928]));
   NOR2_X1 i_0_394 (.A1(n_0_38), .A2(n_0_20), .ZN(normalizedWires[929]));
   NOR2_X1 i_0_395 (.A1(n_0_38), .A2(n_0_21), .ZN(normalizedWires[930]));
   NOR2_X1 i_0_396 (.A1(n_0_38), .A2(n_0_22), .ZN(normalizedWires[931]));
   NOR2_X1 i_0_397 (.A1(n_0_38), .A2(n_0_23), .ZN(normalizedWires[932]));
   NOR2_X1 i_0_398 (.A1(n_0_38), .A2(n_0_24), .ZN(normalizedWires[933]));
   INV_X1 i_0_399 (.A(B[15]), .ZN(n_0_39));
   NOR2_X1 i_0_400 (.A1(n_0_39), .A2(n_0_1), .ZN(normalizedWires[975]));
   NOR2_X1 i_0_401 (.A1(n_0_39), .A2(n_0_2), .ZN(normalizedWires[976]));
   NOR2_X1 i_0_402 (.A1(n_0_39), .A2(n_0_3), .ZN(normalizedWires[977]));
   NOR2_X1 i_0_403 (.A1(n_0_39), .A2(n_0_4), .ZN(normalizedWires[978]));
   NOR2_X1 i_0_404 (.A1(n_0_39), .A2(n_0_5), .ZN(normalizedWires[979]));
   NOR2_X1 i_0_405 (.A1(n_0_39), .A2(n_0_6), .ZN(normalizedWires[980]));
   NOR2_X1 i_0_406 (.A1(n_0_39), .A2(n_0_7), .ZN(normalizedWires[981]));
   NOR2_X1 i_0_407 (.A1(n_0_39), .A2(n_0_8), .ZN(normalizedWires[982]));
   NOR2_X1 i_0_408 (.A1(n_0_39), .A2(n_0_9), .ZN(normalizedWires[983]));
   NOR2_X1 i_0_409 (.A1(n_0_39), .A2(n_0_10), .ZN(normalizedWires[984]));
   NOR2_X1 i_0_410 (.A1(n_0_39), .A2(n_0_11), .ZN(normalizedWires[985]));
   NOR2_X1 i_0_411 (.A1(n_0_39), .A2(n_0_12), .ZN(normalizedWires[986]));
   NOR2_X1 i_0_412 (.A1(n_0_39), .A2(n_0_13), .ZN(normalizedWires[987]));
   NOR2_X1 i_0_413 (.A1(n_0_39), .A2(n_0_14), .ZN(normalizedWires[988]));
   NOR2_X1 i_0_414 (.A1(n_0_39), .A2(n_0_15), .ZN(normalizedWires[989]));
   NOR2_X1 i_0_415 (.A1(n_0_39), .A2(n_0_16), .ZN(normalizedWires[990]));
   NOR2_X1 i_0_416 (.A1(n_0_39), .A2(n_0_17), .ZN(normalizedWires[991]));
   NOR2_X1 i_0_417 (.A1(n_0_39), .A2(n_0_18), .ZN(normalizedWires[992]));
   NOR2_X1 i_0_418 (.A1(n_0_39), .A2(n_0_19), .ZN(normalizedWires[993]));
   NOR2_X1 i_0_419 (.A1(n_0_39), .A2(n_0_20), .ZN(normalizedWires[994]));
   NOR2_X1 i_0_420 (.A1(n_0_39), .A2(n_0_21), .ZN(normalizedWires[995]));
   NOR2_X1 i_0_421 (.A1(n_0_39), .A2(n_0_22), .ZN(normalizedWires[996]));
   NOR2_X1 i_0_422 (.A1(n_0_39), .A2(n_0_23), .ZN(normalizedWires[997]));
   NOR2_X1 i_0_423 (.A1(n_0_39), .A2(n_0_24), .ZN(normalizedWires[998]));
   INV_X1 i_0_424 (.A(B[16]), .ZN(n_0_40));
   NOR2_X1 i_0_425 (.A1(n_0_40), .A2(n_0_1), .ZN(normalizedWires[1040]));
   NOR2_X1 i_0_426 (.A1(n_0_40), .A2(n_0_2), .ZN(normalizedWires[1041]));
   NOR2_X1 i_0_427 (.A1(n_0_40), .A2(n_0_3), .ZN(normalizedWires[1042]));
   NOR2_X1 i_0_428 (.A1(n_0_40), .A2(n_0_4), .ZN(normalizedWires[1043]));
   NOR2_X1 i_0_429 (.A1(n_0_40), .A2(n_0_5), .ZN(normalizedWires[1044]));
   NOR2_X1 i_0_430 (.A1(n_0_40), .A2(n_0_6), .ZN(normalizedWires[1045]));
   NOR2_X1 i_0_431 (.A1(n_0_40), .A2(n_0_7), .ZN(normalizedWires[1046]));
   NOR2_X1 i_0_432 (.A1(n_0_40), .A2(n_0_8), .ZN(normalizedWires[1047]));
   NOR2_X1 i_0_433 (.A1(n_0_40), .A2(n_0_9), .ZN(normalizedWires[1048]));
   NOR2_X1 i_0_434 (.A1(n_0_40), .A2(n_0_10), .ZN(normalizedWires[1049]));
   NOR2_X1 i_0_435 (.A1(n_0_40), .A2(n_0_11), .ZN(normalizedWires[1050]));
   NOR2_X1 i_0_436 (.A1(n_0_40), .A2(n_0_12), .ZN(normalizedWires[1051]));
   NOR2_X1 i_0_437 (.A1(n_0_40), .A2(n_0_13), .ZN(normalizedWires[1052]));
   NOR2_X1 i_0_438 (.A1(n_0_40), .A2(n_0_14), .ZN(normalizedWires[1053]));
   NOR2_X1 i_0_439 (.A1(n_0_40), .A2(n_0_15), .ZN(normalizedWires[1054]));
   NOR2_X1 i_0_440 (.A1(n_0_40), .A2(n_0_16), .ZN(normalizedWires[1055]));
   NOR2_X1 i_0_441 (.A1(n_0_40), .A2(n_0_17), .ZN(normalizedWires[1056]));
   NOR2_X1 i_0_442 (.A1(n_0_40), .A2(n_0_18), .ZN(normalizedWires[1057]));
   NOR2_X1 i_0_443 (.A1(n_0_40), .A2(n_0_19), .ZN(normalizedWires[1058]));
   NOR2_X1 i_0_444 (.A1(n_0_40), .A2(n_0_20), .ZN(normalizedWires[1059]));
   NOR2_X1 i_0_445 (.A1(n_0_40), .A2(n_0_21), .ZN(normalizedWires[1060]));
   NOR2_X1 i_0_446 (.A1(n_0_40), .A2(n_0_22), .ZN(normalizedWires[1061]));
   NOR2_X1 i_0_447 (.A1(n_0_40), .A2(n_0_23), .ZN(normalizedWires[1062]));
   NOR2_X1 i_0_448 (.A1(n_0_40), .A2(n_0_24), .ZN(normalizedWires[1063]));
   INV_X1 i_0_449 (.A(B[17]), .ZN(n_0_41));
   NOR2_X1 i_0_450 (.A1(n_0_41), .A2(n_0_1), .ZN(normalizedWires[1105]));
   NOR2_X1 i_0_451 (.A1(n_0_41), .A2(n_0_2), .ZN(normalizedWires[1106]));
   NOR2_X1 i_0_452 (.A1(n_0_41), .A2(n_0_3), .ZN(normalizedWires[1107]));
   NOR2_X1 i_0_453 (.A1(n_0_41), .A2(n_0_4), .ZN(normalizedWires[1108]));
   NOR2_X1 i_0_454 (.A1(n_0_41), .A2(n_0_5), .ZN(normalizedWires[1109]));
   NOR2_X1 i_0_455 (.A1(n_0_41), .A2(n_0_6), .ZN(normalizedWires[1110]));
   NOR2_X1 i_0_456 (.A1(n_0_41), .A2(n_0_7), .ZN(normalizedWires[1111]));
   NOR2_X1 i_0_457 (.A1(n_0_41), .A2(n_0_8), .ZN(normalizedWires[1112]));
   NOR2_X1 i_0_458 (.A1(n_0_41), .A2(n_0_9), .ZN(normalizedWires[1113]));
   NOR2_X1 i_0_459 (.A1(n_0_41), .A2(n_0_10), .ZN(normalizedWires[1114]));
   NOR2_X1 i_0_460 (.A1(n_0_41), .A2(n_0_11), .ZN(normalizedWires[1115]));
   NOR2_X1 i_0_461 (.A1(n_0_41), .A2(n_0_12), .ZN(normalizedWires[1116]));
   NOR2_X1 i_0_462 (.A1(n_0_41), .A2(n_0_13), .ZN(normalizedWires[1117]));
   NOR2_X1 i_0_463 (.A1(n_0_41), .A2(n_0_14), .ZN(normalizedWires[1118]));
   NOR2_X1 i_0_464 (.A1(n_0_41), .A2(n_0_15), .ZN(normalizedWires[1119]));
   NOR2_X1 i_0_465 (.A1(n_0_41), .A2(n_0_16), .ZN(normalizedWires[1120]));
   NOR2_X1 i_0_466 (.A1(n_0_41), .A2(n_0_17), .ZN(normalizedWires[1121]));
   NOR2_X1 i_0_467 (.A1(n_0_41), .A2(n_0_18), .ZN(normalizedWires[1122]));
   NOR2_X1 i_0_468 (.A1(n_0_41), .A2(n_0_19), .ZN(normalizedWires[1123]));
   NOR2_X1 i_0_469 (.A1(n_0_41), .A2(n_0_20), .ZN(normalizedWires[1124]));
   NOR2_X1 i_0_470 (.A1(n_0_41), .A2(n_0_21), .ZN(normalizedWires[1125]));
   NOR2_X1 i_0_471 (.A1(n_0_41), .A2(n_0_22), .ZN(normalizedWires[1126]));
   NOR2_X1 i_0_472 (.A1(n_0_41), .A2(n_0_23), .ZN(normalizedWires[1127]));
   NOR2_X1 i_0_473 (.A1(n_0_41), .A2(n_0_24), .ZN(normalizedWires[1128]));
   INV_X1 i_0_474 (.A(B[18]), .ZN(n_0_42));
   NOR2_X1 i_0_475 (.A1(n_0_42), .A2(n_0_1), .ZN(normalizedWires[1170]));
   NOR2_X1 i_0_476 (.A1(n_0_42), .A2(n_0_2), .ZN(normalizedWires[1171]));
   NOR2_X1 i_0_477 (.A1(n_0_42), .A2(n_0_3), .ZN(normalizedWires[1172]));
   NOR2_X1 i_0_478 (.A1(n_0_42), .A2(n_0_4), .ZN(normalizedWires[1173]));
   NOR2_X1 i_0_479 (.A1(n_0_42), .A2(n_0_5), .ZN(normalizedWires[1174]));
   NOR2_X1 i_0_480 (.A1(n_0_42), .A2(n_0_6), .ZN(normalizedWires[1175]));
   NOR2_X1 i_0_481 (.A1(n_0_42), .A2(n_0_7), .ZN(normalizedWires[1176]));
   NOR2_X1 i_0_482 (.A1(n_0_42), .A2(n_0_8), .ZN(normalizedWires[1177]));
   NOR2_X1 i_0_483 (.A1(n_0_42), .A2(n_0_9), .ZN(normalizedWires[1178]));
   NOR2_X1 i_0_484 (.A1(n_0_42), .A2(n_0_10), .ZN(normalizedWires[1179]));
   NOR2_X1 i_0_485 (.A1(n_0_42), .A2(n_0_11), .ZN(normalizedWires[1180]));
   NOR2_X1 i_0_486 (.A1(n_0_42), .A2(n_0_12), .ZN(normalizedWires[1181]));
   NOR2_X1 i_0_487 (.A1(n_0_42), .A2(n_0_13), .ZN(normalizedWires[1182]));
   NOR2_X1 i_0_488 (.A1(n_0_42), .A2(n_0_14), .ZN(normalizedWires[1183]));
   NOR2_X1 i_0_489 (.A1(n_0_42), .A2(n_0_15), .ZN(normalizedWires[1184]));
   NOR2_X1 i_0_490 (.A1(n_0_42), .A2(n_0_16), .ZN(normalizedWires[1185]));
   NOR2_X1 i_0_491 (.A1(n_0_42), .A2(n_0_17), .ZN(normalizedWires[1186]));
   NOR2_X1 i_0_492 (.A1(n_0_42), .A2(n_0_18), .ZN(normalizedWires[1187]));
   NOR2_X1 i_0_493 (.A1(n_0_42), .A2(n_0_19), .ZN(normalizedWires[1188]));
   NOR2_X1 i_0_494 (.A1(n_0_42), .A2(n_0_20), .ZN(normalizedWires[1189]));
   NOR2_X1 i_0_495 (.A1(n_0_42), .A2(n_0_21), .ZN(normalizedWires[1190]));
   NOR2_X1 i_0_496 (.A1(n_0_42), .A2(n_0_22), .ZN(normalizedWires[1191]));
   NOR2_X1 i_0_497 (.A1(n_0_42), .A2(n_0_23), .ZN(normalizedWires[1192]));
   NOR2_X1 i_0_498 (.A1(n_0_42), .A2(n_0_24), .ZN(normalizedWires[1193]));
   INV_X1 i_0_499 (.A(B[19]), .ZN(n_0_43));
   NOR2_X1 i_0_500 (.A1(n_0_43), .A2(n_0_1), .ZN(normalizedWires[1235]));
   NOR2_X1 i_0_501 (.A1(n_0_43), .A2(n_0_2), .ZN(normalizedWires[1236]));
   NOR2_X1 i_0_502 (.A1(n_0_43), .A2(n_0_3), .ZN(normalizedWires[1237]));
   NOR2_X1 i_0_503 (.A1(n_0_43), .A2(n_0_4), .ZN(normalizedWires[1238]));
   NOR2_X1 i_0_504 (.A1(n_0_43), .A2(n_0_5), .ZN(normalizedWires[1239]));
   NOR2_X1 i_0_505 (.A1(n_0_43), .A2(n_0_6), .ZN(normalizedWires[1240]));
   NOR2_X1 i_0_506 (.A1(n_0_43), .A2(n_0_7), .ZN(normalizedWires[1241]));
   NOR2_X1 i_0_507 (.A1(n_0_43), .A2(n_0_8), .ZN(normalizedWires[1242]));
   NOR2_X1 i_0_508 (.A1(n_0_43), .A2(n_0_9), .ZN(normalizedWires[1243]));
   NOR2_X1 i_0_509 (.A1(n_0_43), .A2(n_0_10), .ZN(normalizedWires[1244]));
   NOR2_X1 i_0_510 (.A1(n_0_43), .A2(n_0_11), .ZN(normalizedWires[1245]));
   NOR2_X1 i_0_511 (.A1(n_0_43), .A2(n_0_12), .ZN(normalizedWires[1246]));
   NOR2_X1 i_0_512 (.A1(n_0_43), .A2(n_0_13), .ZN(normalizedWires[1247]));
   NOR2_X1 i_0_513 (.A1(n_0_43), .A2(n_0_14), .ZN(normalizedWires[1248]));
   NOR2_X1 i_0_514 (.A1(n_0_43), .A2(n_0_15), .ZN(normalizedWires[1249]));
   NOR2_X1 i_0_515 (.A1(n_0_43), .A2(n_0_16), .ZN(normalizedWires[1250]));
   NOR2_X1 i_0_516 (.A1(n_0_43), .A2(n_0_17), .ZN(normalizedWires[1251]));
   NOR2_X1 i_0_517 (.A1(n_0_43), .A2(n_0_18), .ZN(normalizedWires[1252]));
   NOR2_X1 i_0_518 (.A1(n_0_43), .A2(n_0_19), .ZN(normalizedWires[1253]));
   NOR2_X1 i_0_519 (.A1(n_0_43), .A2(n_0_20), .ZN(normalizedWires[1254]));
   NOR2_X1 i_0_520 (.A1(n_0_43), .A2(n_0_21), .ZN(normalizedWires[1255]));
   NOR2_X1 i_0_521 (.A1(n_0_43), .A2(n_0_22), .ZN(normalizedWires[1256]));
   NOR2_X1 i_0_522 (.A1(n_0_43), .A2(n_0_23), .ZN(normalizedWires[1257]));
   NOR2_X1 i_0_523 (.A1(n_0_43), .A2(n_0_24), .ZN(normalizedWires[1258]));
   INV_X1 i_0_524 (.A(B[20]), .ZN(n_0_44));
   NOR2_X1 i_0_525 (.A1(n_0_44), .A2(n_0_1), .ZN(normalizedWires[1300]));
   NOR2_X1 i_0_526 (.A1(n_0_44), .A2(n_0_2), .ZN(normalizedWires[1301]));
   NOR2_X1 i_0_527 (.A1(n_0_44), .A2(n_0_3), .ZN(normalizedWires[1302]));
   NOR2_X1 i_0_528 (.A1(n_0_44), .A2(n_0_4), .ZN(normalizedWires[1303]));
   NOR2_X1 i_0_529 (.A1(n_0_44), .A2(n_0_5), .ZN(normalizedWires[1304]));
   NOR2_X1 i_0_530 (.A1(n_0_44), .A2(n_0_6), .ZN(normalizedWires[1305]));
   NOR2_X1 i_0_531 (.A1(n_0_44), .A2(n_0_7), .ZN(normalizedWires[1306]));
   NOR2_X1 i_0_532 (.A1(n_0_44), .A2(n_0_8), .ZN(normalizedWires[1307]));
   NOR2_X1 i_0_533 (.A1(n_0_44), .A2(n_0_9), .ZN(normalizedWires[1308]));
   NOR2_X1 i_0_534 (.A1(n_0_44), .A2(n_0_10), .ZN(normalizedWires[1309]));
   NOR2_X1 i_0_535 (.A1(n_0_44), .A2(n_0_11), .ZN(normalizedWires[1310]));
   NOR2_X1 i_0_536 (.A1(n_0_44), .A2(n_0_12), .ZN(normalizedWires[1311]));
   NOR2_X1 i_0_537 (.A1(n_0_44), .A2(n_0_13), .ZN(normalizedWires[1312]));
   NOR2_X1 i_0_538 (.A1(n_0_44), .A2(n_0_14), .ZN(normalizedWires[1313]));
   NOR2_X1 i_0_539 (.A1(n_0_44), .A2(n_0_15), .ZN(normalizedWires[1314]));
   NOR2_X1 i_0_540 (.A1(n_0_44), .A2(n_0_16), .ZN(normalizedWires[1315]));
   NOR2_X1 i_0_541 (.A1(n_0_44), .A2(n_0_17), .ZN(normalizedWires[1316]));
   NOR2_X1 i_0_542 (.A1(n_0_44), .A2(n_0_18), .ZN(normalizedWires[1317]));
   NOR2_X1 i_0_543 (.A1(n_0_44), .A2(n_0_19), .ZN(normalizedWires[1318]));
   NOR2_X1 i_0_544 (.A1(n_0_44), .A2(n_0_20), .ZN(normalizedWires[1319]));
   NOR2_X1 i_0_545 (.A1(n_0_44), .A2(n_0_21), .ZN(normalizedWires[1320]));
   NOR2_X1 i_0_546 (.A1(n_0_44), .A2(n_0_22), .ZN(normalizedWires[1321]));
   NOR2_X1 i_0_547 (.A1(n_0_44), .A2(n_0_23), .ZN(normalizedWires[1322]));
   NOR2_X1 i_0_548 (.A1(n_0_44), .A2(n_0_24), .ZN(normalizedWires[1323]));
   INV_X1 i_0_549 (.A(B[21]), .ZN(n_0_45));
   NOR2_X1 i_0_550 (.A1(n_0_45), .A2(n_0_1), .ZN(normalizedWires[1365]));
   NOR2_X1 i_0_551 (.A1(n_0_45), .A2(n_0_2), .ZN(normalizedWires[1366]));
   NOR2_X1 i_0_552 (.A1(n_0_45), .A2(n_0_3), .ZN(normalizedWires[1367]));
   NOR2_X1 i_0_553 (.A1(n_0_45), .A2(n_0_4), .ZN(normalizedWires[1368]));
   NOR2_X1 i_0_554 (.A1(n_0_45), .A2(n_0_5), .ZN(normalizedWires[1369]));
   NOR2_X1 i_0_555 (.A1(n_0_45), .A2(n_0_6), .ZN(normalizedWires[1370]));
   NOR2_X1 i_0_556 (.A1(n_0_45), .A2(n_0_7), .ZN(normalizedWires[1371]));
   NOR2_X1 i_0_557 (.A1(n_0_45), .A2(n_0_8), .ZN(normalizedWires[1372]));
   NOR2_X1 i_0_558 (.A1(n_0_45), .A2(n_0_9), .ZN(normalizedWires[1373]));
   NOR2_X1 i_0_559 (.A1(n_0_45), .A2(n_0_10), .ZN(normalizedWires[1374]));
   NOR2_X1 i_0_560 (.A1(n_0_45), .A2(n_0_11), .ZN(normalizedWires[1375]));
   NOR2_X1 i_0_561 (.A1(n_0_45), .A2(n_0_12), .ZN(normalizedWires[1376]));
   NOR2_X1 i_0_562 (.A1(n_0_45), .A2(n_0_13), .ZN(normalizedWires[1377]));
   NOR2_X1 i_0_563 (.A1(n_0_45), .A2(n_0_14), .ZN(normalizedWires[1378]));
   NOR2_X1 i_0_564 (.A1(n_0_45), .A2(n_0_15), .ZN(normalizedWires[1379]));
   NOR2_X1 i_0_565 (.A1(n_0_45), .A2(n_0_16), .ZN(normalizedWires[1380]));
   NOR2_X1 i_0_566 (.A1(n_0_45), .A2(n_0_17), .ZN(normalizedWires[1381]));
   NOR2_X1 i_0_567 (.A1(n_0_45), .A2(n_0_18), .ZN(normalizedWires[1382]));
   NOR2_X1 i_0_568 (.A1(n_0_45), .A2(n_0_19), .ZN(normalizedWires[1383]));
   NOR2_X1 i_0_569 (.A1(n_0_45), .A2(n_0_20), .ZN(normalizedWires[1384]));
   NOR2_X1 i_0_570 (.A1(n_0_45), .A2(n_0_21), .ZN(normalizedWires[1385]));
   NOR2_X1 i_0_571 (.A1(n_0_45), .A2(n_0_22), .ZN(normalizedWires[1386]));
   NOR2_X1 i_0_572 (.A1(n_0_45), .A2(n_0_23), .ZN(normalizedWires[1387]));
   NOR2_X1 i_0_573 (.A1(n_0_45), .A2(n_0_24), .ZN(normalizedWires[1388]));
   INV_X1 i_0_574 (.A(B[22]), .ZN(n_0_46));
   NOR2_X1 i_0_575 (.A1(n_0_46), .A2(n_0_1), .ZN(normalizedWires[1430]));
   NOR2_X1 i_0_576 (.A1(n_0_46), .A2(n_0_2), .ZN(normalizedWires[1431]));
   NOR2_X1 i_0_577 (.A1(n_0_46), .A2(n_0_3), .ZN(normalizedWires[1432]));
   NOR2_X1 i_0_578 (.A1(n_0_46), .A2(n_0_4), .ZN(normalizedWires[1433]));
   NOR2_X1 i_0_579 (.A1(n_0_46), .A2(n_0_5), .ZN(normalizedWires[1434]));
   NOR2_X1 i_0_580 (.A1(n_0_46), .A2(n_0_6), .ZN(normalizedWires[1435]));
   NOR2_X1 i_0_581 (.A1(n_0_46), .A2(n_0_7), .ZN(normalizedWires[1436]));
   NOR2_X1 i_0_582 (.A1(n_0_46), .A2(n_0_8), .ZN(normalizedWires[1437]));
   NOR2_X1 i_0_583 (.A1(n_0_46), .A2(n_0_9), .ZN(normalizedWires[1438]));
   NOR2_X1 i_0_584 (.A1(n_0_46), .A2(n_0_10), .ZN(normalizedWires[1439]));
   NOR2_X1 i_0_585 (.A1(n_0_46), .A2(n_0_11), .ZN(normalizedWires[1440]));
   NOR2_X1 i_0_586 (.A1(n_0_46), .A2(n_0_12), .ZN(normalizedWires[1441]));
   NOR2_X1 i_0_587 (.A1(n_0_46), .A2(n_0_13), .ZN(normalizedWires[1442]));
   NOR2_X1 i_0_588 (.A1(n_0_46), .A2(n_0_14), .ZN(normalizedWires[1443]));
   NOR2_X1 i_0_589 (.A1(n_0_46), .A2(n_0_15), .ZN(normalizedWires[1444]));
   NOR2_X1 i_0_590 (.A1(n_0_46), .A2(n_0_16), .ZN(normalizedWires[1445]));
   NOR2_X1 i_0_591 (.A1(n_0_46), .A2(n_0_17), .ZN(normalizedWires[1446]));
   NOR2_X1 i_0_592 (.A1(n_0_46), .A2(n_0_18), .ZN(normalizedWires[1447]));
   NOR2_X1 i_0_593 (.A1(n_0_46), .A2(n_0_19), .ZN(normalizedWires[1448]));
   NOR2_X1 i_0_594 (.A1(n_0_46), .A2(n_0_20), .ZN(normalizedWires[1449]));
   NOR2_X1 i_0_595 (.A1(n_0_46), .A2(n_0_21), .ZN(normalizedWires[1450]));
   NOR2_X1 i_0_596 (.A1(n_0_46), .A2(n_0_22), .ZN(normalizedWires[1451]));
   NOR2_X1 i_0_597 (.A1(n_0_46), .A2(n_0_23), .ZN(normalizedWires[1452]));
   NOR2_X1 i_0_598 (.A1(n_0_46), .A2(n_0_24), .ZN(normalizedWires[1453]));
   NOR2_X1 i_0_599 (.A1(n_0_1), .A2(n_0_24), .ZN(normalizedWires[1495]));
   NOR2_X1 i_0_600 (.A1(n_0_2), .A2(n_0_24), .ZN(normalizedWires[1496]));
   NOR2_X1 i_0_601 (.A1(n_0_3), .A2(n_0_24), .ZN(normalizedWires[1497]));
   NOR2_X1 i_0_602 (.A1(n_0_4), .A2(n_0_24), .ZN(normalizedWires[1498]));
   NOR2_X1 i_0_603 (.A1(n_0_5), .A2(n_0_24), .ZN(normalizedWires[1499]));
   NOR2_X1 i_0_604 (.A1(n_0_6), .A2(n_0_24), .ZN(normalizedWires[1500]));
   NOR2_X1 i_0_605 (.A1(n_0_7), .A2(n_0_24), .ZN(normalizedWires[1501]));
   NOR2_X1 i_0_606 (.A1(n_0_8), .A2(n_0_24), .ZN(normalizedWires[1502]));
   NOR2_X1 i_0_607 (.A1(n_0_9), .A2(n_0_24), .ZN(normalizedWires[1503]));
   NOR2_X1 i_0_608 (.A1(n_0_10), .A2(n_0_24), .ZN(normalizedWires[1504]));
   NOR2_X1 i_0_609 (.A1(n_0_11), .A2(n_0_24), .ZN(normalizedWires[1505]));
   NOR2_X1 i_0_610 (.A1(n_0_12), .A2(n_0_24), .ZN(normalizedWires[1506]));
   NOR2_X1 i_0_611 (.A1(n_0_13), .A2(n_0_24), .ZN(normalizedWires[1507]));
   NOR2_X1 i_0_612 (.A1(n_0_14), .A2(n_0_24), .ZN(normalizedWires[1508]));
   NOR2_X1 i_0_613 (.A1(n_0_15), .A2(n_0_24), .ZN(normalizedWires[1509]));
   NOR2_X1 i_0_614 (.A1(n_0_16), .A2(n_0_24), .ZN(normalizedWires[1510]));
   NOR2_X1 i_0_615 (.A1(n_0_17), .A2(n_0_24), .ZN(normalizedWires[1511]));
   NOR2_X1 i_0_616 (.A1(n_0_18), .A2(n_0_24), .ZN(normalizedWires[1512]));
   NOR2_X1 i_0_617 (.A1(n_0_19), .A2(n_0_24), .ZN(normalizedWires[1513]));
   NOR2_X1 i_0_618 (.A1(n_0_20), .A2(n_0_24), .ZN(normalizedWires[1514]));
   NOR2_X1 i_0_619 (.A1(n_0_21), .A2(n_0_24), .ZN(normalizedWires[1515]));
   NOR2_X1 i_0_620 (.A1(n_0_22), .A2(n_0_24), .ZN(normalizedWires[1516]));
   NOR2_X1 i_0_621 (.A1(n_0_24), .A2(n_0_23), .ZN(normalizedWires[1517]));
endmodule

module datapath(carry_in, Res_in, Res_out);
   input [63:0]carry_in;
   input [63:0]Res_in;
   output [63:0]Res_out;

   XOR2_X1 i_0 (.A(n_4), .B(n_1), .Z(Res_out[24]));
   OAI21_X1 i_1 (.A(n_3), .B1(n_147), .B2(n_137), .ZN(n_1));
   NOR2_X1 i_2 (.A1(n_146), .A2(n_138), .ZN(n_4));
   XOR2_X1 i_3 (.A(n_135), .B(n_11), .Z(Res_out[25]));
   XOR2_X1 i_4 (.A(n_10), .B(n_7), .Z(Res_out[26]));
   XOR2_X1 i_5 (.A(n_8), .B(n_5), .Z(Res_out[27]));
   NOR2_X1 i_6 (.A1(n_106), .A2(n_73), .ZN(n_5));
   XNOR2_X1 i_7 (.A(n_12), .B(n_6), .ZN(Res_out[28]));
   OAI21_X1 i_8 (.A(n_105), .B1(n_73), .B2(n_8), .ZN(n_6));
   NOR2_X1 i_9 (.A1(n_108), .A2(n_75), .ZN(n_7));
   INV_X1 i_10 (.A(n_9), .ZN(n_8));
   OAI21_X1 i_11 (.A(n_107), .B1(n_75), .B2(n_10), .ZN(n_9));
   AOI21_X1 i_12 (.A(n_103), .B1(n_135), .B2(n_77), .ZN(n_10));
   OAI21_X1 i_13 (.A(n_77), .B1(carry_in[25]), .B2(Res_in[25]), .ZN(n_11));
   AOI21_X1 i_14 (.A(n_110), .B1(carry_in[28]), .B2(Res_in[28]), .ZN(n_12));
   XOR2_X1 i_15 (.A(n_40), .B(n_19), .Z(Res_out[29]));
   XOR2_X1 i_16 (.A(n_18), .B(n_15), .Z(Res_out[30]));
   XOR2_X1 i_17 (.A(n_16), .B(n_13), .Z(Res_out[31]));
   NOR2_X1 i_18 (.A1(n_122), .A2(n_89), .ZN(n_13));
   XNOR2_X1 i_19 (.A(n_20), .B(n_14), .ZN(Res_out[32]));
   OAI21_X1 i_20 (.A(n_121), .B1(n_89), .B2(n_16), .ZN(n_14));
   NOR2_X1 i_21 (.A1(n_124), .A2(n_91), .ZN(n_15));
   INV_X1 i_22 (.A(n_17), .ZN(n_16));
   OAI21_X1 i_23 (.A(n_123), .B1(n_91), .B2(n_18), .ZN(n_17));
   AOI21_X1 i_24 (.A(n_127), .B1(n_93), .B2(n_40), .ZN(n_18));
   OAI21_X1 i_25 (.A(n_93), .B1(carry_in[29]), .B2(Res_in[29]), .ZN(n_19));
   AOI21_X1 i_26 (.A(n_126), .B1(carry_in[32]), .B2(Res_in[32]), .ZN(n_20));
   XNOR2_X1 i_27 (.A(n_29), .B(n_28), .ZN(Res_out[33]));
   XOR2_X1 i_28 (.A(n_26), .B(n_25), .Z(Res_out[34]));
   XNOR2_X1 i_29 (.A(n_22), .B(n_21), .ZN(Res_out[35]));
   OAI22_X1 i_30 (.A1(carry_in[34]), .A2(Res_in[34]), .B1(n_98), .B2(n_26), 
      .ZN(n_21));
   NOR2_X1 i_31 (.A1(n_116), .A2(n_95), .ZN(n_22));
   XNOR2_X1 i_32 (.A(n_30), .B(n_23), .ZN(Res_out[36]));
   OAI21_X1 i_33 (.A(n_24), .B1(n_115), .B2(n_95), .ZN(n_23));
   NAND3_X1 i_34 (.A1(n_96), .A2(n_25), .A3(n_27), .ZN(n_24));
   NOR2_X1 i_35 (.A1(n_117), .A2(n_98), .ZN(n_25));
   INV_X1 i_36 (.A(n_27), .ZN(n_26));
   OAI22_X1 i_37 (.A1(carry_in[33]), .A2(Res_in[33]), .B1(n_99), .B2(n_29), 
      .ZN(n_27));
   OAI21_X1 i_38 (.A(n_100), .B1(carry_in[33]), .B2(Res_in[33]), .ZN(n_28));
   OAI21_X1 i_39 (.A(n_88), .B1(n_119), .B2(n_40), .ZN(n_29));
   AOI21_X1 i_40 (.A(n_118), .B1(carry_in[36]), .B2(Res_in[36]), .ZN(n_30));
   XNOR2_X1 i_41 (.A(n_39), .B(n_38), .ZN(Res_out[37]));
   XOR2_X1 i_42 (.A(n_36), .B(n_35), .Z(Res_out[38]));
   XNOR2_X1 i_43 (.A(n_32), .B(n_31), .ZN(Res_out[39]));
   OAI22_X1 i_44 (.A1(carry_in[38]), .A2(Res_in[38]), .B1(n_83), .B2(n_36), 
      .ZN(n_31));
   NOR2_X1 i_45 (.A1(n_131), .A2(n_80), .ZN(n_32));
   XNOR2_X1 i_50 (.A(n_42), .B(n_33), .ZN(Res_out[40]));
   OAI21_X1 i_51 (.A(n_34), .B1(n_130), .B2(n_80), .ZN(n_33));
   NAND3_X1 i_52 (.A1(n_81), .A2(n_35), .A3(n_37), .ZN(n_34));
   NOR2_X1 i_46 (.A1(n_132), .A2(n_83), .ZN(n_35));
   INV_X1 i_47 (.A(n_37), .ZN(n_36));
   OAI22_X1 i_48 (.A1(carry_in[37]), .A2(Res_in[37]), .B1(n_84), .B2(n_39), 
      .ZN(n_37));
   OAI21_X1 i_49 (.A(n_85), .B1(carry_in[37]), .B2(Res_in[37]), .ZN(n_38));
   OAI21_X1 i_53 (.A(n_86), .B1(n_112), .B2(n_40), .ZN(n_39));
   INV_X1 i_54 (.A(n_41), .ZN(n_40));
   OAI21_X1 i_55 (.A(n_72), .B1(n_135), .B2(n_102), .ZN(n_41));
   AOI21_X1 i_60 (.A(n_133), .B1(carry_in[40]), .B2(Res_in[40]), .ZN(n_42));
   XOR2_X1 i_61 (.A(n_70), .B(n_49), .Z(Res_out[41]));
   XOR2_X1 i_62 (.A(n_48), .B(n_45), .Z(Res_out[42]));
   XOR2_X1 i_63 (.A(n_46), .B(n_43), .Z(Res_out[43]));
   NOR2_X1 i_64 (.A1(n_66), .A2(n_58), .ZN(n_43));
   XNOR2_X1 i_65 (.A(n_50), .B(n_44), .ZN(Res_out[44]));
   OAI22_X1 i_66 (.A1(carry_in[43]), .A2(Res_in[43]), .B1(n_58), .B2(n_46), 
      .ZN(n_44));
   AOI21_X1 i_67 (.A(n_67), .B1(carry_in[42]), .B2(Res_in[42]), .ZN(n_45));
   AOI21_X1 i_68 (.A(n_67), .B1(n_62), .B2(n_47), .ZN(n_46));
   INV_X1 i_69 (.A(n_48), .ZN(n_47));
   AOI21_X1 i_70 (.A(n_69), .B1(n_70), .B2(n_63), .ZN(n_48));
   OAI21_X1 i_71 (.A(n_63), .B1(carry_in[41]), .B2(Res_in[41]), .ZN(n_49));
   NOR2_X1 i_72 (.A1(n_68), .A2(n_60), .ZN(n_50));
   XOR2_X1 i_73 (.A(n_56), .B(n_51), .Z(Res_out[45]));
   OAI22_X1 i_74 (.A1(carry_in[45]), .A2(Res_in[45]), .B1(n_175), .B2(n_173), 
      .ZN(n_51));
   XNOR2_X1 i_75 (.A(n_55), .B(n_52), .ZN(Res_out[46]));
   OAI21_X1 i_76 (.A(n_172), .B1(n_0), .B2(n_174), .ZN(n_52));
   XNOR2_X1 i_77 (.A(n_54), .B(n_53), .ZN(Res_out[47]));
   XOR2_X1 i_78 (.A(carry_in[47]), .B(Res_in[47]), .Z(n_53));
   AOI22_X1 i_79 (.A1(carry_in[46]), .A2(Res_in[46]), .B1(n_172), .B2(n_55), 
      .ZN(n_54));
   OAI22_X1 i_80 (.A1(n_175), .A2(n_173), .B1(n_171), .B2(n_56), .ZN(n_55));
   NOR4_X1 i_81 (.A1(n_60), .A2(n_57), .A3(n_61), .A4(n_64), .ZN(n_56));
   NOR2_X1 i_56 (.A1(n_68), .A2(n_59), .ZN(n_57));
   INV_X1 i_83 (.A(n_59), .ZN(n_58));
   NAND2_X1 i_57 (.A1(carry_in[43]), .A2(Res_in[43]), .ZN(n_59));
   AND2_X1 i_85 (.A1(carry_in[44]), .A2(Res_in[44]), .ZN(n_60));
   AOI21_X1 i_58 (.A(n_65), .B1(n_63), .B2(n_62), .ZN(n_61));
   NAND2_X1 i_59 (.A1(carry_in[42]), .A2(Res_in[42]), .ZN(n_62));
   NAND2_X1 i_82 (.A1(carry_in[41]), .A2(Res_in[41]), .ZN(n_63));
   NOR3_X1 i_89 (.A1(n_69), .A2(n_65), .A3(n_70), .ZN(n_64));
   OR3_X1 i_84 (.A1(n_68), .A2(n_66), .A3(n_67), .ZN(n_65));
   NOR2_X1 i_86 (.A1(carry_in[43]), .A2(Res_in[43]), .ZN(n_66));
   NOR2_X1 i_87 (.A1(carry_in[42]), .A2(Res_in[42]), .ZN(n_67));
   NOR2_X1 i_88 (.A1(carry_in[44]), .A2(Res_in[44]), .ZN(n_68));
   NOR2_X1 i_94 (.A1(carry_in[41]), .A2(Res_in[41]), .ZN(n_69));
   AOI21_X1 i_95 (.A(n_71), .B1(n_134), .B2(n_101), .ZN(n_70));
   OAI221_X1 i_90 (.A(n_78), .B1(n_111), .B2(n_72), .C1(n_128), .C2(n_86), 
      .ZN(n_71));
   AOI221_X1 i_91 (.A(n_74), .B1(carry_in[28]), .B2(Res_in[28]), .C1(n_109), 
      .C2(n_73), .ZN(n_72));
   AND2_X1 i_92 (.A1(carry_in[27]), .A2(Res_in[27]), .ZN(n_73));
   AOI21_X1 i_93 (.A(n_104), .B1(n_77), .B2(n_76), .ZN(n_74));
   INV_X1 i_96 (.A(n_76), .ZN(n_75));
   NAND2_X1 i_97 (.A1(carry_in[26]), .A2(Res_in[26]), .ZN(n_76));
   NAND2_X1 i_98 (.A1(carry_in[25]), .A2(Res_in[25]), .ZN(n_77));
   AOI21_X1 i_99 (.A(n_79), .B1(carry_in[40]), .B2(Res_in[40]), .ZN(n_78));
   OAI21_X1 i_100 (.A(n_82), .B1(n_133), .B2(n_81), .ZN(n_79));
   INV_X1 i_101 (.A(n_81), .ZN(n_80));
   NAND2_X1 i_102 (.A1(carry_in[39]), .A2(Res_in[39]), .ZN(n_81));
   OAI21_X1 i_103 (.A(n_129), .B1(n_84), .B2(n_83), .ZN(n_82));
   AND2_X1 i_104 (.A1(carry_in[38]), .A2(Res_in[38]), .ZN(n_83));
   INV_X1 i_105 (.A(n_85), .ZN(n_84));
   NAND2_X1 i_106 (.A1(carry_in[37]), .A2(Res_in[37]), .ZN(n_85));
   AOI211_X1 i_107 (.A(n_94), .B(n_87), .C1(carry_in[36]), .C2(Res_in[36]), 
      .ZN(n_86));
   NOR2_X1 i_108 (.A1(n_113), .A2(n_88), .ZN(n_87));
   AOI221_X1 i_109 (.A(n_90), .B1(carry_in[32]), .B2(Res_in[32]), .C1(n_125), 
      .C2(n_89), .ZN(n_88));
   AND2_X1 i_110 (.A1(carry_in[31]), .A2(Res_in[31]), .ZN(n_89));
   AOI21_X1 i_111 (.A(n_120), .B1(n_93), .B2(n_92), .ZN(n_90));
   INV_X1 i_112 (.A(n_92), .ZN(n_91));
   NAND2_X1 i_113 (.A1(carry_in[30]), .A2(Res_in[30]), .ZN(n_92));
   NAND2_X1 i_114 (.A1(carry_in[29]), .A2(Res_in[29]), .ZN(n_93));
   OAI21_X1 i_115 (.A(n_97), .B1(n_118), .B2(n_96), .ZN(n_94));
   INV_X1 i_116 (.A(n_96), .ZN(n_95));
   NAND2_X1 i_117 (.A1(carry_in[35]), .A2(Res_in[35]), .ZN(n_96));
   OAI21_X1 i_118 (.A(n_114), .B1(n_99), .B2(n_98), .ZN(n_97));
   AND2_X1 i_119 (.A1(carry_in[34]), .A2(Res_in[34]), .ZN(n_98));
   INV_X1 i_120 (.A(n_100), .ZN(n_99));
   NAND2_X1 i_121 (.A1(carry_in[33]), .A2(Res_in[33]), .ZN(n_100));
   NOR2_X1 i_126 (.A1(n_111), .A2(n_102), .ZN(n_101));
   OR2_X1 i_122 (.A1(n_104), .A2(n_103), .ZN(n_102));
   NOR2_X1 i_123 (.A1(carry_in[25]), .A2(Res_in[25]), .ZN(n_103));
   NAND3_X1 i_124 (.A1(n_109), .A2(n_105), .A3(n_107), .ZN(n_104));
   INV_X1 i_125 (.A(n_106), .ZN(n_105));
   NOR2_X1 i_127 (.A1(carry_in[27]), .A2(Res_in[27]), .ZN(n_106));
   INV_X1 i_128 (.A(n_108), .ZN(n_107));
   NOR2_X1 i_129 (.A1(carry_in[26]), .A2(Res_in[26]), .ZN(n_108));
   INV_X1 i_130 (.A(n_110), .ZN(n_109));
   NOR2_X1 i_131 (.A1(carry_in[28]), .A2(Res_in[28]), .ZN(n_110));
   OR2_X1 i_132 (.A1(n_128), .A2(n_112), .ZN(n_111));
   OR2_X1 i_133 (.A1(n_119), .A2(n_113), .ZN(n_112));
   OAI21_X1 i_134 (.A(n_114), .B1(carry_in[33]), .B2(Res_in[33]), .ZN(n_113));
   NOR3_X1 i_135 (.A1(n_118), .A2(n_116), .A3(n_117), .ZN(n_114));
   NOR2_X1 i_136 (.A1(n_117), .A2(n_116), .ZN(n_115));
   NOR2_X1 i_137 (.A1(carry_in[35]), .A2(Res_in[35]), .ZN(n_116));
   NOR2_X1 i_138 (.A1(carry_in[34]), .A2(Res_in[34]), .ZN(n_117));
   NOR2_X1 i_139 (.A1(carry_in[36]), .A2(Res_in[36]), .ZN(n_118));
   OR2_X1 i_140 (.A1(n_127), .A2(n_120), .ZN(n_119));
   NAND3_X1 i_141 (.A1(n_125), .A2(n_121), .A3(n_123), .ZN(n_120));
   INV_X1 i_142 (.A(n_122), .ZN(n_121));
   NOR2_X1 i_143 (.A1(carry_in[31]), .A2(Res_in[31]), .ZN(n_122));
   INV_X1 i_144 (.A(n_124), .ZN(n_123));
   NOR2_X1 i_145 (.A1(carry_in[30]), .A2(Res_in[30]), .ZN(n_124));
   INV_X1 i_146 (.A(n_126), .ZN(n_125));
   NOR2_X1 i_147 (.A1(carry_in[32]), .A2(Res_in[32]), .ZN(n_126));
   NOR2_X1 i_148 (.A1(carry_in[29]), .A2(Res_in[29]), .ZN(n_127));
   OAI21_X1 i_149 (.A(n_129), .B1(carry_in[37]), .B2(Res_in[37]), .ZN(n_128));
   NOR3_X1 i_150 (.A1(n_133), .A2(n_131), .A3(n_132), .ZN(n_129));
   NOR2_X1 i_155 (.A1(n_132), .A2(n_131), .ZN(n_130));
   NOR2_X1 i_151 (.A1(carry_in[39]), .A2(Res_in[39]), .ZN(n_131));
   NOR2_X1 i_152 (.A1(carry_in[38]), .A2(Res_in[38]), .ZN(n_132));
   NOR2_X1 i_153 (.A1(carry_in[40]), .A2(Res_in[40]), .ZN(n_133));
   INV_X1 i_159 (.A(n_135), .ZN(n_134));
   NOR4_X1 i_154 (.A1(n_138), .A2(n_136), .A3(n_139), .A4(n_143), .ZN(n_135));
   NOR2_X1 i_156 (.A1(n_146), .A2(n_3), .ZN(n_136));
   AND2_X1 i_157 (.A1(carry_in[24]), .A2(Res_in[24]), .ZN(n_138));
   AOI21_X1 i_158 (.A(n_145), .B1(n_141), .B2(n_162), .ZN(n_139));
   NOR3_X1 i_160 (.A1(n_145), .A2(n_161), .A3(n_142), .ZN(n_143));
   OAI221_X1 i_161 (.A(n_164), .B1(carry_in[23]), .B2(Res_in[23]), .C1(
      carry_in[24]), .C2(Res_in[24]), .ZN(n_145));
   NOR2_X1 i_162 (.A1(carry_in[24]), .A2(Res_in[24]), .ZN(n_146));
   NOR2_X1 i_163 (.A1(carry_in[23]), .A2(Res_in[23]), .ZN(n_147));
   NOR2_X1 i_196 (.A1(carry_in[45]), .A2(Res_in[45]), .ZN(n_171));
   NAND2_X1 i_164 (.A1(n_0), .A2(n_174), .ZN(n_172));
   INV_X1 i_198 (.A(Res_in[45]), .ZN(n_173));
   INV_X1 i_165 (.A(Res_in[46]), .ZN(n_174));
   INV_X1 i_200 (.A(carry_in[45]), .ZN(n_175));
   INV_X1 i_166 (.A(carry_in[46]), .ZN(n_0));
   XOR2_X1 i_167 (.A(n_137), .B(n_2), .Z(Res_out[23]));
   OAI21_X1 i_168 (.A(n_3), .B1(carry_in[23]), .B2(Res_in[23]), .ZN(n_2));
   NAND2_X1 i_169 (.A1(carry_in[23]), .A2(Res_in[23]), .ZN(n_3));
   OAI21_X1 i_170 (.A(n_164), .B1(n_163), .B2(n_140), .ZN(n_137));
   AOI21_X1 i_171 (.A(n_161), .B1(n_142), .B2(n_141), .ZN(n_140));
   NAND2_X1 i_172 (.A1(carry_in[21]), .A2(Res_in[21]), .ZN(n_141));
   INV_X1 i_173 (.A(n_144), .ZN(n_142));
   OAI21_X1 i_174 (.A(n_149), .B1(n_151), .B2(n_148), .ZN(n_144));
   AOI22_X1 i_175 (.A1(carry_in[20]), .A2(Res_in[20]), .B1(carry_in[19]), 
      .B2(Res_in[19]), .ZN(n_148));
   OR3_X1 i_176 (.A1(n_151), .A2(n_150), .A3(n_152), .ZN(n_149));
   OAI22_X1 i_177 (.A1(carry_in[18]), .A2(Res_in[18]), .B1(carry_in[19]), 
      .B2(Res_in[19]), .ZN(n_150));
   NOR2_X1 i_178 (.A1(carry_in[20]), .A2(Res_in[20]), .ZN(n_151));
   AOI221_X1 i_179 (.A(n_153), .B1(carry_in[18]), .B2(Res_in[18]), .C1(
      carry_in[17]), .C2(Res_in[17]), .ZN(n_152));
   AOI21_X1 i_180 (.A(n_154), .B1(n_160), .B2(n_155), .ZN(n_153));
   OAI22_X1 i_181 (.A1(carry_in[17]), .A2(Res_in[17]), .B1(carry_in[16]), 
      .B2(Res_in[16]), .ZN(n_154));
   OAI221_X1 i_182 (.A(n_156), .B1(carry_in[14]), .B2(Res_in[14]), .C1(
      carry_in[15]), .C2(Res_in[15]), .ZN(n_155));
   OAI21_X1 i_183 (.A(n_159), .B1(n_158), .B2(n_157), .ZN(n_156));
   OAI22_X1 i_184 (.A1(carry_in[12]), .A2(Res_in[12]), .B1(carry_in[13]), 
      .B2(Res_in[13]), .ZN(n_157));
   AOI221_X1 i_185 (.A(n_165), .B1(carry_in[11]), .B2(Res_in[11]), .C1(
      carry_in[12]), .C2(Res_in[12]), .ZN(n_158));
   AOI22_X1 i_186 (.A1(carry_in[13]), .A2(Res_in[13]), .B1(carry_in[14]), 
      .B2(Res_in[14]), .ZN(n_159));
   AOI22_X1 i_187 (.A1(carry_in[16]), .A2(Res_in[16]), .B1(carry_in[15]), 
      .B2(Res_in[15]), .ZN(n_160));
   NOR2_X1 i_188 (.A1(carry_in[21]), .A2(Res_in[21]), .ZN(n_161));
   INV_X1 i_189 (.A(n_163), .ZN(n_162));
   NOR2_X1 i_190 (.A1(n_167), .A2(n_166), .ZN(n_163));
   NAND2_X1 i_191 (.A1(n_167), .A2(n_166), .ZN(n_164));
   INV_X1 i_192 (.A(n_168), .ZN(n_165));
   INV_X1 i_193 (.A(Res_in[22]), .ZN(n_166));
   INV_X1 i_194 (.A(carry_in[22]), .ZN(n_167));
   OAI221_X1 i_195 (.A(n_169), .B1(carry_in[11]), .B2(Res_in[11]), .C1(
      carry_in[10]), .C2(Res_in[10]), .ZN(n_168));
   INV_X1 i_197 (.A(n_170), .ZN(n_169));
   AOI22_X1 i_199 (.A1(carry_in[9]), .A2(Res_in[9]), .B1(carry_in[10]), .B2(
      Res_in[10]), .ZN(n_170));
endmodule

module addResWithCarry(Res_out, Res_in, carry_in);
   output [63:0]Res_out;
   input [63:0]Res_in;
   input [63:0]carry_in;

   datapath i_0 (.carry_in({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, 
      uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, carry_in[47], carry_in[46], 
      carry_in[45], carry_in[44], carry_in[43], carry_in[42], carry_in[41], 
      carry_in[40], carry_in[39], carry_in[38], carry_in[37], carry_in[36], 
      carry_in[35], carry_in[34], carry_in[33], carry_in[32], carry_in[31], 
      carry_in[30], carry_in[29], carry_in[28], carry_in[27], carry_in[26], 
      carry_in[25], carry_in[24], carry_in[23], carry_in[22], carry_in[21], 
      carry_in[20], carry_in[19], carry_in[18], carry_in[17], carry_in[16], 
      carry_in[15], carry_in[14], carry_in[13], carry_in[12], carry_in[11], 
      carry_in[10], carry_in[9], uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, 
      uc_23, uc_24}), .Res_in({uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, 
      uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, Res_in[47], 
      Res_in[46], Res_in[45], Res_in[44], Res_in[43], Res_in[42], Res_in[41], 
      Res_in[40], Res_in[39], Res_in[38], Res_in[37], Res_in[36], Res_in[35], 
      Res_in[34], Res_in[33], Res_in[32], Res_in[31], Res_in[30], Res_in[29], 
      Res_in[28], Res_in[27], Res_in[26], Res_in[25], Res_in[24], Res_in[23], 
      Res_in[22], Res_in[21], Res_in[20], Res_in[19], Res_in[18], Res_in[17], 
      Res_in[16], Res_in[15], Res_in[14], Res_in[13], Res_in[12], Res_in[11], 
      Res_in[10], Res_in[9], uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, 
      uc_48, uc_49}), .Res_out({uc_50, uc_51, uc_52, uc_53, uc_54, uc_55, uc_56, 
      uc_57, uc_58, uc_59, uc_60, uc_61, uc_62, uc_63, uc_64, uc_65, Res_out[47], 
      Res_out[46], Res_out[45], Res_out[44], Res_out[43], Res_out[42], 
      Res_out[41], Res_out[40], Res_out[39], Res_out[38], Res_out[37], 
      Res_out[36], Res_out[35], Res_out[34], Res_out[33], Res_out[32], 
      Res_out[31], Res_out[30], Res_out[29], Res_out[28], Res_out[27], 
      Res_out[26], Res_out[25], Res_out[24], Res_out[23], uc_66, uc_67, uc_68, 
      uc_69, uc_70, uc_71, uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, 
      uc_79, uc_80, uc_81, uc_82, uc_83, uc_84, uc_85, uc_86, uc_87, uc_88}));
endmodule

module multiplierTree(Res, OVF, A, B, clk, reset, enable);
   output [63:0]Res;
   output OVF;
   input [31:0]A;
   input [31:0]B;
   input clk;
   input reset;
   input enable;

   wire [63:0]secondStage_carry;
   wire [63:0]secondStage_Res;
   wire [2047:0]normalizedWires;
   wire [63:0]Res_imm;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_0;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_1;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_0_0;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_119;
   wire n_0_118;

   addIntermedaiteWires secondStage (.Res({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, 
      uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, 
      secondStage_Res[47], secondStage_Res[46], secondStage_Res[45], 
      secondStage_Res[44], secondStage_Res[43], secondStage_Res[42], 
      secondStage_Res[41], secondStage_Res[40], secondStage_Res[39], 
      secondStage_Res[38], secondStage_Res[37], secondStage_Res[36], 
      secondStage_Res[35], secondStage_Res[34], secondStage_Res[33], 
      secondStage_Res[32], secondStage_Res[31], secondStage_Res[30], 
      secondStage_Res[29], secondStage_Res[28], secondStage_Res[27], 
      secondStage_Res[26], secondStage_Res[25], secondStage_Res[24], 
      secondStage_Res[23], secondStage_Res[22], secondStage_Res[21], 
      secondStage_Res[20], secondStage_Res[19], secondStage_Res[18], 
      secondStage_Res[17], secondStage_Res[16], secondStage_Res[15], 
      secondStage_Res[14], secondStage_Res[13], secondStage_Res[12], 
      secondStage_Res[11], secondStage_Res[10], secondStage_Res[9], uc_16, uc_17, 
      uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24}), .carry({uc_25, uc_26, 
      uc_27, uc_28, uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, 
      uc_37, uc_38, uc_39, uc_40, secondStage_carry[47], secondStage_carry[46], 
      secondStage_carry[45], secondStage_carry[44], secondStage_carry[43], 
      secondStage_carry[42], secondStage_carry[41], secondStage_carry[40], 
      secondStage_carry[39], secondStage_carry[38], secondStage_carry[37], 
      secondStage_carry[36], secondStage_carry[35], secondStage_carry[34], 
      secondStage_carry[33], secondStage_carry[32], secondStage_carry[31], 
      secondStage_carry[30], secondStage_carry[29], secondStage_carry[28], 
      secondStage_carry[27], secondStage_carry[26], secondStage_carry[25], 
      secondStage_carry[24], secondStage_carry[23], secondStage_carry[22], 
      secondStage_carry[21], secondStage_carry[20], secondStage_carry[19], 
      secondStage_carry[18], secondStage_carry[17], secondStage_carry[16], 
      secondStage_carry[15], secondStage_carry[14], secondStage_carry[13], 
      secondStage_carry[12], secondStage_carry[11], secondStage_carry[10], 
      secondStage_carry[9], uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, 
      uc_48, uc_49}), .normalizedWires({uc_50, uc_51, 1'b0, uc_52, uc_53, uc_54, 
      uc_55, uc_56, uc_57, uc_58, uc_59, uc_60, uc_61, uc_62, uc_63, uc_64, 
      uc_65, uc_66, uc_67, uc_68, uc_69, uc_70, uc_71, uc_72, uc_73, uc_74, 
      uc_75, uc_76, uc_77, uc_78, uc_79, uc_80, uc_81, uc_82, uc_83, uc_84, 
      uc_85, uc_86, uc_87, uc_88, uc_89, uc_90, uc_91, uc_92, uc_93, uc_94, 
      uc_95, uc_96, uc_97, uc_98, uc_99, uc_100, uc_101, uc_102, uc_103, uc_104, 
      uc_105, uc_106, uc_107, uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, 
      uc_114, uc_115, uc_116, uc_117, uc_118, uc_119, uc_120, uc_121, uc_122, 
      uc_123, uc_124, uc_125, uc_126, uc_127, uc_128, uc_129, uc_130, uc_131, 
      uc_132, uc_133, uc_134, uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, 
      uc_141, uc_142, uc_143, uc_144, uc_145, uc_146, uc_147, uc_148, uc_149, 
      uc_150, uc_151, uc_152, uc_153, uc_154, uc_155, uc_156, uc_157, uc_158, 
      uc_159, uc_160, uc_161, uc_162, uc_163, uc_164, uc_165, uc_166, uc_167, 
      uc_168, uc_169, uc_170, uc_171, uc_172, uc_173, uc_174, uc_175, uc_176, 
      uc_177, uc_178, uc_179, uc_180, uc_181, uc_182, uc_183, uc_184, uc_185, 
      uc_186, uc_187, uc_188, uc_189, uc_190, uc_191, uc_192, uc_193, uc_194, 
      uc_195, uc_196, uc_197, uc_198, uc_199, uc_200, uc_201, uc_202, uc_203, 
      uc_204, uc_205, uc_206, uc_207, uc_208, uc_209, uc_210, uc_211, uc_212, 
      uc_213, uc_214, uc_215, uc_216, uc_217, uc_218, uc_219, uc_220, uc_221, 
      uc_222, uc_223, uc_224, uc_225, uc_226, uc_227, uc_228, uc_229, uc_230, 
      uc_231, uc_232, uc_233, uc_234, uc_235, uc_236, uc_237, uc_238, uc_239, 
      uc_240, uc_241, uc_242, uc_243, uc_244, uc_245, uc_246, uc_247, uc_248, 
      uc_249, uc_250, uc_251, uc_252, uc_253, uc_254, uc_255, uc_256, uc_257, 
      uc_258, uc_259, uc_260, uc_261, uc_262, uc_263, uc_264, uc_265, uc_266, 
      uc_267, uc_268, uc_269, uc_270, uc_271, uc_272, uc_273, uc_274, uc_275, 
      uc_276, uc_277, uc_278, uc_279, uc_280, uc_281, uc_282, uc_283, uc_284, 
      uc_285, uc_286, uc_287, uc_288, uc_289, uc_290, uc_291, uc_292, uc_293, 
      uc_294, uc_295, uc_296, uc_297, uc_298, uc_299, uc_300, uc_301, uc_302, 
      uc_303, uc_304, uc_305, uc_306, uc_307, uc_308, uc_309, uc_310, uc_311, 
      uc_312, uc_313, uc_314, uc_315, uc_316, uc_317, uc_318, uc_319, uc_320, 
      uc_321, uc_322, uc_323, uc_324, uc_325, uc_326, uc_327, uc_328, uc_329, 
      uc_330, uc_331, uc_332, uc_333, uc_334, uc_335, uc_336, uc_337, uc_338, 
      uc_339, uc_340, uc_341, uc_342, uc_343, uc_344, uc_345, uc_346, uc_347, 
      uc_348, uc_349, uc_350, uc_351, uc_352, uc_353, uc_354, uc_355, uc_356, 
      uc_357, uc_358, uc_359, uc_360, uc_361, uc_362, uc_363, uc_364, uc_365, 
      uc_366, uc_367, uc_368, uc_369, uc_370, uc_371, uc_372, uc_373, uc_374, 
      uc_375, uc_376, uc_377, uc_378, uc_379, uc_380, uc_381, uc_382, uc_383, 
      uc_384, uc_385, uc_386, uc_387, uc_388, uc_389, uc_390, uc_391, uc_392, 
      uc_393, uc_394, uc_395, uc_396, uc_397, uc_398, uc_399, uc_400, uc_401, 
      uc_402, uc_403, uc_404, uc_405, uc_406, uc_407, uc_408, uc_409, uc_410, 
      uc_411, uc_412, uc_413, uc_414, uc_415, uc_416, uc_417, uc_418, uc_419, 
      uc_420, uc_421, uc_422, uc_423, uc_424, uc_425, uc_426, uc_427, uc_428, 
      uc_429, uc_430, uc_431, uc_432, uc_433, uc_434, uc_435, uc_436, uc_437, 
      uc_438, uc_439, uc_440, uc_441, uc_442, uc_443, uc_444, uc_445, uc_446, 
      uc_447, uc_448, uc_449, uc_450, uc_451, uc_452, uc_453, uc_454, uc_455, 
      uc_456, uc_457, uc_458, uc_459, uc_460, uc_461, uc_462, uc_463, uc_464, 
      uc_465, uc_466, uc_467, uc_468, uc_469, uc_470, uc_471, uc_472, uc_473, 
      uc_474, uc_475, uc_476, uc_477, uc_478, uc_479, uc_480, uc_481, uc_482, 
      uc_483, uc_484, uc_485, uc_486, uc_487, uc_488, uc_489, uc_490, uc_491, 
      uc_492, uc_493, uc_494, uc_495, uc_496, uc_497, uc_498, uc_499, uc_500, 
      uc_501, uc_502, uc_503, uc_504, uc_505, uc_506, uc_507, uc_508, uc_509, 
      uc_510, uc_511, uc_512, uc_513, uc_514, uc_515, uc_516, uc_517, uc_518, 
      uc_519, uc_520, uc_521, uc_522, uc_523, uc_524, uc_525, uc_526, uc_527, 
      uc_528, uc_529, uc_530, uc_531, uc_532, uc_533, uc_534, uc_535, uc_536, 
      uc_537, uc_538, uc_539, uc_540, uc_541, uc_542, uc_543, uc_544, uc_545, 
      uc_546, uc_547, uc_548, uc_549, uc_550, uc_551, uc_552, uc_553, uc_554, 
      uc_555, uc_556, uc_557, uc_558, uc_559, uc_560, uc_561, uc_562, uc_563, 
      uc_564, uc_565, uc_566, uc_567, uc_568, uc_569, uc_570, 1'b0, uc_571, 
      uc_572, uc_573, uc_574, uc_575, uc_576, normalizedWires[1518], 
      normalizedWires[1517], normalizedWires[1516], normalizedWires[1515], 
      normalizedWires[1514], normalizedWires[1513], normalizedWires[1512], 
      normalizedWires[1511], normalizedWires[1510], normalizedWires[1509], 
      normalizedWires[1508], normalizedWires[1507], normalizedWires[1506], 
      normalizedWires[1505], normalizedWires[1504], normalizedWires[1503], 
      normalizedWires[1502], normalizedWires[1501], normalizedWires[1500], 
      normalizedWires[1499], normalizedWires[1498], normalizedWires[1497], 
      normalizedWires[1496], normalizedWires[1495], uc_577, uc_578, uc_579, 
      uc_580, uc_581, uc_582, uc_583, uc_584, uc_585, uc_586, uc_587, uc_588, 
      uc_589, uc_590, uc_591, uc_592, uc_593, uc_594, uc_595, uc_596, uc_597, 
      uc_598, uc_599, uc_600, uc_601, uc_602, uc_603, uc_604, uc_605, uc_606, 
      uc_607, uc_608, uc_609, uc_610, uc_611, uc_612, uc_613, uc_614, uc_615, 
      uc_616, uc_617, normalizedWires[1453], normalizedWires[1452], 
      normalizedWires[1451], normalizedWires[1450], normalizedWires[1449], 
      normalizedWires[1448], normalizedWires[1447], normalizedWires[1446], 
      normalizedWires[1445], normalizedWires[1444], normalizedWires[1443], 
      normalizedWires[1442], normalizedWires[1441], normalizedWires[1440], 
      normalizedWires[1439], normalizedWires[1438], normalizedWires[1437], 
      normalizedWires[1436], normalizedWires[1435], normalizedWires[1434], 
      normalizedWires[1433], normalizedWires[1432], normalizedWires[1431], 
      normalizedWires[1430], uc_618, uc_619, uc_620, uc_621, uc_622, uc_623, 
      uc_624, uc_625, uc_626, uc_627, uc_628, uc_629, uc_630, uc_631, uc_632, 
      uc_633, uc_634, uc_635, uc_636, uc_637, uc_638, uc_639, uc_640, uc_641, 
      uc_642, uc_643, uc_644, uc_645, uc_646, uc_647, uc_648, uc_649, uc_650, 
      uc_651, uc_652, uc_653, uc_654, uc_655, uc_656, uc_657, uc_658, 
      normalizedWires[1388], normalizedWires[1387], normalizedWires[1386], 
      normalizedWires[1385], normalizedWires[1384], normalizedWires[1383], 
      normalizedWires[1382], normalizedWires[1381], normalizedWires[1380], 
      normalizedWires[1379], normalizedWires[1378], normalizedWires[1377], 
      normalizedWires[1376], normalizedWires[1375], normalizedWires[1374], 
      normalizedWires[1373], normalizedWires[1372], normalizedWires[1371], 
      normalizedWires[1370], normalizedWires[1369], normalizedWires[1368], 
      normalizedWires[1367], normalizedWires[1366], normalizedWires[1365], 
      uc_659, uc_660, uc_661, uc_662, uc_663, uc_664, uc_665, uc_666, uc_667, 
      uc_668, uc_669, uc_670, uc_671, uc_672, uc_673, uc_674, uc_675, uc_676, 
      uc_677, uc_678, uc_679, uc_680, uc_681, uc_682, uc_683, uc_684, uc_685, 
      uc_686, uc_687, uc_688, uc_689, uc_690, uc_691, uc_692, uc_693, uc_694, 
      uc_695, uc_696, uc_697, uc_698, uc_699, normalizedWires[1323], 
      normalizedWires[1322], normalizedWires[1321], normalizedWires[1320], 
      normalizedWires[1319], normalizedWires[1318], normalizedWires[1317], 
      normalizedWires[1316], normalizedWires[1315], normalizedWires[1314], 
      normalizedWires[1313], normalizedWires[1312], normalizedWires[1311], 
      normalizedWires[1310], normalizedWires[1309], normalizedWires[1308], 
      normalizedWires[1307], normalizedWires[1306], normalizedWires[1305], 
      normalizedWires[1304], normalizedWires[1303], normalizedWires[1302], 
      normalizedWires[1301], normalizedWires[1300], uc_700, uc_701, uc_702, 
      uc_703, uc_704, uc_705, uc_706, uc_707, uc_708, uc_709, uc_710, uc_711, 
      uc_712, uc_713, uc_714, uc_715, uc_716, uc_717, uc_718, uc_719, uc_720, 
      uc_721, uc_722, uc_723, uc_724, uc_725, uc_726, uc_727, uc_728, uc_729, 
      uc_730, uc_731, uc_732, uc_733, uc_734, uc_735, uc_736, uc_737, uc_738, 
      uc_739, uc_740, normalizedWires[1258], normalizedWires[1257], 
      normalizedWires[1256], normalizedWires[1255], normalizedWires[1254], 
      normalizedWires[1253], normalizedWires[1252], normalizedWires[1251], 
      normalizedWires[1250], normalizedWires[1249], normalizedWires[1248], 
      normalizedWires[1247], normalizedWires[1246], normalizedWires[1245], 
      normalizedWires[1244], normalizedWires[1243], normalizedWires[1242], 
      normalizedWires[1241], normalizedWires[1240], normalizedWires[1239], 
      normalizedWires[1238], normalizedWires[1237], normalizedWires[1236], 
      normalizedWires[1235], uc_741, uc_742, uc_743, uc_744, uc_745, uc_746, 
      uc_747, uc_748, uc_749, uc_750, uc_751, uc_752, uc_753, uc_754, uc_755, 
      uc_756, uc_757, uc_758, uc_759, uc_760, uc_761, uc_762, uc_763, uc_764, 
      uc_765, uc_766, uc_767, uc_768, uc_769, uc_770, uc_771, uc_772, uc_773, 
      uc_774, uc_775, uc_776, uc_777, uc_778, uc_779, uc_780, uc_781, 
      normalizedWires[1193], normalizedWires[1192], normalizedWires[1191], 
      normalizedWires[1190], normalizedWires[1189], normalizedWires[1188], 
      normalizedWires[1187], normalizedWires[1186], normalizedWires[1185], 
      normalizedWires[1184], normalizedWires[1183], normalizedWires[1182], 
      normalizedWires[1181], normalizedWires[1180], normalizedWires[1179], 
      normalizedWires[1178], normalizedWires[1177], normalizedWires[1176], 
      normalizedWires[1175], normalizedWires[1174], normalizedWires[1173], 
      normalizedWires[1172], normalizedWires[1171], normalizedWires[1170], 
      uc_782, uc_783, uc_784, uc_785, uc_786, uc_787, uc_788, uc_789, uc_790, 
      uc_791, uc_792, uc_793, uc_794, uc_795, uc_796, uc_797, uc_798, uc_799, 
      uc_800, uc_801, uc_802, uc_803, uc_804, uc_805, uc_806, uc_807, uc_808, 
      uc_809, uc_810, uc_811, uc_812, uc_813, uc_814, uc_815, uc_816, uc_817, 
      uc_818, uc_819, uc_820, uc_821, uc_822, normalizedWires[1128], 
      normalizedWires[1127], normalizedWires[1126], normalizedWires[1125], 
      normalizedWires[1124], normalizedWires[1123], normalizedWires[1122], 
      normalizedWires[1121], normalizedWires[1120], normalizedWires[1119], 
      normalizedWires[1118], normalizedWires[1117], normalizedWires[1116], 
      normalizedWires[1115], normalizedWires[1114], normalizedWires[1113], 
      normalizedWires[1112], normalizedWires[1111], normalizedWires[1110], 
      normalizedWires[1109], normalizedWires[1108], normalizedWires[1107], 
      normalizedWires[1106], normalizedWires[1105], uc_823, uc_824, uc_825, 
      uc_826, uc_827, uc_828, uc_829, uc_830, uc_831, uc_832, uc_833, uc_834, 
      uc_835, uc_836, uc_837, uc_838, uc_839, uc_840, uc_841, uc_842, uc_843, 
      uc_844, uc_845, uc_846, uc_847, uc_848, uc_849, uc_850, uc_851, uc_852, 
      uc_853, uc_854, uc_855, uc_856, uc_857, uc_858, uc_859, uc_860, uc_861, 
      uc_862, uc_863, normalizedWires[1063], normalizedWires[1062], 
      normalizedWires[1061], normalizedWires[1060], normalizedWires[1059], 
      normalizedWires[1058], normalizedWires[1057], normalizedWires[1056], 
      normalizedWires[1055], normalizedWires[1054], normalizedWires[1053], 
      normalizedWires[1052], normalizedWires[1051], normalizedWires[1050], 
      normalizedWires[1049], normalizedWires[1048], normalizedWires[1047], 
      normalizedWires[1046], normalizedWires[1045], normalizedWires[1044], 
      normalizedWires[1043], normalizedWires[1042], normalizedWires[1041], 
      normalizedWires[1040], uc_864, uc_865, uc_866, uc_867, uc_868, uc_869, 
      uc_870, uc_871, uc_872, uc_873, uc_874, uc_875, uc_876, uc_877, uc_878, 
      uc_879, uc_880, uc_881, uc_882, uc_883, uc_884, uc_885, uc_886, uc_887, 
      uc_888, uc_889, uc_890, uc_891, uc_892, uc_893, uc_894, uc_895, uc_896, 
      uc_897, uc_898, uc_899, uc_900, uc_901, uc_902, uc_903, uc_904, 
      normalizedWires[998], normalizedWires[997], normalizedWires[996], 
      normalizedWires[995], normalizedWires[994], normalizedWires[993], 
      normalizedWires[992], normalizedWires[991], normalizedWires[990], 
      normalizedWires[989], normalizedWires[988], normalizedWires[987], 
      normalizedWires[986], normalizedWires[985], normalizedWires[984], 
      normalizedWires[983], normalizedWires[982], normalizedWires[981], 
      normalizedWires[980], normalizedWires[979], normalizedWires[978], 
      normalizedWires[977], normalizedWires[976], normalizedWires[975], uc_905, 
      uc_906, uc_907, uc_908, uc_909, uc_910, uc_911, uc_912, uc_913, uc_914, 
      uc_915, uc_916, uc_917, uc_918, uc_919, uc_920, uc_921, uc_922, uc_923, 
      uc_924, uc_925, uc_926, uc_927, uc_928, uc_929, uc_930, uc_931, uc_932, 
      uc_933, uc_934, uc_935, uc_936, uc_937, uc_938, uc_939, uc_940, uc_941, 
      uc_942, uc_943, uc_944, uc_945, normalizedWires[933], normalizedWires[932], 
      normalizedWires[931], normalizedWires[930], normalizedWires[929], 
      normalizedWires[928], normalizedWires[927], normalizedWires[926], 
      normalizedWires[925], normalizedWires[924], normalizedWires[923], 
      normalizedWires[922], normalizedWires[921], normalizedWires[920], 
      normalizedWires[919], normalizedWires[918], normalizedWires[917], 
      normalizedWires[916], normalizedWires[915], normalizedWires[914], 
      normalizedWires[913], normalizedWires[912], normalizedWires[911], 
      normalizedWires[910], uc_946, uc_947, uc_948, uc_949, uc_950, uc_951, 
      uc_952, uc_953, uc_954, uc_955, uc_956, uc_957, uc_958, uc_959, uc_960, 
      uc_961, uc_962, uc_963, uc_964, uc_965, uc_966, uc_967, uc_968, uc_969, 
      uc_970, uc_971, uc_972, uc_973, uc_974, uc_975, uc_976, uc_977, uc_978, 
      uc_979, uc_980, uc_981, uc_982, uc_983, uc_984, uc_985, uc_986, 
      normalizedWires[868], normalizedWires[867], normalizedWires[866], 
      normalizedWires[865], normalizedWires[864], normalizedWires[863], 
      normalizedWires[862], normalizedWires[861], normalizedWires[860], 
      normalizedWires[859], normalizedWires[858], normalizedWires[857], 
      normalizedWires[856], normalizedWires[855], normalizedWires[854], 
      normalizedWires[853], normalizedWires[852], normalizedWires[851], 
      normalizedWires[850], normalizedWires[849], normalizedWires[848], 
      normalizedWires[847], normalizedWires[846], normalizedWires[845], uc_987, 
      uc_988, uc_989, uc_990, uc_991, uc_992, uc_993, uc_994, uc_995, uc_996, 
      uc_997, uc_998, uc_999, uc_1000, uc_1001, uc_1002, uc_1003, uc_1004, 
      uc_1005, uc_1006, uc_1007, uc_1008, uc_1009, uc_1010, uc_1011, uc_1012, 
      uc_1013, uc_1014, uc_1015, uc_1016, uc_1017, uc_1018, uc_1019, uc_1020, 
      uc_1021, uc_1022, uc_1023, uc_1024, uc_1025, uc_1026, uc_1027, 
      normalizedWires[803], normalizedWires[802], normalizedWires[801], 
      normalizedWires[800], normalizedWires[799], normalizedWires[798], 
      normalizedWires[797], normalizedWires[796], normalizedWires[795], 
      normalizedWires[794], normalizedWires[793], normalizedWires[792], 
      normalizedWires[791], normalizedWires[790], normalizedWires[789], 
      normalizedWires[788], normalizedWires[787], normalizedWires[786], 
      normalizedWires[785], normalizedWires[784], normalizedWires[783], 
      normalizedWires[782], normalizedWires[781], normalizedWires[780], uc_1028, 
      uc_1029, uc_1030, uc_1031, uc_1032, uc_1033, uc_1034, uc_1035, uc_1036, 
      uc_1037, uc_1038, uc_1039, uc_1040, uc_1041, uc_1042, uc_1043, uc_1044, 
      uc_1045, uc_1046, uc_1047, uc_1048, uc_1049, uc_1050, uc_1051, uc_1052, 
      uc_1053, uc_1054, uc_1055, uc_1056, uc_1057, uc_1058, uc_1059, uc_1060, 
      uc_1061, uc_1062, uc_1063, uc_1064, uc_1065, uc_1066, uc_1067, uc_1068, 
      normalizedWires[738], normalizedWires[737], normalizedWires[736], 
      normalizedWires[735], normalizedWires[734], normalizedWires[733], 
      normalizedWires[732], normalizedWires[731], normalizedWires[730], 
      normalizedWires[729], normalizedWires[728], normalizedWires[727], 
      normalizedWires[726], normalizedWires[725], normalizedWires[724], 
      normalizedWires[723], normalizedWires[722], normalizedWires[721], 
      normalizedWires[720], normalizedWires[719], normalizedWires[718], 
      normalizedWires[717], normalizedWires[716], normalizedWires[715], uc_1069, 
      uc_1070, uc_1071, uc_1072, uc_1073, uc_1074, uc_1075, uc_1076, uc_1077, 
      uc_1078, uc_1079, uc_1080, uc_1081, uc_1082, uc_1083, uc_1084, uc_1085, 
      uc_1086, uc_1087, uc_1088, uc_1089, uc_1090, uc_1091, uc_1092, uc_1093, 
      uc_1094, uc_1095, uc_1096, uc_1097, uc_1098, uc_1099, uc_1100, uc_1101, 
      uc_1102, uc_1103, uc_1104, uc_1105, uc_1106, uc_1107, uc_1108, uc_1109, 
      normalizedWires[673], normalizedWires[672], normalizedWires[671], 
      normalizedWires[670], normalizedWires[669], normalizedWires[668], 
      normalizedWires[667], normalizedWires[666], normalizedWires[665], 
      normalizedWires[664], normalizedWires[663], normalizedWires[662], 
      normalizedWires[661], normalizedWires[660], normalizedWires[659], 
      normalizedWires[658], normalizedWires[657], normalizedWires[656], 
      normalizedWires[655], normalizedWires[654], normalizedWires[653], 
      normalizedWires[652], normalizedWires[651], normalizedWires[650], uc_1110, 
      uc_1111, uc_1112, uc_1113, uc_1114, uc_1115, uc_1116, uc_1117, uc_1118, 
      uc_1119, uc_1120, uc_1121, uc_1122, uc_1123, uc_1124, uc_1125, uc_1126, 
      uc_1127, uc_1128, uc_1129, uc_1130, uc_1131, uc_1132, uc_1133, uc_1134, 
      uc_1135, uc_1136, uc_1137, uc_1138, uc_1139, uc_1140, uc_1141, uc_1142, 
      uc_1143, uc_1144, uc_1145, uc_1146, uc_1147, uc_1148, uc_1149, uc_1150, 
      normalizedWires[608], normalizedWires[607], normalizedWires[606], 
      normalizedWires[605], normalizedWires[604], normalizedWires[603], 
      normalizedWires[602], normalizedWires[601], normalizedWires[600], 
      normalizedWires[599], normalizedWires[598], normalizedWires[597], 
      normalizedWires[596], normalizedWires[595], normalizedWires[594], 
      normalizedWires[593], normalizedWires[592], normalizedWires[591], 
      normalizedWires[590], normalizedWires[589], normalizedWires[588], 
      normalizedWires[587], normalizedWires[586], normalizedWires[585], uc_1151, 
      uc_1152, uc_1153, uc_1154, uc_1155, uc_1156, uc_1157, uc_1158, uc_1159, 
      uc_1160, uc_1161, uc_1162, uc_1163, uc_1164, uc_1165, uc_1166, uc_1167, 
      uc_1168, uc_1169, uc_1170, uc_1171, uc_1172, uc_1173, uc_1174, uc_1175, 
      uc_1176, uc_1177, uc_1178, uc_1179, uc_1180, uc_1181, uc_1182, uc_1183, 
      uc_1184, uc_1185, uc_1186, uc_1187, uc_1188, uc_1189, uc_1190, uc_1191, 
      normalizedWires[543], normalizedWires[542], normalizedWires[541], 
      normalizedWires[540], normalizedWires[539], normalizedWires[538], 
      normalizedWires[537], normalizedWires[536], normalizedWires[535], 
      normalizedWires[534], normalizedWires[533], normalizedWires[532], 
      normalizedWires[531], normalizedWires[530], normalizedWires[529], 
      normalizedWires[528], normalizedWires[527], normalizedWires[526], 
      normalizedWires[525], normalizedWires[524], normalizedWires[523], 
      normalizedWires[522], normalizedWires[521], normalizedWires[520], uc_1192, 
      uc_1193, uc_1194, uc_1195, uc_1196, uc_1197, uc_1198, uc_1199, uc_1200, 
      uc_1201, uc_1202, uc_1203, uc_1204, uc_1205, uc_1206, uc_1207, uc_1208, 
      uc_1209, uc_1210, uc_1211, uc_1212, uc_1213, uc_1214, uc_1215, uc_1216, 
      uc_1217, uc_1218, uc_1219, uc_1220, uc_1221, uc_1222, uc_1223, uc_1224, 
      uc_1225, uc_1226, uc_1227, uc_1228, uc_1229, uc_1230, uc_1231, uc_1232, 
      normalizedWires[478], normalizedWires[477], normalizedWires[476], 
      normalizedWires[475], normalizedWires[474], normalizedWires[473], 
      normalizedWires[472], normalizedWires[471], normalizedWires[470], 
      normalizedWires[469], normalizedWires[468], normalizedWires[467], 
      normalizedWires[466], normalizedWires[465], normalizedWires[464], 
      normalizedWires[463], normalizedWires[462], normalizedWires[461], 
      normalizedWires[460], normalizedWires[459], normalizedWires[458], 
      normalizedWires[457], normalizedWires[456], normalizedWires[455], uc_1233, 
      uc_1234, uc_1235, uc_1236, uc_1237, uc_1238, uc_1239, uc_1240, uc_1241, 
      uc_1242, uc_1243, uc_1244, uc_1245, uc_1246, uc_1247, uc_1248, uc_1249, 
      uc_1250, uc_1251, uc_1252, uc_1253, uc_1254, uc_1255, uc_1256, uc_1257, 
      uc_1258, uc_1259, uc_1260, uc_1261, uc_1262, uc_1263, uc_1264, uc_1265, 
      uc_1266, uc_1267, uc_1268, uc_1269, uc_1270, uc_1271, uc_1272, uc_1273, 
      normalizedWires[413], normalizedWires[412], normalizedWires[411], 
      normalizedWires[410], normalizedWires[409], normalizedWires[408], 
      normalizedWires[407], normalizedWires[406], normalizedWires[405], 
      normalizedWires[404], normalizedWires[403], normalizedWires[402], 
      normalizedWires[401], normalizedWires[400], normalizedWires[399], 
      normalizedWires[398], normalizedWires[397], normalizedWires[396], 
      normalizedWires[395], normalizedWires[394], normalizedWires[393], 
      normalizedWires[392], normalizedWires[391], normalizedWires[390], uc_1274, 
      uc_1275, uc_1276, uc_1277, uc_1278, uc_1279, uc_1280, uc_1281, uc_1282, 
      uc_1283, uc_1284, uc_1285, uc_1286, uc_1287, uc_1288, uc_1289, uc_1290, 
      uc_1291, uc_1292, uc_1293, uc_1294, uc_1295, uc_1296, uc_1297, uc_1298, 
      uc_1299, uc_1300, uc_1301, uc_1302, uc_1303, uc_1304, uc_1305, uc_1306, 
      uc_1307, uc_1308, uc_1309, uc_1310, uc_1311, uc_1312, uc_1313, uc_1314, 
      normalizedWires[348], normalizedWires[347], normalizedWires[346], 
      normalizedWires[345], normalizedWires[344], normalizedWires[343], 
      normalizedWires[342], normalizedWires[341], normalizedWires[340], 
      normalizedWires[339], normalizedWires[338], normalizedWires[337], 
      normalizedWires[336], normalizedWires[335], normalizedWires[334], 
      normalizedWires[333], normalizedWires[332], normalizedWires[331], 
      normalizedWires[330], normalizedWires[329], normalizedWires[328], 
      normalizedWires[327], normalizedWires[326], normalizedWires[325], uc_1315, 
      uc_1316, uc_1317, uc_1318, uc_1319, uc_1320, uc_1321, uc_1322, uc_1323, 
      uc_1324, uc_1325, uc_1326, uc_1327, uc_1328, uc_1329, uc_1330, uc_1331, 
      uc_1332, uc_1333, uc_1334, uc_1335, uc_1336, uc_1337, uc_1338, uc_1339, 
      uc_1340, uc_1341, uc_1342, uc_1343, uc_1344, uc_1345, uc_1346, uc_1347, 
      uc_1348, uc_1349, uc_1350, uc_1351, uc_1352, uc_1353, uc_1354, uc_1355, 
      normalizedWires[283], normalizedWires[282], normalizedWires[281], 
      normalizedWires[280], normalizedWires[279], normalizedWires[278], 
      normalizedWires[277], normalizedWires[276], normalizedWires[275], 
      normalizedWires[274], normalizedWires[273], normalizedWires[272], 
      normalizedWires[271], normalizedWires[270], normalizedWires[269], 
      normalizedWires[268], normalizedWires[267], normalizedWires[266], 
      normalizedWires[265], normalizedWires[264], normalizedWires[263], 
      normalizedWires[262], normalizedWires[261], normalizedWires[260], uc_1356, 
      uc_1357, uc_1358, uc_1359, uc_1360, uc_1361, uc_1362, uc_1363, uc_1364, 
      uc_1365, uc_1366, uc_1367, uc_1368, uc_1369, uc_1370, uc_1371, uc_1372, 
      uc_1373, uc_1374, uc_1375, uc_1376, uc_1377, uc_1378, uc_1379, uc_1380, 
      uc_1381, uc_1382, uc_1383, uc_1384, uc_1385, uc_1386, uc_1387, uc_1388, 
      uc_1389, uc_1390, uc_1391, uc_1392, uc_1393, uc_1394, uc_1395, uc_1396, 
      normalizedWires[218], normalizedWires[217], normalizedWires[216], 
      normalizedWires[215], normalizedWires[214], normalizedWires[213], 
      normalizedWires[212], normalizedWires[211], normalizedWires[210], 
      normalizedWires[209], normalizedWires[208], normalizedWires[207], 
      normalizedWires[206], normalizedWires[205], normalizedWires[204], 
      normalizedWires[203], normalizedWires[202], normalizedWires[201], 
      normalizedWires[200], normalizedWires[199], normalizedWires[198], 
      normalizedWires[197], normalizedWires[196], normalizedWires[195], uc_1397, 
      uc_1398, uc_1399, uc_1400, uc_1401, uc_1402, uc_1403, uc_1404, uc_1405, 
      uc_1406, uc_1407, uc_1408, uc_1409, uc_1410, uc_1411, uc_1412, uc_1413, 
      uc_1414, uc_1415, uc_1416, uc_1417, uc_1418, uc_1419, uc_1420, uc_1421, 
      uc_1422, uc_1423, uc_1424, uc_1425, uc_1426, uc_1427, uc_1428, uc_1429, 
      uc_1430, uc_1431, uc_1432, uc_1433, uc_1434, uc_1435, uc_1436, uc_1437, 
      normalizedWires[153], normalizedWires[152], normalizedWires[151], 
      normalizedWires[150], normalizedWires[149], normalizedWires[148], 
      normalizedWires[147], normalizedWires[146], normalizedWires[145], 
      normalizedWires[144], normalizedWires[143], normalizedWires[142], 
      normalizedWires[141], normalizedWires[140], normalizedWires[139], 
      normalizedWires[138], normalizedWires[137], normalizedWires[136], 
      normalizedWires[135], normalizedWires[134], normalizedWires[133], 
      normalizedWires[132], normalizedWires[131], normalizedWires[130], uc_1438, 
      uc_1439, uc_1440, uc_1441, uc_1442, uc_1443, uc_1444, uc_1445, uc_1446, 
      uc_1447, uc_1448, uc_1449, uc_1450, uc_1451, uc_1452, uc_1453, uc_1454, 
      uc_1455, uc_1456, uc_1457, uc_1458, uc_1459, uc_1460, uc_1461, uc_1462, 
      uc_1463, uc_1464, uc_1465, uc_1466, uc_1467, uc_1468, uc_1469, uc_1470, 
      uc_1471, uc_1472, uc_1473, uc_1474, uc_1475, uc_1476, uc_1477, uc_1478, 
      normalizedWires[88], normalizedWires[87], normalizedWires[86], 
      normalizedWires[85], normalizedWires[84], normalizedWires[83], 
      normalizedWires[82], normalizedWires[81], normalizedWires[80], 
      normalizedWires[79], normalizedWires[78], normalizedWires[77], 
      normalizedWires[76], normalizedWires[75], normalizedWires[74], 
      normalizedWires[73], normalizedWires[72], normalizedWires[71], 
      normalizedWires[70], normalizedWires[69], normalizedWires[68], 
      normalizedWires[67], normalizedWires[66], normalizedWires[65], uc_1479, 
      uc_1480, uc_1481, uc_1482, uc_1483, uc_1484, uc_1485, uc_1486, uc_1487, 
      uc_1488, uc_1489, uc_1490, uc_1491, uc_1492, uc_1493, uc_1494, uc_1495, 
      uc_1496, uc_1497, uc_1498, uc_1499, uc_1500, uc_1501, uc_1502, uc_1503, 
      uc_1504, uc_1505, uc_1506, uc_1507, uc_1508, uc_1509, uc_1510, uc_1511, 
      uc_1512, uc_1513, uc_1514, uc_1515, uc_1516, uc_1517, uc_1518, uc_1519, 
      normalizedWires[23], normalizedWires[22], normalizedWires[21], 
      normalizedWires[20], normalizedWires[19], normalizedWires[18], 
      normalizedWires[17], normalizedWires[16], normalizedWires[15], 
      normalizedWires[14], normalizedWires[13], normalizedWires[12], 
      normalizedWires[11], normalizedWires[10], normalizedWires[9], 
      normalizedWires[8], normalizedWires[7], normalizedWires[6], 
      normalizedWires[5], normalizedWires[4], normalizedWires[3], 
      normalizedWires[2], normalizedWires[1], uc_1520}));
   multiplyAllBits firstStage (.normalizedWires({uc_1521, uc_1522, uc_1523, 
      uc_1524, uc_1525, uc_1526, uc_1527, uc_1528, uc_1529, uc_1530, uc_1531, 
      uc_1532, uc_1533, uc_1534, uc_1535, uc_1536, uc_1537, uc_1538, uc_1539, 
      uc_1540, uc_1541, uc_1542, uc_1543, uc_1544, uc_1545, uc_1546, uc_1547, 
      uc_1548, uc_1549, uc_1550, uc_1551, uc_1552, uc_1553, uc_1554, uc_1555, 
      uc_1556, uc_1557, uc_1558, uc_1559, uc_1560, uc_1561, uc_1562, uc_1563, 
      uc_1564, uc_1565, uc_1566, uc_1567, uc_1568, uc_1569, uc_1570, uc_1571, 
      uc_1572, uc_1573, uc_1574, uc_1575, uc_1576, uc_1577, uc_1578, uc_1579, 
      uc_1580, uc_1581, uc_1582, uc_1583, uc_1584, uc_1585, uc_1586, uc_1587, 
      uc_1588, uc_1589, uc_1590, uc_1591, uc_1592, uc_1593, uc_1594, uc_1595, 
      uc_1596, uc_1597, uc_1598, uc_1599, uc_1600, uc_1601, uc_1602, uc_1603, 
      uc_1604, uc_1605, uc_1606, uc_1607, uc_1608, uc_1609, uc_1610, uc_1611, 
      uc_1612, uc_1613, uc_1614, uc_1615, uc_1616, uc_1617, uc_1618, uc_1619, 
      uc_1620, uc_1621, uc_1622, uc_1623, uc_1624, uc_1625, uc_1626, uc_1627, 
      uc_1628, uc_1629, uc_1630, uc_1631, uc_1632, uc_1633, uc_1634, uc_1635, 
      uc_1636, uc_1637, uc_1638, uc_1639, uc_1640, uc_1641, uc_1642, uc_1643, 
      uc_1644, uc_1645, uc_1646, uc_1647, uc_1648, uc_1649, uc_1650, uc_1651, 
      uc_1652, uc_1653, uc_1654, uc_1655, uc_1656, uc_1657, uc_1658, uc_1659, 
      uc_1660, uc_1661, uc_1662, uc_1663, uc_1664, uc_1665, uc_1666, uc_1667, 
      uc_1668, uc_1669, uc_1670, uc_1671, uc_1672, uc_1673, uc_1674, uc_1675, 
      uc_1676, uc_1677, uc_1678, uc_1679, uc_1680, uc_1681, uc_1682, uc_1683, 
      uc_1684, uc_1685, uc_1686, uc_1687, uc_1688, uc_1689, uc_1690, uc_1691, 
      uc_1692, uc_1693, uc_1694, uc_1695, uc_1696, uc_1697, uc_1698, uc_1699, 
      uc_1700, uc_1701, uc_1702, uc_1703, uc_1704, uc_1705, uc_1706, uc_1707, 
      uc_1708, uc_1709, uc_1710, uc_1711, uc_1712, uc_1713, uc_1714, uc_1715, 
      uc_1716, uc_1717, uc_1718, uc_1719, uc_1720, uc_1721, uc_1722, uc_1723, 
      uc_1724, uc_1725, uc_1726, uc_1727, uc_1728, uc_1729, uc_1730, uc_1731, 
      uc_1732, uc_1733, uc_1734, uc_1735, uc_1736, uc_1737, uc_1738, uc_1739, 
      uc_1740, uc_1741, uc_1742, uc_1743, uc_1744, uc_1745, uc_1746, uc_1747, 
      uc_1748, uc_1749, uc_1750, uc_1751, uc_1752, uc_1753, uc_1754, uc_1755, 
      uc_1756, uc_1757, uc_1758, uc_1759, uc_1760, uc_1761, uc_1762, uc_1763, 
      uc_1764, uc_1765, uc_1766, uc_1767, uc_1768, uc_1769, uc_1770, uc_1771, 
      uc_1772, uc_1773, uc_1774, uc_1775, uc_1776, uc_1777, uc_1778, uc_1779, 
      uc_1780, uc_1781, uc_1782, uc_1783, uc_1784, uc_1785, uc_1786, uc_1787, 
      uc_1788, uc_1789, uc_1790, uc_1791, uc_1792, uc_1793, uc_1794, uc_1795, 
      uc_1796, uc_1797, uc_1798, uc_1799, uc_1800, uc_1801, uc_1802, uc_1803, 
      uc_1804, uc_1805, uc_1806, uc_1807, uc_1808, uc_1809, uc_1810, uc_1811, 
      uc_1812, uc_1813, uc_1814, uc_1815, uc_1816, uc_1817, uc_1818, uc_1819, 
      uc_1820, uc_1821, uc_1822, uc_1823, uc_1824, uc_1825, uc_1826, uc_1827, 
      uc_1828, uc_1829, uc_1830, uc_1831, uc_1832, uc_1833, uc_1834, uc_1835, 
      uc_1836, uc_1837, uc_1838, uc_1839, uc_1840, uc_1841, uc_1842, uc_1843, 
      uc_1844, uc_1845, uc_1846, uc_1847, uc_1848, uc_1849, uc_1850, uc_1851, 
      uc_1852, uc_1853, uc_1854, uc_1855, uc_1856, uc_1857, uc_1858, uc_1859, 
      uc_1860, uc_1861, uc_1862, uc_1863, uc_1864, uc_1865, uc_1866, uc_1867, 
      uc_1868, uc_1869, uc_1870, uc_1871, uc_1872, uc_1873, uc_1874, uc_1875, 
      uc_1876, uc_1877, uc_1878, uc_1879, uc_1880, uc_1881, uc_1882, uc_1883, 
      uc_1884, uc_1885, uc_1886, uc_1887, uc_1888, uc_1889, uc_1890, uc_1891, 
      uc_1892, uc_1893, uc_1894, uc_1895, uc_1896, uc_1897, uc_1898, uc_1899, 
      uc_1900, uc_1901, uc_1902, uc_1903, uc_1904, uc_1905, uc_1906, uc_1907, 
      uc_1908, uc_1909, uc_1910, uc_1911, uc_1912, uc_1913, uc_1914, uc_1915, 
      uc_1916, uc_1917, uc_1918, uc_1919, uc_1920, uc_1921, uc_1922, uc_1923, 
      uc_1924, uc_1925, uc_1926, uc_1927, uc_1928, uc_1929, uc_1930, uc_1931, 
      uc_1932, uc_1933, uc_1934, uc_1935, uc_1936, uc_1937, uc_1938, uc_1939, 
      uc_1940, uc_1941, uc_1942, uc_1943, uc_1944, uc_1945, uc_1946, uc_1947, 
      uc_1948, uc_1949, uc_1950, uc_1951, uc_1952, uc_1953, uc_1954, uc_1955, 
      uc_1956, uc_1957, uc_1958, uc_1959, uc_1960, uc_1961, uc_1962, uc_1963, 
      uc_1964, uc_1965, uc_1966, uc_1967, uc_1968, uc_1969, uc_1970, uc_1971, 
      uc_1972, uc_1973, uc_1974, uc_1975, uc_1976, uc_1977, uc_1978, uc_1979, 
      uc_1980, uc_1981, uc_1982, uc_1983, uc_1984, uc_1985, uc_1986, uc_1987, 
      uc_1988, uc_1989, uc_1990, uc_1991, uc_1992, uc_1993, uc_1994, uc_1995, 
      uc_1996, uc_1997, uc_1998, uc_1999, uc_2000, uc_2001, uc_2002, uc_2003, 
      uc_2004, uc_2005, uc_2006, uc_2007, uc_2008, uc_2009, uc_2010, uc_2011, 
      uc_2012, uc_2013, uc_2014, uc_2015, uc_2016, uc_2017, uc_2018, uc_2019, 
      uc_2020, uc_2021, uc_2022, uc_2023, uc_2024, uc_2025, uc_2026, uc_2027, 
      uc_2028, uc_2029, uc_2030, uc_2031, uc_2032, uc_2033, uc_2034, uc_2035, 
      uc_2036, uc_2037, uc_2038, uc_2039, uc_2040, uc_2041, uc_2042, uc_2043, 
      uc_2044, uc_2045, uc_2046, uc_2047, uc_2048, uc_2049, uc_2050, 
      normalizedWires[1517], normalizedWires[1516], normalizedWires[1515], 
      normalizedWires[1514], normalizedWires[1513], normalizedWires[1512], 
      normalizedWires[1511], normalizedWires[1510], normalizedWires[1509], 
      normalizedWires[1508], normalizedWires[1507], normalizedWires[1506], 
      normalizedWires[1505], normalizedWires[1504], normalizedWires[1503], 
      normalizedWires[1502], normalizedWires[1501], normalizedWires[1500], 
      normalizedWires[1499], normalizedWires[1498], normalizedWires[1497], 
      normalizedWires[1496], normalizedWires[1495], uc_2051, uc_2052, uc_2053, 
      uc_2054, uc_2055, uc_2056, uc_2057, uc_2058, uc_2059, uc_2060, uc_2061, 
      uc_2062, uc_2063, uc_2064, uc_2065, uc_2066, uc_2067, uc_2068, uc_2069, 
      uc_2070, uc_2071, uc_2072, uc_2073, uc_2074, uc_2075, uc_2076, uc_2077, 
      uc_2078, uc_2079, uc_2080, uc_2081, uc_2082, uc_2083, uc_2084, uc_2085, 
      uc_2086, uc_2087, uc_2088, uc_2089, uc_2090, uc_2091, 
      normalizedWires[1453], normalizedWires[1452], normalizedWires[1451], 
      normalizedWires[1450], normalizedWires[1449], normalizedWires[1448], 
      normalizedWires[1447], normalizedWires[1446], normalizedWires[1445], 
      normalizedWires[1444], normalizedWires[1443], normalizedWires[1442], 
      normalizedWires[1441], normalizedWires[1440], normalizedWires[1439], 
      normalizedWires[1438], normalizedWires[1437], normalizedWires[1436], 
      normalizedWires[1435], normalizedWires[1434], normalizedWires[1433], 
      normalizedWires[1432], normalizedWires[1431], normalizedWires[1430], 
      uc_2092, uc_2093, uc_2094, uc_2095, uc_2096, uc_2097, uc_2098, uc_2099, 
      uc_2100, uc_2101, uc_2102, uc_2103, uc_2104, uc_2105, uc_2106, uc_2107, 
      uc_2108, uc_2109, uc_2110, uc_2111, uc_2112, uc_2113, uc_2114, uc_2115, 
      uc_2116, uc_2117, uc_2118, uc_2119, uc_2120, uc_2121, uc_2122, uc_2123, 
      uc_2124, uc_2125, uc_2126, uc_2127, uc_2128, uc_2129, uc_2130, uc_2131, 
      uc_2132, normalizedWires[1388], normalizedWires[1387], 
      normalizedWires[1386], normalizedWires[1385], normalizedWires[1384], 
      normalizedWires[1383], normalizedWires[1382], normalizedWires[1381], 
      normalizedWires[1380], normalizedWires[1379], normalizedWires[1378], 
      normalizedWires[1377], normalizedWires[1376], normalizedWires[1375], 
      normalizedWires[1374], normalizedWires[1373], normalizedWires[1372], 
      normalizedWires[1371], normalizedWires[1370], normalizedWires[1369], 
      normalizedWires[1368], normalizedWires[1367], normalizedWires[1366], 
      normalizedWires[1365], uc_2133, uc_2134, uc_2135, uc_2136, uc_2137, 
      uc_2138, uc_2139, uc_2140, uc_2141, uc_2142, uc_2143, uc_2144, uc_2145, 
      uc_2146, uc_2147, uc_2148, uc_2149, uc_2150, uc_2151, uc_2152, uc_2153, 
      uc_2154, uc_2155, uc_2156, uc_2157, uc_2158, uc_2159, uc_2160, uc_2161, 
      uc_2162, uc_2163, uc_2164, uc_2165, uc_2166, uc_2167, uc_2168, uc_2169, 
      uc_2170, uc_2171, uc_2172, uc_2173, normalizedWires[1323], 
      normalizedWires[1322], normalizedWires[1321], normalizedWires[1320], 
      normalizedWires[1319], normalizedWires[1318], normalizedWires[1317], 
      normalizedWires[1316], normalizedWires[1315], normalizedWires[1314], 
      normalizedWires[1313], normalizedWires[1312], normalizedWires[1311], 
      normalizedWires[1310], normalizedWires[1309], normalizedWires[1308], 
      normalizedWires[1307], normalizedWires[1306], normalizedWires[1305], 
      normalizedWires[1304], normalizedWires[1303], normalizedWires[1302], 
      normalizedWires[1301], normalizedWires[1300], uc_2174, uc_2175, uc_2176, 
      uc_2177, uc_2178, uc_2179, uc_2180, uc_2181, uc_2182, uc_2183, uc_2184, 
      uc_2185, uc_2186, uc_2187, uc_2188, uc_2189, uc_2190, uc_2191, uc_2192, 
      uc_2193, uc_2194, uc_2195, uc_2196, uc_2197, uc_2198, uc_2199, uc_2200, 
      uc_2201, uc_2202, uc_2203, uc_2204, uc_2205, uc_2206, uc_2207, uc_2208, 
      uc_2209, uc_2210, uc_2211, uc_2212, uc_2213, uc_2214, 
      normalizedWires[1258], normalizedWires[1257], normalizedWires[1256], 
      normalizedWires[1255], normalizedWires[1254], normalizedWires[1253], 
      normalizedWires[1252], normalizedWires[1251], normalizedWires[1250], 
      normalizedWires[1249], normalizedWires[1248], normalizedWires[1247], 
      normalizedWires[1246], normalizedWires[1245], normalizedWires[1244], 
      normalizedWires[1243], normalizedWires[1242], normalizedWires[1241], 
      normalizedWires[1240], normalizedWires[1239], normalizedWires[1238], 
      normalizedWires[1237], normalizedWires[1236], normalizedWires[1235], 
      uc_2215, uc_2216, uc_2217, uc_2218, uc_2219, uc_2220, uc_2221, uc_2222, 
      uc_2223, uc_2224, uc_2225, uc_2226, uc_2227, uc_2228, uc_2229, uc_2230, 
      uc_2231, uc_2232, uc_2233, uc_2234, uc_2235, uc_2236, uc_2237, uc_2238, 
      uc_2239, uc_2240, uc_2241, uc_2242, uc_2243, uc_2244, uc_2245, uc_2246, 
      uc_2247, uc_2248, uc_2249, uc_2250, uc_2251, uc_2252, uc_2253, uc_2254, 
      uc_2255, normalizedWires[1193], normalizedWires[1192], 
      normalizedWires[1191], normalizedWires[1190], normalizedWires[1189], 
      normalizedWires[1188], normalizedWires[1187], normalizedWires[1186], 
      normalizedWires[1185], normalizedWires[1184], normalizedWires[1183], 
      normalizedWires[1182], normalizedWires[1181], normalizedWires[1180], 
      normalizedWires[1179], normalizedWires[1178], normalizedWires[1177], 
      normalizedWires[1176], normalizedWires[1175], normalizedWires[1174], 
      normalizedWires[1173], normalizedWires[1172], normalizedWires[1171], 
      normalizedWires[1170], uc_2256, uc_2257, uc_2258, uc_2259, uc_2260, 
      uc_2261, uc_2262, uc_2263, uc_2264, uc_2265, uc_2266, uc_2267, uc_2268, 
      uc_2269, uc_2270, uc_2271, uc_2272, uc_2273, uc_2274, uc_2275, uc_2276, 
      uc_2277, uc_2278, uc_2279, uc_2280, uc_2281, uc_2282, uc_2283, uc_2284, 
      uc_2285, uc_2286, uc_2287, uc_2288, uc_2289, uc_2290, uc_2291, uc_2292, 
      uc_2293, uc_2294, uc_2295, uc_2296, normalizedWires[1128], 
      normalizedWires[1127], normalizedWires[1126], normalizedWires[1125], 
      normalizedWires[1124], normalizedWires[1123], normalizedWires[1122], 
      normalizedWires[1121], normalizedWires[1120], normalizedWires[1119], 
      normalizedWires[1118], normalizedWires[1117], normalizedWires[1116], 
      normalizedWires[1115], normalizedWires[1114], normalizedWires[1113], 
      normalizedWires[1112], normalizedWires[1111], normalizedWires[1110], 
      normalizedWires[1109], normalizedWires[1108], normalizedWires[1107], 
      normalizedWires[1106], normalizedWires[1105], uc_2297, uc_2298, uc_2299, 
      uc_2300, uc_2301, uc_2302, uc_2303, uc_2304, uc_2305, uc_2306, uc_2307, 
      uc_2308, uc_2309, uc_2310, uc_2311, uc_2312, uc_2313, uc_2314, uc_2315, 
      uc_2316, uc_2317, uc_2318, uc_2319, uc_2320, uc_2321, uc_2322, uc_2323, 
      uc_2324, uc_2325, uc_2326, uc_2327, uc_2328, uc_2329, uc_2330, uc_2331, 
      uc_2332, uc_2333, uc_2334, uc_2335, uc_2336, uc_2337, 
      normalizedWires[1063], normalizedWires[1062], normalizedWires[1061], 
      normalizedWires[1060], normalizedWires[1059], normalizedWires[1058], 
      normalizedWires[1057], normalizedWires[1056], normalizedWires[1055], 
      normalizedWires[1054], normalizedWires[1053], normalizedWires[1052], 
      normalizedWires[1051], normalizedWires[1050], normalizedWires[1049], 
      normalizedWires[1048], normalizedWires[1047], normalizedWires[1046], 
      normalizedWires[1045], normalizedWires[1044], normalizedWires[1043], 
      normalizedWires[1042], normalizedWires[1041], normalizedWires[1040], 
      uc_2338, uc_2339, uc_2340, uc_2341, uc_2342, uc_2343, uc_2344, uc_2345, 
      uc_2346, uc_2347, uc_2348, uc_2349, uc_2350, uc_2351, uc_2352, uc_2353, 
      uc_2354, uc_2355, uc_2356, uc_2357, uc_2358, uc_2359, uc_2360, uc_2361, 
      uc_2362, uc_2363, uc_2364, uc_2365, uc_2366, uc_2367, uc_2368, uc_2369, 
      uc_2370, uc_2371, uc_2372, uc_2373, uc_2374, uc_2375, uc_2376, uc_2377, 
      uc_2378, normalizedWires[998], normalizedWires[997], normalizedWires[996], 
      normalizedWires[995], normalizedWires[994], normalizedWires[993], 
      normalizedWires[992], normalizedWires[991], normalizedWires[990], 
      normalizedWires[989], normalizedWires[988], normalizedWires[987], 
      normalizedWires[986], normalizedWires[985], normalizedWires[984], 
      normalizedWires[983], normalizedWires[982], normalizedWires[981], 
      normalizedWires[980], normalizedWires[979], normalizedWires[978], 
      normalizedWires[977], normalizedWires[976], normalizedWires[975], uc_2379, 
      uc_2380, uc_2381, uc_2382, uc_2383, uc_2384, uc_2385, uc_2386, uc_2387, 
      uc_2388, uc_2389, uc_2390, uc_2391, uc_2392, uc_2393, uc_2394, uc_2395, 
      uc_2396, uc_2397, uc_2398, uc_2399, uc_2400, uc_2401, uc_2402, uc_2403, 
      uc_2404, uc_2405, uc_2406, uc_2407, uc_2408, uc_2409, uc_2410, uc_2411, 
      uc_2412, uc_2413, uc_2414, uc_2415, uc_2416, uc_2417, uc_2418, uc_2419, 
      normalizedWires[933], normalizedWires[932], normalizedWires[931], 
      normalizedWires[930], normalizedWires[929], normalizedWires[928], 
      normalizedWires[927], normalizedWires[926], normalizedWires[925], 
      normalizedWires[924], normalizedWires[923], normalizedWires[922], 
      normalizedWires[921], normalizedWires[920], normalizedWires[919], 
      normalizedWires[918], normalizedWires[917], normalizedWires[916], 
      normalizedWires[915], normalizedWires[914], normalizedWires[913], 
      normalizedWires[912], normalizedWires[911], normalizedWires[910], uc_2420, 
      uc_2421, uc_2422, uc_2423, uc_2424, uc_2425, uc_2426, uc_2427, uc_2428, 
      uc_2429, uc_2430, uc_2431, uc_2432, uc_2433, uc_2434, uc_2435, uc_2436, 
      uc_2437, uc_2438, uc_2439, uc_2440, uc_2441, uc_2442, uc_2443, uc_2444, 
      uc_2445, uc_2446, uc_2447, uc_2448, uc_2449, uc_2450, uc_2451, uc_2452, 
      uc_2453, uc_2454, uc_2455, uc_2456, uc_2457, uc_2458, uc_2459, uc_2460, 
      normalizedWires[868], normalizedWires[867], normalizedWires[866], 
      normalizedWires[865], normalizedWires[864], normalizedWires[863], 
      normalizedWires[862], normalizedWires[861], normalizedWires[860], 
      normalizedWires[859], normalizedWires[858], normalizedWires[857], 
      normalizedWires[856], normalizedWires[855], normalizedWires[854], 
      normalizedWires[853], normalizedWires[852], normalizedWires[851], 
      normalizedWires[850], normalizedWires[849], normalizedWires[848], 
      normalizedWires[847], normalizedWires[846], normalizedWires[845], uc_2461, 
      uc_2462, uc_2463, uc_2464, uc_2465, uc_2466, uc_2467, uc_2468, uc_2469, 
      uc_2470, uc_2471, uc_2472, uc_2473, uc_2474, uc_2475, uc_2476, uc_2477, 
      uc_2478, uc_2479, uc_2480, uc_2481, uc_2482, uc_2483, uc_2484, uc_2485, 
      uc_2486, uc_2487, uc_2488, uc_2489, uc_2490, uc_2491, uc_2492, uc_2493, 
      uc_2494, uc_2495, uc_2496, uc_2497, uc_2498, uc_2499, uc_2500, uc_2501, 
      normalizedWires[803], normalizedWires[802], normalizedWires[801], 
      normalizedWires[800], normalizedWires[799], normalizedWires[798], 
      normalizedWires[797], normalizedWires[796], normalizedWires[795], 
      normalizedWires[794], normalizedWires[793], normalizedWires[792], 
      normalizedWires[791], normalizedWires[790], normalizedWires[789], 
      normalizedWires[788], normalizedWires[787], normalizedWires[786], 
      normalizedWires[785], normalizedWires[784], normalizedWires[783], 
      normalizedWires[782], normalizedWires[781], normalizedWires[780], uc_2502, 
      uc_2503, uc_2504, uc_2505, uc_2506, uc_2507, uc_2508, uc_2509, uc_2510, 
      uc_2511, uc_2512, uc_2513, uc_2514, uc_2515, uc_2516, uc_2517, uc_2518, 
      uc_2519, uc_2520, uc_2521, uc_2522, uc_2523, uc_2524, uc_2525, uc_2526, 
      uc_2527, uc_2528, uc_2529, uc_2530, uc_2531, uc_2532, uc_2533, uc_2534, 
      uc_2535, uc_2536, uc_2537, uc_2538, uc_2539, uc_2540, uc_2541, uc_2542, 
      normalizedWires[738], normalizedWires[737], normalizedWires[736], 
      normalizedWires[735], normalizedWires[734], normalizedWires[733], 
      normalizedWires[732], normalizedWires[731], normalizedWires[730], 
      normalizedWires[729], normalizedWires[728], normalizedWires[727], 
      normalizedWires[726], normalizedWires[725], normalizedWires[724], 
      normalizedWires[723], normalizedWires[722], normalizedWires[721], 
      normalizedWires[720], normalizedWires[719], normalizedWires[718], 
      normalizedWires[717], normalizedWires[716], normalizedWires[715], uc_2543, 
      uc_2544, uc_2545, uc_2546, uc_2547, uc_2548, uc_2549, uc_2550, uc_2551, 
      uc_2552, uc_2553, uc_2554, uc_2555, uc_2556, uc_2557, uc_2558, uc_2559, 
      uc_2560, uc_2561, uc_2562, uc_2563, uc_2564, uc_2565, uc_2566, uc_2567, 
      uc_2568, uc_2569, uc_2570, uc_2571, uc_2572, uc_2573, uc_2574, uc_2575, 
      uc_2576, uc_2577, uc_2578, uc_2579, uc_2580, uc_2581, uc_2582, uc_2583, 
      normalizedWires[673], normalizedWires[672], normalizedWires[671], 
      normalizedWires[670], normalizedWires[669], normalizedWires[668], 
      normalizedWires[667], normalizedWires[666], normalizedWires[665], 
      normalizedWires[664], normalizedWires[663], normalizedWires[662], 
      normalizedWires[661], normalizedWires[660], normalizedWires[659], 
      normalizedWires[658], normalizedWires[657], normalizedWires[656], 
      normalizedWires[655], normalizedWires[654], normalizedWires[653], 
      normalizedWires[652], normalizedWires[651], normalizedWires[650], uc_2584, 
      uc_2585, uc_2586, uc_2587, uc_2588, uc_2589, uc_2590, uc_2591, uc_2592, 
      uc_2593, uc_2594, uc_2595, uc_2596, uc_2597, uc_2598, uc_2599, uc_2600, 
      uc_2601, uc_2602, uc_2603, uc_2604, uc_2605, uc_2606, uc_2607, uc_2608, 
      uc_2609, uc_2610, uc_2611, uc_2612, uc_2613, uc_2614, uc_2615, uc_2616, 
      uc_2617, uc_2618, uc_2619, uc_2620, uc_2621, uc_2622, uc_2623, uc_2624, 
      normalizedWires[608], normalizedWires[607], normalizedWires[606], 
      normalizedWires[605], normalizedWires[604], normalizedWires[603], 
      normalizedWires[602], normalizedWires[601], normalizedWires[600], 
      normalizedWires[599], normalizedWires[598], normalizedWires[597], 
      normalizedWires[596], normalizedWires[595], normalizedWires[594], 
      normalizedWires[593], normalizedWires[592], normalizedWires[591], 
      normalizedWires[590], normalizedWires[589], normalizedWires[588], 
      normalizedWires[587], normalizedWires[586], normalizedWires[585], uc_2625, 
      uc_2626, uc_2627, uc_2628, uc_2629, uc_2630, uc_2631, uc_2632, uc_2633, 
      uc_2634, uc_2635, uc_2636, uc_2637, uc_2638, uc_2639, uc_2640, uc_2641, 
      uc_2642, uc_2643, uc_2644, uc_2645, uc_2646, uc_2647, uc_2648, uc_2649, 
      uc_2650, uc_2651, uc_2652, uc_2653, uc_2654, uc_2655, uc_2656, uc_2657, 
      uc_2658, uc_2659, uc_2660, uc_2661, uc_2662, uc_2663, uc_2664, uc_2665, 
      normalizedWires[543], normalizedWires[542], normalizedWires[541], 
      normalizedWires[540], normalizedWires[539], normalizedWires[538], 
      normalizedWires[537], normalizedWires[536], normalizedWires[535], 
      normalizedWires[534], normalizedWires[533], normalizedWires[532], 
      normalizedWires[531], normalizedWires[530], normalizedWires[529], 
      normalizedWires[528], normalizedWires[527], normalizedWires[526], 
      normalizedWires[525], normalizedWires[524], normalizedWires[523], 
      normalizedWires[522], normalizedWires[521], normalizedWires[520], uc_2666, 
      uc_2667, uc_2668, uc_2669, uc_2670, uc_2671, uc_2672, uc_2673, uc_2674, 
      uc_2675, uc_2676, uc_2677, uc_2678, uc_2679, uc_2680, uc_2681, uc_2682, 
      uc_2683, uc_2684, uc_2685, uc_2686, uc_2687, uc_2688, uc_2689, uc_2690, 
      uc_2691, uc_2692, uc_2693, uc_2694, uc_2695, uc_2696, uc_2697, uc_2698, 
      uc_2699, uc_2700, uc_2701, uc_2702, uc_2703, uc_2704, uc_2705, uc_2706, 
      normalizedWires[478], normalizedWires[477], normalizedWires[476], 
      normalizedWires[475], normalizedWires[474], normalizedWires[473], 
      normalizedWires[472], normalizedWires[471], normalizedWires[470], 
      normalizedWires[469], normalizedWires[468], normalizedWires[467], 
      normalizedWires[466], normalizedWires[465], normalizedWires[464], 
      normalizedWires[463], normalizedWires[462], normalizedWires[461], 
      normalizedWires[460], normalizedWires[459], normalizedWires[458], 
      normalizedWires[457], normalizedWires[456], normalizedWires[455], uc_2707, 
      uc_2708, uc_2709, uc_2710, uc_2711, uc_2712, uc_2713, uc_2714, uc_2715, 
      uc_2716, uc_2717, uc_2718, uc_2719, uc_2720, uc_2721, uc_2722, uc_2723, 
      uc_2724, uc_2725, uc_2726, uc_2727, uc_2728, uc_2729, uc_2730, uc_2731, 
      uc_2732, uc_2733, uc_2734, uc_2735, uc_2736, uc_2737, uc_2738, uc_2739, 
      uc_2740, uc_2741, uc_2742, uc_2743, uc_2744, uc_2745, uc_2746, uc_2747, 
      normalizedWires[413], normalizedWires[412], normalizedWires[411], 
      normalizedWires[410], normalizedWires[409], normalizedWires[408], 
      normalizedWires[407], normalizedWires[406], normalizedWires[405], 
      normalizedWires[404], normalizedWires[403], normalizedWires[402], 
      normalizedWires[401], normalizedWires[400], normalizedWires[399], 
      normalizedWires[398], normalizedWires[397], normalizedWires[396], 
      normalizedWires[395], normalizedWires[394], normalizedWires[393], 
      normalizedWires[392], normalizedWires[391], normalizedWires[390], uc_2748, 
      uc_2749, uc_2750, uc_2751, uc_2752, uc_2753, uc_2754, uc_2755, uc_2756, 
      uc_2757, uc_2758, uc_2759, uc_2760, uc_2761, uc_2762, uc_2763, uc_2764, 
      uc_2765, uc_2766, uc_2767, uc_2768, uc_2769, uc_2770, uc_2771, uc_2772, 
      uc_2773, uc_2774, uc_2775, uc_2776, uc_2777, uc_2778, uc_2779, uc_2780, 
      uc_2781, uc_2782, uc_2783, uc_2784, uc_2785, uc_2786, uc_2787, uc_2788, 
      normalizedWires[348], normalizedWires[347], normalizedWires[346], 
      normalizedWires[345], normalizedWires[344], normalizedWires[343], 
      normalizedWires[342], normalizedWires[341], normalizedWires[340], 
      normalizedWires[339], normalizedWires[338], normalizedWires[337], 
      normalizedWires[336], normalizedWires[335], normalizedWires[334], 
      normalizedWires[333], normalizedWires[332], normalizedWires[331], 
      normalizedWires[330], normalizedWires[329], normalizedWires[328], 
      normalizedWires[327], normalizedWires[326], normalizedWires[325], uc_2789, 
      uc_2790, uc_2791, uc_2792, uc_2793, uc_2794, uc_2795, uc_2796, uc_2797, 
      uc_2798, uc_2799, uc_2800, uc_2801, uc_2802, uc_2803, uc_2804, uc_2805, 
      uc_2806, uc_2807, uc_2808, uc_2809, uc_2810, uc_2811, uc_2812, uc_2813, 
      uc_2814, uc_2815, uc_2816, uc_2817, uc_2818, uc_2819, uc_2820, uc_2821, 
      uc_2822, uc_2823, uc_2824, uc_2825, uc_2826, uc_2827, uc_2828, uc_2829, 
      normalizedWires[283], normalizedWires[282], normalizedWires[281], 
      normalizedWires[280], normalizedWires[279], normalizedWires[278], 
      normalizedWires[277], normalizedWires[276], normalizedWires[275], 
      normalizedWires[274], normalizedWires[273], normalizedWires[272], 
      normalizedWires[271], normalizedWires[270], normalizedWires[269], 
      normalizedWires[268], normalizedWires[267], normalizedWires[266], 
      normalizedWires[265], normalizedWires[264], normalizedWires[263], 
      normalizedWires[262], normalizedWires[261], normalizedWires[260], uc_2830, 
      uc_2831, uc_2832, uc_2833, uc_2834, uc_2835, uc_2836, uc_2837, uc_2838, 
      uc_2839, uc_2840, uc_2841, uc_2842, uc_2843, uc_2844, uc_2845, uc_2846, 
      uc_2847, uc_2848, uc_2849, uc_2850, uc_2851, uc_2852, uc_2853, uc_2854, 
      uc_2855, uc_2856, uc_2857, uc_2858, uc_2859, uc_2860, uc_2861, uc_2862, 
      uc_2863, uc_2864, uc_2865, uc_2866, uc_2867, uc_2868, uc_2869, uc_2870, 
      normalizedWires[218], normalizedWires[217], normalizedWires[216], 
      normalizedWires[215], normalizedWires[214], normalizedWires[213], 
      normalizedWires[212], normalizedWires[211], normalizedWires[210], 
      normalizedWires[209], normalizedWires[208], normalizedWires[207], 
      normalizedWires[206], normalizedWires[205], normalizedWires[204], 
      normalizedWires[203], normalizedWires[202], normalizedWires[201], 
      normalizedWires[200], normalizedWires[199], normalizedWires[198], 
      normalizedWires[197], normalizedWires[196], normalizedWires[195], uc_2871, 
      uc_2872, uc_2873, uc_2874, uc_2875, uc_2876, uc_2877, uc_2878, uc_2879, 
      uc_2880, uc_2881, uc_2882, uc_2883, uc_2884, uc_2885, uc_2886, uc_2887, 
      uc_2888, uc_2889, uc_2890, uc_2891, uc_2892, uc_2893, uc_2894, uc_2895, 
      uc_2896, uc_2897, uc_2898, uc_2899, uc_2900, uc_2901, uc_2902, uc_2903, 
      uc_2904, uc_2905, uc_2906, uc_2907, uc_2908, uc_2909, uc_2910, uc_2911, 
      normalizedWires[153], normalizedWires[152], normalizedWires[151], 
      normalizedWires[150], normalizedWires[149], normalizedWires[148], 
      normalizedWires[147], normalizedWires[146], normalizedWires[145], 
      normalizedWires[144], normalizedWires[143], normalizedWires[142], 
      normalizedWires[141], normalizedWires[140], normalizedWires[139], 
      normalizedWires[138], normalizedWires[137], normalizedWires[136], 
      normalizedWires[135], normalizedWires[134], normalizedWires[133], 
      normalizedWires[132], normalizedWires[131], normalizedWires[130], uc_2912, 
      uc_2913, uc_2914, uc_2915, uc_2916, uc_2917, uc_2918, uc_2919, uc_2920, 
      uc_2921, uc_2922, uc_2923, uc_2924, uc_2925, uc_2926, uc_2927, uc_2928, 
      uc_2929, uc_2930, uc_2931, uc_2932, uc_2933, uc_2934, uc_2935, uc_2936, 
      uc_2937, uc_2938, uc_2939, uc_2940, uc_2941, uc_2942, uc_2943, uc_2944, 
      uc_2945, uc_2946, uc_2947, uc_2948, uc_2949, uc_2950, uc_2951, uc_2952, 
      normalizedWires[88], normalizedWires[87], normalizedWires[86], 
      normalizedWires[85], normalizedWires[84], normalizedWires[83], 
      normalizedWires[82], normalizedWires[81], normalizedWires[80], 
      normalizedWires[79], normalizedWires[78], normalizedWires[77], 
      normalizedWires[76], normalizedWires[75], normalizedWires[74], 
      normalizedWires[73], normalizedWires[72], normalizedWires[71], 
      normalizedWires[70], normalizedWires[69], normalizedWires[68], 
      normalizedWires[67], normalizedWires[66], normalizedWires[65], uc_2953, 
      uc_2954, uc_2955, uc_2956, uc_2957, uc_2958, uc_2959, uc_2960, uc_2961, 
      uc_2962, uc_2963, uc_2964, uc_2965, uc_2966, uc_2967, uc_2968, uc_2969, 
      uc_2970, uc_2971, uc_2972, uc_2973, uc_2974, uc_2975, uc_2976, uc_2977, 
      uc_2978, uc_2979, uc_2980, uc_2981, uc_2982, uc_2983, uc_2984, uc_2985, 
      uc_2986, uc_2987, uc_2988, uc_2989, uc_2990, uc_2991, uc_2992, uc_2993, 
      normalizedWires[23], normalizedWires[22], normalizedWires[21], 
      normalizedWires[20], normalizedWires[19], normalizedWires[18], 
      normalizedWires[17], normalizedWires[16], normalizedWires[15], 
      normalizedWires[14], normalizedWires[13], normalizedWires[12], 
      normalizedWires[11], normalizedWires[10], normalizedWires[9], 
      normalizedWires[8], normalizedWires[7], normalizedWires[6], 
      normalizedWires[5], normalizedWires[4], normalizedWires[3], 
      normalizedWires[2], normalizedWires[1], uc_2994}), .A({uc_2995, uc_2996, 
      uc_2997, uc_2998, uc_2999, uc_3000, uc_3001, uc_3002, 
      normalizedWires[1518], n_0_24, n_0_25, n_0_26, n_0_27, n_0_28, n_0_29, 
      n_0_30, n_0_31, n_0_32, n_0_33, n_0_34, n_0_35, n_0_36, n_0_37, n_0_38, 
      n_0_39, n_0_40, n_0_41, n_0_42, n_0_43, n_0_44, n_0_45, n_0_1}), .B({
      uc_3003, uc_3004, uc_3005, uc_3006, uc_3007, uc_3008, uc_3009, uc_3010, 
      uc_3011, n_0_2, n_0_3, n_0_4, n_0_5, n_0_6, n_0_7, n_0_8, n_0_9, n_0_10, 
      n_0_11, n_0_12, n_0_13, n_0_14, n_0_15, n_0_16, n_0_17, n_0_18, n_0_19, 
      n_0_20, n_0_21, n_0_22, n_0_23, n_0_0}));
   addResWithCarry thirdStage (.Res_out({uc_3012, uc_3013, uc_3014, uc_3015, 
      uc_3016, uc_3017, uc_3018, uc_3019, uc_3020, uc_3021, uc_3022, uc_3023, 
      uc_3024, uc_3025, uc_3026, uc_3027, Res_imm[47], Res_imm[46], Res_imm[45], 
      Res_imm[44], Res_imm[43], Res_imm[42], Res_imm[41], Res_imm[40], 
      Res_imm[39], Res_imm[38], Res_imm[37], Res_imm[36], Res_imm[35], 
      Res_imm[34], Res_imm[33], Res_imm[32], Res_imm[31], Res_imm[30], 
      Res_imm[29], Res_imm[28], Res_imm[27], Res_imm[26], Res_imm[25], 
      Res_imm[24], Res_imm[23], uc_3028, uc_3029, uc_3030, uc_3031, uc_3032, 
      uc_3033, uc_3034, uc_3035, uc_3036, uc_3037, uc_3038, uc_3039, uc_3040, 
      uc_3041, uc_3042, uc_3043, uc_3044, uc_3045, uc_3046, uc_3047, uc_3048, 
      uc_3049, uc_3050}), .Res_in({uc_3051, uc_3052, uc_3053, uc_3054, uc_3055, 
      uc_3056, uc_3057, uc_3058, uc_3059, uc_3060, uc_3061, uc_3062, uc_3063, 
      uc_3064, uc_3065, uc_3066, secondStage_Res[47], secondStage_Res[46], 
      secondStage_Res[45], secondStage_Res[44], secondStage_Res[43], 
      secondStage_Res[42], secondStage_Res[41], secondStage_Res[40], 
      secondStage_Res[39], secondStage_Res[38], secondStage_Res[37], 
      secondStage_Res[36], secondStage_Res[35], secondStage_Res[34], 
      secondStage_Res[33], secondStage_Res[32], secondStage_Res[31], 
      secondStage_Res[30], secondStage_Res[29], secondStage_Res[28], 
      secondStage_Res[27], secondStage_Res[26], secondStage_Res[25], 
      secondStage_Res[24], secondStage_Res[23], secondStage_Res[22], 
      secondStage_Res[21], secondStage_Res[20], secondStage_Res[19], 
      secondStage_Res[18], secondStage_Res[17], secondStage_Res[16], 
      secondStage_Res[15], secondStage_Res[14], secondStage_Res[13], 
      secondStage_Res[12], secondStage_Res[11], secondStage_Res[10], 
      secondStage_Res[9], uc_3067, uc_3068, uc_3069, uc_3070, uc_3071, uc_3072, 
      uc_3073, uc_3074, uc_3075}), .carry_in({uc_3076, uc_3077, uc_3078, uc_3079, 
      uc_3080, uc_3081, uc_3082, uc_3083, uc_3084, uc_3085, uc_3086, uc_3087, 
      uc_3088, uc_3089, uc_3090, uc_3091, secondStage_carry[47], 
      secondStage_carry[46], secondStage_carry[45], secondStage_carry[44], 
      secondStage_carry[43], secondStage_carry[42], secondStage_carry[41], 
      secondStage_carry[40], secondStage_carry[39], secondStage_carry[38], 
      secondStage_carry[37], secondStage_carry[36], secondStage_carry[35], 
      secondStage_carry[34], secondStage_carry[33], secondStage_carry[32], 
      secondStage_carry[31], secondStage_carry[30], secondStage_carry[29], 
      secondStage_carry[28], secondStage_carry[27], secondStage_carry[26], 
      secondStage_carry[25], secondStage_carry[24], secondStage_carry[23], 
      secondStage_carry[22], secondStage_carry[21], secondStage_carry[20], 
      secondStage_carry[19], secondStage_carry[18], secondStage_carry[17], 
      secondStage_carry[16], secondStage_carry[15], secondStage_carry[14], 
      secondStage_carry[13], secondStage_carry[12], secondStage_carry[11], 
      secondStage_carry[10], secondStage_carry[9], uc_3092, uc_3093, uc_3094, 
      uc_3095, uc_3096, uc_3097, uc_3098, uc_3099, uc_3100}));
   DLH_X1 \Res_reg[47]  (.D(n_0_70), .G(n_0_119), .Q(Res[47]));
   DLH_X1 \Res_reg[46]  (.D(n_0_69), .G(n_0_119), .Q(Res[46]));
   DLH_X1 \Res_reg[45]  (.D(n_0_68), .G(n_0_119), .Q(Res[45]));
   DLH_X1 \Res_reg[44]  (.D(n_0_67), .G(n_0_119), .Q(Res[44]));
   DLH_X1 \Res_reg[43]  (.D(n_0_66), .G(n_0_119), .Q(Res[43]));
   DLH_X1 \Res_reg[42]  (.D(n_0_65), .G(n_0_119), .Q(Res[42]));
   DLH_X1 \Res_reg[41]  (.D(n_0_64), .G(n_0_119), .Q(Res[41]));
   DLH_X1 \Res_reg[40]  (.D(n_0_63), .G(n_0_119), .Q(Res[40]));
   DLH_X1 \Res_reg[39]  (.D(n_0_62), .G(n_0_119), .Q(Res[39]));
   DLH_X1 \Res_reg[38]  (.D(n_0_61), .G(n_0_119), .Q(Res[38]));
   DLH_X1 \Res_reg[37]  (.D(n_0_60), .G(n_0_119), .Q(Res[37]));
   DLH_X1 \Res_reg[36]  (.D(n_0_59), .G(n_0_119), .Q(Res[36]));
   DLH_X1 \Res_reg[35]  (.D(n_0_58), .G(n_0_119), .Q(Res[35]));
   DLH_X1 \Res_reg[34]  (.D(n_0_57), .G(n_0_119), .Q(Res[34]));
   DLH_X1 \Res_reg[33]  (.D(n_0_56), .G(n_0_119), .Q(Res[33]));
   DLH_X1 \Res_reg[32]  (.D(n_0_55), .G(n_0_119), .Q(Res[32]));
   DLH_X1 \Res_reg[31]  (.D(n_0_54), .G(n_0_119), .Q(Res[31]));
   DLH_X1 \Res_reg[30]  (.D(n_0_53), .G(n_0_119), .Q(Res[30]));
   DLH_X1 \Res_reg[29]  (.D(n_0_52), .G(n_0_119), .Q(Res[29]));
   DLH_X1 \Res_reg[28]  (.D(n_0_51), .G(n_0_119), .Q(Res[28]));
   DLH_X1 \Res_reg[27]  (.D(n_0_50), .G(n_0_119), .Q(Res[27]));
   DLH_X1 \Res_reg[26]  (.D(n_0_49), .G(n_0_119), .Q(Res[26]));
   DLH_X1 \Res_reg[25]  (.D(n_0_48), .G(n_0_119), .Q(Res[25]));
   DLH_X1 \Res_reg[24]  (.D(n_0_47), .G(n_0_119), .Q(Res[24]));
   DLH_X1 \Res_reg[23]  (.D(n_0_46), .G(n_0_119), .Q(Res[23]));
   DLH_X1 \B_in_reg[22]  (.D(n_0_117), .G(n_0_94), .Q(n_0_2));
   DLH_X1 \B_in_reg[21]  (.D(n_0_116), .G(n_0_94), .Q(n_0_3));
   DLH_X1 \B_in_reg[20]  (.D(n_0_115), .G(n_0_94), .Q(n_0_4));
   DLH_X1 \B_in_reg[19]  (.D(n_0_114), .G(n_0_94), .Q(n_0_5));
   DLH_X1 \B_in_reg[18]  (.D(n_0_113), .G(n_0_94), .Q(n_0_6));
   DLH_X1 \B_in_reg[17]  (.D(n_0_112), .G(n_0_94), .Q(n_0_7));
   DLH_X1 \B_in_reg[16]  (.D(n_0_111), .G(n_0_94), .Q(n_0_8));
   DLH_X1 \B_in_reg[15]  (.D(n_0_110), .G(n_0_94), .Q(n_0_9));
   DLH_X1 \B_in_reg[14]  (.D(n_0_109), .G(n_0_94), .Q(n_0_10));
   DLH_X1 \B_in_reg[13]  (.D(n_0_108), .G(n_0_94), .Q(n_0_11));
   DLH_X1 \B_in_reg[12]  (.D(n_0_107), .G(n_0_94), .Q(n_0_12));
   DLH_X1 \B_in_reg[11]  (.D(n_0_106), .G(n_0_94), .Q(n_0_13));
   DLH_X1 \B_in_reg[10]  (.D(n_0_105), .G(n_0_94), .Q(n_0_14));
   DLH_X1 \B_in_reg[9]  (.D(n_0_104), .G(n_0_94), .Q(n_0_15));
   DLH_X1 \B_in_reg[8]  (.D(n_0_103), .G(n_0_94), .Q(n_0_16));
   DLH_X1 \B_in_reg[7]  (.D(n_0_102), .G(n_0_94), .Q(n_0_17));
   DLH_X1 \B_in_reg[6]  (.D(n_0_101), .G(n_0_94), .Q(n_0_18));
   DLH_X1 \B_in_reg[5]  (.D(n_0_100), .G(n_0_94), .Q(n_0_19));
   DLH_X1 \B_in_reg[4]  (.D(n_0_99), .G(n_0_94), .Q(n_0_20));
   DLH_X1 \B_in_reg[3]  (.D(n_0_98), .G(n_0_94), .Q(n_0_21));
   DLH_X1 \B_in_reg[2]  (.D(n_0_97), .G(n_0_94), .Q(n_0_22));
   DLH_X1 \B_in_reg[1]  (.D(n_0_96), .G(n_0_94), .Q(n_0_23));
   DLH_X1 \B_in_reg[0]  (.D(n_0_95), .G(n_0_94), .Q(n_0_0));
   DLH_X1 \A_in_reg[22]  (.D(n_0_93), .G(n_0_94), .Q(n_0_24));
   DLH_X1 \A_in_reg[21]  (.D(n_0_92), .G(n_0_94), .Q(n_0_25));
   DLH_X1 \A_in_reg[20]  (.D(n_0_91), .G(n_0_94), .Q(n_0_26));
   DLH_X1 \A_in_reg[19]  (.D(n_0_90), .G(n_0_94), .Q(n_0_27));
   DLH_X1 \A_in_reg[18]  (.D(n_0_89), .G(n_0_94), .Q(n_0_28));
   DLH_X1 \A_in_reg[17]  (.D(n_0_88), .G(n_0_94), .Q(n_0_29));
   DLH_X1 \A_in_reg[16]  (.D(n_0_87), .G(n_0_94), .Q(n_0_30));
   DLH_X1 \A_in_reg[15]  (.D(n_0_86), .G(n_0_94), .Q(n_0_31));
   DLH_X1 \A_in_reg[14]  (.D(n_0_85), .G(n_0_94), .Q(n_0_32));
   DLH_X1 \A_in_reg[13]  (.D(n_0_84), .G(n_0_94), .Q(n_0_33));
   DLH_X1 \A_in_reg[12]  (.D(n_0_83), .G(n_0_94), .Q(n_0_34));
   DLH_X1 \A_in_reg[11]  (.D(n_0_82), .G(n_0_94), .Q(n_0_35));
   DLH_X1 \A_in_reg[10]  (.D(n_0_81), .G(n_0_94), .Q(n_0_36));
   DLH_X1 \A_in_reg[9]  (.D(n_0_80), .G(n_0_94), .Q(n_0_37));
   DLH_X1 \A_in_reg[8]  (.D(n_0_79), .G(n_0_94), .Q(n_0_38));
   DLH_X1 \A_in_reg[7]  (.D(n_0_78), .G(n_0_94), .Q(n_0_39));
   DLH_X1 \A_in_reg[6]  (.D(n_0_77), .G(n_0_94), .Q(n_0_40));
   DLH_X1 \A_in_reg[5]  (.D(n_0_76), .G(n_0_94), .Q(n_0_41));
   DLH_X1 \A_in_reg[4]  (.D(n_0_75), .G(n_0_94), .Q(n_0_42));
   DLH_X1 \A_in_reg[3]  (.D(n_0_74), .G(n_0_94), .Q(n_0_43));
   DLH_X1 \A_in_reg[2]  (.D(n_0_73), .G(n_0_94), .Q(n_0_44));
   DLH_X1 \A_in_reg[1]  (.D(n_0_72), .G(n_0_94), .Q(n_0_45));
   DLH_X1 \A_in_reg[0]  (.D(n_0_71), .G(n_0_94), .Q(n_0_1));
   DLH_X1 \B_in_reg[23]  (.D(n_0_118), .G(n_0_94), .Q(normalizedWires[1518]));
   AND2_X1 i_0_0_0 (.A1(n_0_118), .A2(Res_imm[23]), .ZN(n_0_46));
   AND2_X1 i_0_0_1 (.A1(n_0_118), .A2(Res_imm[24]), .ZN(n_0_47));
   AND2_X1 i_0_0_2 (.A1(n_0_118), .A2(Res_imm[25]), .ZN(n_0_48));
   AND2_X1 i_0_0_3 (.A1(n_0_118), .A2(Res_imm[26]), .ZN(n_0_49));
   AND2_X1 i_0_0_4 (.A1(n_0_118), .A2(Res_imm[27]), .ZN(n_0_50));
   AND2_X1 i_0_0_5 (.A1(n_0_118), .A2(Res_imm[28]), .ZN(n_0_51));
   AND2_X1 i_0_0_6 (.A1(n_0_118), .A2(Res_imm[29]), .ZN(n_0_52));
   AND2_X1 i_0_0_7 (.A1(n_0_118), .A2(Res_imm[30]), .ZN(n_0_53));
   AND2_X1 i_0_0_8 (.A1(n_0_118), .A2(Res_imm[31]), .ZN(n_0_54));
   AND2_X1 i_0_0_9 (.A1(n_0_118), .A2(Res_imm[32]), .ZN(n_0_55));
   AND2_X1 i_0_0_10 (.A1(n_0_118), .A2(Res_imm[33]), .ZN(n_0_56));
   AND2_X1 i_0_0_11 (.A1(n_0_118), .A2(Res_imm[34]), .ZN(n_0_57));
   AND2_X1 i_0_0_12 (.A1(n_0_118), .A2(Res_imm[35]), .ZN(n_0_58));
   AND2_X1 i_0_0_13 (.A1(n_0_118), .A2(Res_imm[36]), .ZN(n_0_59));
   AND2_X1 i_0_0_14 (.A1(n_0_118), .A2(Res_imm[37]), .ZN(n_0_60));
   AND2_X1 i_0_0_15 (.A1(n_0_118), .A2(Res_imm[38]), .ZN(n_0_61));
   AND2_X1 i_0_0_16 (.A1(n_0_118), .A2(Res_imm[39]), .ZN(n_0_62));
   AND2_X1 i_0_0_17 (.A1(n_0_118), .A2(Res_imm[40]), .ZN(n_0_63));
   AND2_X1 i_0_0_18 (.A1(n_0_118), .A2(Res_imm[41]), .ZN(n_0_64));
   AND2_X1 i_0_0_19 (.A1(n_0_118), .A2(Res_imm[42]), .ZN(n_0_65));
   AND2_X1 i_0_0_20 (.A1(n_0_118), .A2(Res_imm[43]), .ZN(n_0_66));
   AND2_X1 i_0_0_21 (.A1(n_0_118), .A2(Res_imm[44]), .ZN(n_0_67));
   AND2_X1 i_0_0_22 (.A1(n_0_118), .A2(Res_imm[45]), .ZN(n_0_68));
   AND2_X1 i_0_0_23 (.A1(n_0_118), .A2(Res_imm[46]), .ZN(n_0_69));
   AND2_X1 i_0_0_24 (.A1(n_0_118), .A2(Res_imm[47]), .ZN(n_0_70));
   AND2_X1 i_0_0_25 (.A1(n_0_118), .A2(A[0]), .ZN(n_0_71));
   AND2_X1 i_0_0_26 (.A1(n_0_118), .A2(A[1]), .ZN(n_0_72));
   AND2_X1 i_0_0_27 (.A1(n_0_118), .A2(A[2]), .ZN(n_0_73));
   AND2_X1 i_0_0_28 (.A1(n_0_118), .A2(A[3]), .ZN(n_0_74));
   AND2_X1 i_0_0_29 (.A1(n_0_118), .A2(A[4]), .ZN(n_0_75));
   AND2_X1 i_0_0_30 (.A1(n_0_118), .A2(A[5]), .ZN(n_0_76));
   AND2_X1 i_0_0_31 (.A1(n_0_118), .A2(A[6]), .ZN(n_0_77));
   AND2_X1 i_0_0_32 (.A1(n_0_118), .A2(A[7]), .ZN(n_0_78));
   AND2_X1 i_0_0_33 (.A1(n_0_118), .A2(A[8]), .ZN(n_0_79));
   AND2_X1 i_0_0_34 (.A1(n_0_118), .A2(A[9]), .ZN(n_0_80));
   AND2_X1 i_0_0_35 (.A1(n_0_118), .A2(A[10]), .ZN(n_0_81));
   AND2_X1 i_0_0_36 (.A1(n_0_118), .A2(A[11]), .ZN(n_0_82));
   AND2_X1 i_0_0_37 (.A1(n_0_118), .A2(A[12]), .ZN(n_0_83));
   AND2_X1 i_0_0_38 (.A1(n_0_118), .A2(A[13]), .ZN(n_0_84));
   AND2_X1 i_0_0_39 (.A1(n_0_118), .A2(A[14]), .ZN(n_0_85));
   AND2_X1 i_0_0_40 (.A1(n_0_118), .A2(A[15]), .ZN(n_0_86));
   AND2_X1 i_0_0_41 (.A1(n_0_118), .A2(A[16]), .ZN(n_0_87));
   AND2_X1 i_0_0_42 (.A1(n_0_118), .A2(A[17]), .ZN(n_0_88));
   AND2_X1 i_0_0_43 (.A1(n_0_118), .A2(A[18]), .ZN(n_0_89));
   AND2_X1 i_0_0_44 (.A1(n_0_118), .A2(A[19]), .ZN(n_0_90));
   AND2_X1 i_0_0_45 (.A1(n_0_118), .A2(A[20]), .ZN(n_0_91));
   AND2_X1 i_0_0_46 (.A1(n_0_118), .A2(A[21]), .ZN(n_0_92));
   AND2_X1 i_0_0_47 (.A1(n_0_118), .A2(A[22]), .ZN(n_0_93));
   INV_X1 i_0_0_48 (.A(n_0_0_0), .ZN(n_0_94));
   AOI21_X1 i_0_0_49 (.A(reset), .B1(clk), .B2(enable), .ZN(n_0_0_0));
   AND2_X1 i_0_0_50 (.A1(n_0_118), .A2(B[0]), .ZN(n_0_95));
   AND2_X1 i_0_0_51 (.A1(n_0_118), .A2(B[1]), .ZN(n_0_96));
   AND2_X1 i_0_0_52 (.A1(n_0_118), .A2(B[2]), .ZN(n_0_97));
   AND2_X1 i_0_0_53 (.A1(n_0_118), .A2(B[3]), .ZN(n_0_98));
   AND2_X1 i_0_0_54 (.A1(n_0_118), .A2(B[4]), .ZN(n_0_99));
   AND2_X1 i_0_0_55 (.A1(n_0_118), .A2(B[5]), .ZN(n_0_100));
   AND2_X1 i_0_0_56 (.A1(n_0_118), .A2(B[6]), .ZN(n_0_101));
   AND2_X1 i_0_0_57 (.A1(n_0_118), .A2(B[7]), .ZN(n_0_102));
   AND2_X1 i_0_0_58 (.A1(n_0_118), .A2(B[8]), .ZN(n_0_103));
   AND2_X1 i_0_0_59 (.A1(n_0_118), .A2(B[9]), .ZN(n_0_104));
   AND2_X1 i_0_0_60 (.A1(n_0_118), .A2(B[10]), .ZN(n_0_105));
   AND2_X1 i_0_0_61 (.A1(n_0_118), .A2(B[11]), .ZN(n_0_106));
   AND2_X1 i_0_0_62 (.A1(n_0_118), .A2(B[12]), .ZN(n_0_107));
   AND2_X1 i_0_0_63 (.A1(n_0_118), .A2(B[13]), .ZN(n_0_108));
   AND2_X1 i_0_0_64 (.A1(n_0_118), .A2(B[14]), .ZN(n_0_109));
   AND2_X1 i_0_0_65 (.A1(n_0_118), .A2(B[15]), .ZN(n_0_110));
   AND2_X1 i_0_0_66 (.A1(n_0_118), .A2(B[16]), .ZN(n_0_111));
   AND2_X1 i_0_0_67 (.A1(n_0_118), .A2(B[17]), .ZN(n_0_112));
   AND2_X1 i_0_0_68 (.A1(n_0_118), .A2(B[18]), .ZN(n_0_113));
   AND2_X1 i_0_0_69 (.A1(n_0_118), .A2(B[19]), .ZN(n_0_114));
   AND2_X1 i_0_0_70 (.A1(n_0_118), .A2(B[20]), .ZN(n_0_115));
   AND2_X1 i_0_0_71 (.A1(n_0_118), .A2(B[21]), .ZN(n_0_116));
   AND2_X1 i_0_0_72 (.A1(n_0_118), .A2(B[22]), .ZN(n_0_117));
   NAND2_X1 i_0_0_73 (.A1(n_0_118), .A2(clk), .ZN(n_0_119));
   INV_X1 i_0_0_74 (.A(reset), .ZN(n_0_118));
endmodule

module datapath__0_133(M_multiplied, p_0, M_resultTruncated);
   input M_multiplied;
   input [22:0]p_0;
   output [22:0]M_resultTruncated;

   HA_X1 i_0 (.A(M_multiplied), .B(p_0[0]), .CO(n_0), .S(M_resultTruncated[0]));
   HA_X1 i_1 (.A(p_0[1]), .B(n_0), .CO(n_1), .S(M_resultTruncated[1]));
   HA_X1 i_2 (.A(p_0[2]), .B(n_1), .CO(n_2), .S(M_resultTruncated[2]));
   HA_X1 i_3 (.A(p_0[3]), .B(n_2), .CO(n_3), .S(M_resultTruncated[3]));
   HA_X1 i_4 (.A(p_0[4]), .B(n_3), .CO(n_4), .S(M_resultTruncated[4]));
   HA_X1 i_5 (.A(p_0[5]), .B(n_4), .CO(n_5), .S(M_resultTruncated[5]));
   HA_X1 i_6 (.A(p_0[6]), .B(n_5), .CO(n_6), .S(M_resultTruncated[6]));
   HA_X1 i_7 (.A(p_0[7]), .B(n_6), .CO(n_7), .S(M_resultTruncated[7]));
   HA_X1 i_8 (.A(p_0[8]), .B(n_7), .CO(n_8), .S(M_resultTruncated[8]));
   HA_X1 i_9 (.A(p_0[9]), .B(n_8), .CO(n_9), .S(M_resultTruncated[9]));
   HA_X1 i_10 (.A(p_0[10]), .B(n_9), .CO(n_10), .S(M_resultTruncated[10]));
   HA_X1 i_11 (.A(p_0[11]), .B(n_10), .CO(n_11), .S(M_resultTruncated[11]));
   HA_X1 i_12 (.A(p_0[12]), .B(n_11), .CO(n_12), .S(M_resultTruncated[12]));
   HA_X1 i_13 (.A(p_0[13]), .B(n_12), .CO(n_13), .S(M_resultTruncated[13]));
   HA_X1 i_14 (.A(p_0[14]), .B(n_13), .CO(n_14), .S(M_resultTruncated[14]));
   HA_X1 i_15 (.A(p_0[15]), .B(n_14), .CO(n_15), .S(M_resultTruncated[15]));
   HA_X1 i_16 (.A(p_0[16]), .B(n_15), .CO(n_16), .S(M_resultTruncated[16]));
   HA_X1 i_17 (.A(p_0[17]), .B(n_16), .CO(n_17), .S(M_resultTruncated[17]));
   HA_X1 i_18 (.A(p_0[18]), .B(n_17), .CO(n_18), .S(M_resultTruncated[18]));
   HA_X1 i_19 (.A(p_0[19]), .B(n_18), .CO(n_19), .S(M_resultTruncated[19]));
   HA_X1 i_20 (.A(p_0[20]), .B(n_19), .CO(n_20), .S(M_resultTruncated[20]));
   HA_X1 i_21 (.A(p_0[21]), .B(n_20), .CO(n_21), .S(M_resultTruncated[21]));
   XOR2_X1 i_22 (.A(p_0[22]), .B(n_21), .Z(M_resultTruncated[22]));
endmodule

module FPU_multiplierTree(Res, A, B, clk, reset, enable);
   output [31:0]Res;
   input [31:0]A;
   input [31:0]B;
   input clk;
   input reset;
   input enable;

   wire [22:0]M_resultTruncated;
   wire [7:0]EA;
   wire [7:0]EB;
   wire A_reg;
   wire B_reg;
   wire n_0_1_2;
   wire n_0_1_3;
   wire n_0_1_4;
   wire n_0_1_5;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_1_8;
   wire n_0_1_9;
   wire n_0_1_10;
   wire n_0_1_11;
   wire n_0_1_12;
   wire n_0_1_13;
   wire n_0_1_14;
   wire n_0_1_15;
   wire n_0_1_22;
   wire n_0_1_16;
   wire n_0_1_23;
   wire n_0_1_17;
   wire n_0_1_24;
   wire n_0_1_18;
   wire n_0_1_25;
   wire n_0_1_19;
   wire n_0_1_26;
   wire n_0_1_20;
   wire n_0_1_27;
   wire n_0_1_21;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_1;
   wire n_0_1_32;
   wire n_0_2;
   wire n_0_1_33;
   wire n_0_3;
   wire n_0_1_34;
   wire n_0_4;
   wire n_0_1_35;
   wire n_0_5;
   wire n_0_1_36;
   wire n_0_6;
   wire n_0_1_37;
   wire n_0_7;
   wire n_0_1_38;
   wire n_0_8;
   wire n_0_1_39;
   wire n_0_9;
   wire n_0_1_40;
   wire n_0_10;
   wire n_0_1_41;
   wire n_0_11;
   wire n_0_1_42;
   wire n_0_12;
   wire n_0_1_43;
   wire n_0_13;
   wire n_0_1_44;
   wire n_0_14;
   wire n_0_1_45;
   wire n_0_15;
   wire n_0_1_46;
   wire n_0_16;
   wire n_0_1_47;
   wire n_0_17;
   wire n_0_1_48;
   wire n_0_18;
   wire n_0_1_49;
   wire n_0_19;
   wire n_0_1_50;
   wire n_0_20;
   wire n_0_1_51;
   wire n_0_21;
   wire n_0_1_52;
   wire n_0_22;
   wire n_0_1_53;
   wire n_0_1_54;
   wire n_0_1_55;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_1_56;
   wire n_0_1_57;
   wire n_0_1_58;
   wire n_0_1_59;
   wire n_0_1_60;
   wire n_0_1_62;
   wire n_0_1_64;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_1_105;
   wire n_0_1_106;
   wire n_0_1_107;
   wire n_0_1_108;
   wire n_0_1_109;
   wire n_0_1_110;
   wire n_0_1_111;
   wire n_0_1_112;
   wire n_0_1_28;
   wire n_0_1_29;
   wire n_0_0;
   wire n_0_1_30;
   wire n_0_1_31;
   wire n_0_1_61;
   wire n_0_1_63;
   wire n_0_1_65;
   wire n_0_1_66;
   wire n_0_1_67;
   wire n_0_1_68;
   wire n_0_1_69;
   wire n_0_1_70;
   wire n_0_1_71;
   wire n_0_1_72;
   wire n_0_1_73;
   wire n_0_1_74;
   wire n_0_1_75;
   wire n_0_1_76;
   wire n_0_1_77;
   wire n_0_1_78;
   wire n_0_1_79;
   wire n_0_1_80;
   wire n_0_1_81;
   wire n_0_1_82;
   wire n_0_1_83;
   wire n_0_1_84;
   wire n_0_1_85;
   wire n_0_1_86;
   wire n_0_1_87;
   wire n_0_1_88;
   wire n_0_1_89;
   wire n_0_1_90;
   wire n_0_1_91;
   wire n_0_1_92;
   wire n_0_1_93;
   wire n_0_1_94;
   wire n_0_1_95;
   wire n_0_1_96;
   wire n_0_1_97;
   wire n_0_1_98;
   wire n_0_1_99;
   wire n_0_1_100;
   wire n_0_1_101;
   wire n_0_1_102;
   wire n_0_1_103;
   wire n_0_31;
   wire n_0_1_104;

   multiplierTree multiplier (.Res({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, 
      uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, n_24, n_23, 
      n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, 
      n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, uc_16, uc_17, 
      uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, 
      uc_28, uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, 
      uc_38}), .OVF(), .A({uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, 
      uc_46, uc_47, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, 
      n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, 
      n_47}), .B({uc_48, uc_49, uc_50, uc_51, uc_52, uc_53, uc_54, uc_55, uc_56, 
      n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, 
      n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70}), 
      .clk(clk), .reset(reset), .enable(enable));
   datapath__0_133 i_0_0 (.M_multiplied(n_0), .p_0({n_23, n_22, n_21, n_20, n_19, 
      n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, 
      n_5, n_4, n_3, n_2, n_1}), .M_resultTruncated(M_resultTruncated));
   DLH_X1 \Res_reg[31]  (.D(n_0_31), .G(n_0_97), .Q(Res[31]));
   DLH_X1 \Res_reg[30]  (.D(n_0_30), .G(n_0_97), .Q(Res[30]));
   DLH_X1 \Res_reg[29]  (.D(n_0_29), .G(n_0_97), .Q(Res[29]));
   DLH_X1 \Res_reg[28]  (.D(n_0_28), .G(n_0_97), .Q(Res[28]));
   DLH_X1 \Res_reg[27]  (.D(n_0_27), .G(n_0_97), .Q(Res[27]));
   DLH_X1 \Res_reg[26]  (.D(n_0_26), .G(n_0_97), .Q(Res[26]));
   DLH_X1 \Res_reg[25]  (.D(n_0_25), .G(n_0_97), .Q(Res[25]));
   DLH_X1 \Res_reg[24]  (.D(n_0_24), .G(n_0_97), .Q(Res[24]));
   DLH_X1 \Res_reg[23]  (.D(n_0_23), .G(n_0_97), .Q(Res[23]));
   DLH_X1 \Res_reg[22]  (.D(n_0_22), .G(n_0_97), .Q(Res[22]));
   DLH_X1 \Res_reg[21]  (.D(n_0_21), .G(n_0_97), .Q(Res[21]));
   DLH_X1 \Res_reg[20]  (.D(n_0_20), .G(n_0_97), .Q(Res[20]));
   DLH_X1 \Res_reg[19]  (.D(n_0_19), .G(n_0_97), .Q(Res[19]));
   DLH_X1 \Res_reg[18]  (.D(n_0_18), .G(n_0_97), .Q(Res[18]));
   DLH_X1 \Res_reg[17]  (.D(n_0_17), .G(n_0_97), .Q(Res[17]));
   DLH_X1 \Res_reg[16]  (.D(n_0_16), .G(n_0_97), .Q(Res[16]));
   DLH_X1 \Res_reg[15]  (.D(n_0_15), .G(n_0_97), .Q(Res[15]));
   DLH_X1 \Res_reg[14]  (.D(n_0_14), .G(n_0_97), .Q(Res[14]));
   DLH_X1 \Res_reg[13]  (.D(n_0_13), .G(n_0_97), .Q(Res[13]));
   DLH_X1 \Res_reg[12]  (.D(n_0_12), .G(n_0_97), .Q(Res[12]));
   DLH_X1 \Res_reg[11]  (.D(n_0_11), .G(n_0_97), .Q(Res[11]));
   DLH_X1 \Res_reg[10]  (.D(n_0_10), .G(n_0_97), .Q(Res[10]));
   DLH_X1 \Res_reg[9]  (.D(n_0_9), .G(n_0_97), .Q(Res[9]));
   DLH_X1 \Res_reg[8]  (.D(n_0_8), .G(n_0_97), .Q(Res[8]));
   DLH_X1 \Res_reg[7]  (.D(n_0_7), .G(n_0_97), .Q(Res[7]));
   DLH_X1 \Res_reg[6]  (.D(n_0_6), .G(n_0_97), .Q(Res[6]));
   DLH_X1 \Res_reg[5]  (.D(n_0_5), .G(n_0_97), .Q(Res[5]));
   DLH_X1 \Res_reg[4]  (.D(n_0_4), .G(n_0_97), .Q(Res[4]));
   DLH_X1 \Res_reg[3]  (.D(n_0_3), .G(n_0_97), .Q(Res[3]));
   DLH_X1 \Res_reg[2]  (.D(n_0_2), .G(n_0_97), .Q(Res[2]));
   DLH_X1 \Res_reg[1]  (.D(n_0_1), .G(n_0_97), .Q(Res[1]));
   DLH_X1 \Res_reg[0]  (.D(n_0_0), .G(n_0_97), .Q(Res[0]));
   DLH_X1 \A_reg_reg[30]  (.D(n_0_65), .G(n_0_33), .Q(EA[7]));
   DLH_X1 \A_reg_reg[29]  (.D(n_0_64), .G(n_0_33), .Q(EA[6]));
   DLH_X1 \A_reg_reg[28]  (.D(n_0_63), .G(n_0_33), .Q(EA[5]));
   DLH_X1 \A_reg_reg[27]  (.D(n_0_62), .G(n_0_33), .Q(EA[4]));
   DLH_X1 \A_reg_reg[26]  (.D(n_0_61), .G(n_0_33), .Q(EA[3]));
   DLH_X1 \A_reg_reg[25]  (.D(n_0_60), .G(n_0_33), .Q(EA[2]));
   DLH_X1 \A_reg_reg[24]  (.D(n_0_59), .G(n_0_33), .Q(EA[1]));
   DLH_X1 \A_reg_reg[23]  (.D(n_0_58), .G(n_0_33), .Q(EA[0]));
   DLH_X1 \A_reg_reg[22]  (.D(n_0_57), .G(n_0_33), .Q(n_25));
   DLH_X1 \A_reg_reg[21]  (.D(n_0_56), .G(n_0_33), .Q(n_26));
   DLH_X1 \A_reg_reg[20]  (.D(n_0_55), .G(n_0_33), .Q(n_27));
   DLH_X1 \A_reg_reg[19]  (.D(n_0_54), .G(n_0_33), .Q(n_28));
   DLH_X1 \A_reg_reg[18]  (.D(n_0_53), .G(n_0_33), .Q(n_29));
   DLH_X1 \A_reg_reg[17]  (.D(n_0_52), .G(n_0_33), .Q(n_30));
   DLH_X1 \A_reg_reg[16]  (.D(n_0_51), .G(n_0_33), .Q(n_31));
   DLH_X1 \A_reg_reg[15]  (.D(n_0_50), .G(n_0_33), .Q(n_32));
   DLH_X1 \A_reg_reg[14]  (.D(n_0_49), .G(n_0_33), .Q(n_33));
   DLH_X1 \A_reg_reg[13]  (.D(n_0_48), .G(n_0_33), .Q(n_34));
   DLH_X1 \A_reg_reg[12]  (.D(n_0_47), .G(n_0_33), .Q(n_35));
   DLH_X1 \A_reg_reg[11]  (.D(n_0_46), .G(n_0_33), .Q(n_36));
   DLH_X1 \A_reg_reg[10]  (.D(n_0_45), .G(n_0_33), .Q(n_37));
   DLH_X1 \A_reg_reg[9]  (.D(n_0_44), .G(n_0_33), .Q(n_38));
   DLH_X1 \A_reg_reg[8]  (.D(n_0_43), .G(n_0_33), .Q(n_39));
   DLH_X1 \A_reg_reg[7]  (.D(n_0_42), .G(n_0_33), .Q(n_40));
   DLH_X1 \A_reg_reg[6]  (.D(n_0_41), .G(n_0_33), .Q(n_41));
   DLH_X1 \A_reg_reg[5]  (.D(n_0_40), .G(n_0_33), .Q(n_42));
   DLH_X1 \A_reg_reg[4]  (.D(n_0_39), .G(n_0_33), .Q(n_43));
   DLH_X1 \A_reg_reg[3]  (.D(n_0_38), .G(n_0_33), .Q(n_44));
   DLH_X1 \A_reg_reg[2]  (.D(n_0_37), .G(n_0_33), .Q(n_45));
   DLH_X1 \A_reg_reg[1]  (.D(n_0_36), .G(n_0_33), .Q(n_46));
   DLH_X1 \A_reg_reg[0]  (.D(n_0_35), .G(n_0_33), .Q(n_47));
   DLH_X1 \B_reg_reg[30]  (.D(n_0_96), .G(n_0_33), .Q(EB[7]));
   DLH_X1 \B_reg_reg[29]  (.D(n_0_95), .G(n_0_33), .Q(EB[6]));
   DLH_X1 \B_reg_reg[28]  (.D(n_0_94), .G(n_0_33), .Q(EB[5]));
   DLH_X1 \B_reg_reg[27]  (.D(n_0_93), .G(n_0_33), .Q(EB[4]));
   DLH_X1 \B_reg_reg[26]  (.D(n_0_92), .G(n_0_33), .Q(EB[3]));
   DLH_X1 \B_reg_reg[25]  (.D(n_0_91), .G(n_0_33), .Q(EB[2]));
   DLH_X1 \B_reg_reg[24]  (.D(n_0_90), .G(n_0_33), .Q(EB[1]));
   DLH_X1 \B_reg_reg[23]  (.D(n_0_89), .G(n_0_33), .Q(EB[0]));
   DLH_X1 \B_reg_reg[22]  (.D(n_0_88), .G(n_0_33), .Q(n_48));
   DLH_X1 \B_reg_reg[21]  (.D(n_0_87), .G(n_0_33), .Q(n_49));
   DLH_X1 \B_reg_reg[20]  (.D(n_0_86), .G(n_0_33), .Q(n_50));
   DLH_X1 \B_reg_reg[19]  (.D(n_0_85), .G(n_0_33), .Q(n_51));
   DLH_X1 \B_reg_reg[18]  (.D(n_0_84), .G(n_0_33), .Q(n_52));
   DLH_X1 \B_reg_reg[17]  (.D(n_0_83), .G(n_0_33), .Q(n_53));
   DLH_X1 \B_reg_reg[16]  (.D(n_0_82), .G(n_0_33), .Q(n_54));
   DLH_X1 \B_reg_reg[15]  (.D(n_0_81), .G(n_0_33), .Q(n_55));
   DLH_X1 \B_reg_reg[14]  (.D(n_0_80), .G(n_0_33), .Q(n_56));
   DLH_X1 \B_reg_reg[13]  (.D(n_0_79), .G(n_0_33), .Q(n_57));
   DLH_X1 \B_reg_reg[12]  (.D(n_0_78), .G(n_0_33), .Q(n_58));
   DLH_X1 \B_reg_reg[11]  (.D(n_0_77), .G(n_0_33), .Q(n_59));
   DLH_X1 \B_reg_reg[10]  (.D(n_0_76), .G(n_0_33), .Q(n_60));
   DLH_X1 \B_reg_reg[9]  (.D(n_0_75), .G(n_0_33), .Q(n_61));
   DLH_X1 \B_reg_reg[8]  (.D(n_0_74), .G(n_0_33), .Q(n_62));
   DLH_X1 \B_reg_reg[7]  (.D(n_0_73), .G(n_0_33), .Q(n_63));
   DLH_X1 \B_reg_reg[6]  (.D(n_0_72), .G(n_0_33), .Q(n_64));
   DLH_X1 \B_reg_reg[5]  (.D(n_0_71), .G(n_0_33), .Q(n_65));
   DLH_X1 \B_reg_reg[4]  (.D(n_0_70), .G(n_0_33), .Q(n_66));
   DLH_X1 \B_reg_reg[3]  (.D(n_0_69), .G(n_0_33), .Q(n_67));
   DLH_X1 \B_reg_reg[2]  (.D(n_0_68), .G(n_0_33), .Q(n_68));
   DLH_X1 \B_reg_reg[1]  (.D(n_0_67), .G(n_0_33), .Q(n_69));
   DLH_X1 \B_reg_reg[0]  (.D(n_0_66), .G(n_0_33), .Q(n_70));
   DLH_X1 \A_reg_reg[31]  (.D(n_0_32), .G(n_0_33), .Q(A_reg));
   DLH_X1 \B_reg_reg[31]  (.D(n_0_34), .G(n_0_33), .Q(B_reg));
   HA_X1 i_0_1_0 (.A(EB[1]), .B(EA[1]), .CO(n_0_1_3), .S(n_0_1_2));
   HA_X1 i_0_1_1 (.A(EB[2]), .B(EA[2]), .CO(n_0_1_5), .S(n_0_1_4));
   HA_X1 i_0_1_2 (.A(EB[3]), .B(EA[3]), .CO(n_0_1_7), .S(n_0_1_6));
   HA_X1 i_0_1_3 (.A(EB[4]), .B(EA[4]), .CO(n_0_1_9), .S(n_0_1_8));
   HA_X1 i_0_1_4 (.A(EB[5]), .B(EA[5]), .CO(n_0_1_11), .S(n_0_1_10));
   HA_X1 i_0_1_5 (.A(EB[6]), .B(EA[6]), .CO(n_0_1_13), .S(n_0_1_12));
   HA_X1 i_0_1_6 (.A(EA[0]), .B(n_0_1_0), .CO(n_0_1_15), .S(n_0_1_14));
   FA_X1 i_0_1_7 (.A(n_0_1_1), .B(n_0_1_2), .CI(n_0_1_15), .CO(n_0_1_16), 
      .S(n_0_1_22));
   FA_X1 i_0_1_8 (.A(n_0_1_3), .B(n_0_1_4), .CI(n_0_1_16), .CO(n_0_1_17), 
      .S(n_0_1_23));
   FA_X1 i_0_1_9 (.A(n_0_1_5), .B(n_0_1_6), .CI(n_0_1_17), .CO(n_0_1_18), 
      .S(n_0_1_24));
   FA_X1 i_0_1_10 (.A(n_0_1_7), .B(n_0_1_8), .CI(n_0_1_18), .CO(n_0_1_19), 
      .S(n_0_1_25));
   FA_X1 i_0_1_11 (.A(n_0_1_9), .B(n_0_1_10), .CI(n_0_1_19), .CO(n_0_1_20), 
      .S(n_0_1_26));
   FA_X1 i_0_1_12 (.A(n_0_1_11), .B(n_0_1_12), .CI(n_0_1_20), .CO(n_0_1_21), 
      .S(n_0_1_27));
   XNOR2_X1 i_0_1_13 (.A(EB[0]), .B(n_24), .ZN(n_0_1_0));
   OR2_X1 i_0_1_14 (.A1(EB[0]), .A2(n_24), .ZN(n_0_1_1));
   INV_X1 i_0_1_15 (.A(n_0_1_32), .ZN(n_0_1));
   AOI22_X1 i_0_1_16 (.A1(M_resultTruncated[1]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_1), .ZN(n_0_1_32));
   INV_X1 i_0_1_22 (.A(n_0_1_33), .ZN(n_0_2));
   AOI22_X1 i_0_1_23 (.A1(M_resultTruncated[2]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_2), .ZN(n_0_1_33));
   INV_X1 i_0_1_24 (.A(n_0_1_34), .ZN(n_0_3));
   AOI22_X1 i_0_1_25 (.A1(M_resultTruncated[3]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_3), .ZN(n_0_1_34));
   INV_X1 i_0_1_26 (.A(n_0_1_35), .ZN(n_0_4));
   AOI22_X1 i_0_1_27 (.A1(M_resultTruncated[4]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_4), .ZN(n_0_1_35));
   INV_X1 i_0_1_28 (.A(n_0_1_36), .ZN(n_0_5));
   AOI22_X1 i_0_1_29 (.A1(M_resultTruncated[5]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_5), .ZN(n_0_1_36));
   INV_X1 i_0_1_30 (.A(n_0_1_37), .ZN(n_0_6));
   AOI22_X1 i_0_1_31 (.A1(M_resultTruncated[6]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_6), .ZN(n_0_1_37));
   INV_X1 i_0_1_32 (.A(n_0_1_38), .ZN(n_0_7));
   AOI22_X1 i_0_1_33 (.A1(M_resultTruncated[7]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_7), .ZN(n_0_1_38));
   INV_X1 i_0_1_34 (.A(n_0_1_39), .ZN(n_0_8));
   AOI22_X1 i_0_1_35 (.A1(M_resultTruncated[8]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_8), .ZN(n_0_1_39));
   INV_X1 i_0_1_36 (.A(n_0_1_40), .ZN(n_0_9));
   AOI22_X1 i_0_1_37 (.A1(M_resultTruncated[9]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_9), .ZN(n_0_1_40));
   INV_X1 i_0_1_38 (.A(n_0_1_41), .ZN(n_0_10));
   AOI22_X1 i_0_1_39 (.A1(M_resultTruncated[10]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_10), .ZN(n_0_1_41));
   INV_X1 i_0_1_40 (.A(n_0_1_42), .ZN(n_0_11));
   AOI22_X1 i_0_1_41 (.A1(M_resultTruncated[11]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_11), .ZN(n_0_1_42));
   INV_X1 i_0_1_42 (.A(n_0_1_43), .ZN(n_0_12));
   AOI22_X1 i_0_1_43 (.A1(M_resultTruncated[12]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_12), .ZN(n_0_1_43));
   INV_X1 i_0_1_44 (.A(n_0_1_44), .ZN(n_0_13));
   AOI22_X1 i_0_1_45 (.A1(M_resultTruncated[13]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_13), .ZN(n_0_1_44));
   INV_X1 i_0_1_46 (.A(n_0_1_45), .ZN(n_0_14));
   AOI22_X1 i_0_1_47 (.A1(M_resultTruncated[14]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_14), .ZN(n_0_1_45));
   INV_X1 i_0_1_48 (.A(n_0_1_46), .ZN(n_0_15));
   AOI22_X1 i_0_1_49 (.A1(M_resultTruncated[15]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_15), .ZN(n_0_1_46));
   INV_X1 i_0_1_50 (.A(n_0_1_47), .ZN(n_0_16));
   AOI22_X1 i_0_1_51 (.A1(M_resultTruncated[16]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_16), .ZN(n_0_1_47));
   INV_X1 i_0_1_52 (.A(n_0_1_48), .ZN(n_0_17));
   AOI22_X1 i_0_1_53 (.A1(M_resultTruncated[17]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_17), .ZN(n_0_1_48));
   INV_X1 i_0_1_54 (.A(n_0_1_49), .ZN(n_0_18));
   AOI22_X1 i_0_1_55 (.A1(M_resultTruncated[18]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_18), .ZN(n_0_1_49));
   INV_X1 i_0_1_56 (.A(n_0_1_50), .ZN(n_0_19));
   AOI22_X1 i_0_1_57 (.A1(M_resultTruncated[19]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_19), .ZN(n_0_1_50));
   INV_X1 i_0_1_58 (.A(n_0_1_51), .ZN(n_0_20));
   AOI22_X1 i_0_1_59 (.A1(M_resultTruncated[20]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_20), .ZN(n_0_1_51));
   INV_X1 i_0_1_60 (.A(n_0_1_52), .ZN(n_0_21));
   AOI22_X1 i_0_1_61 (.A1(M_resultTruncated[21]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_21), .ZN(n_0_1_52));
   INV_X1 i_0_1_62 (.A(n_0_1_53), .ZN(n_0_22));
   AOI22_X1 i_0_1_63 (.A1(M_resultTruncated[22]), .A2(n_0_1_55), .B1(n_0_1_54), 
      .B2(n_22), .ZN(n_0_1_53));
   NOR3_X1 i_0_1_17 (.A1(n_0_1_60), .A2(n_24), .A3(n_0_1_64), .ZN(n_0_1_54));
   NOR3_X1 i_0_1_18 (.A1(n_0_1_29), .A2(n_0_1_64), .A3(n_0_1_60), .ZN(n_0_1_55));
   OAI21_X1 i_0_1_19 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_111), .ZN(n_0_23));
   OAI21_X1 i_0_1_67 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_110), .ZN(n_0_24));
   OAI21_X1 i_0_1_68 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_109), .ZN(n_0_25));
   OAI21_X1 i_0_1_69 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_108), .ZN(n_0_26));
   OAI21_X1 i_0_1_70 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_107), .ZN(n_0_27));
   OAI21_X1 i_0_1_71 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_106), .ZN(n_0_28));
   OAI21_X1 i_0_1_72 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_105), .ZN(n_0_29));
   OAI21_X1 i_0_1_73 (.A(n_0_1_62), .B1(n_0_1_60), .B2(n_0_1_56), .ZN(n_0_30));
   XNOR2_X1 i_0_1_74 (.A(n_0_1_58), .B(n_0_1_57), .ZN(n_0_1_56));
   XNOR2_X1 i_0_1_75 (.A(n_0_1_13), .B(n_0_1_21), .ZN(n_0_1_57));
   NOR2_X1 i_0_1_76 (.A1(n_0_1_68), .A2(n_0_1_59), .ZN(n_0_1_58));
   NOR2_X1 i_0_1_77 (.A1(EB[7]), .A2(EA[7]), .ZN(n_0_1_59));
   NAND2_X1 i_0_1_20 (.A1(n_0_1_69), .A2(n_0_1_66), .ZN(n_0_1_60));
   AOI21_X1 i_0_1_21 (.A(n_0_1_72), .B1(n_0_1_69), .B2(n_0_1_64), .ZN(n_0_1_62));
   NAND3_X1 i_0_1_64 (.A1(n_0_1_100), .A2(n_0_1_97), .A3(n_0_1_67), .ZN(n_0_1_64));
   AND2_X1 i_0_1_65 (.A1(n_0_1_112), .A2(A[31]), .ZN(n_0_32));
   OAI21_X1 i_0_1_125 (.A(n_0_1_112), .B1(n_0_1_28), .B2(clk), .ZN(n_0_33));
   AND2_X1 i_0_1_126 (.A1(n_0_1_112), .A2(B[31]), .ZN(n_0_34));
   AND2_X1 i_0_1_127 (.A1(n_0_1_112), .A2(A[0]), .ZN(n_0_35));
   AND2_X1 i_0_1_128 (.A1(n_0_1_112), .A2(A[1]), .ZN(n_0_36));
   AND2_X1 i_0_1_129 (.A1(n_0_1_112), .A2(A[2]), .ZN(n_0_37));
   AND2_X1 i_0_1_130 (.A1(n_0_1_112), .A2(A[3]), .ZN(n_0_38));
   AND2_X1 i_0_1_131 (.A1(n_0_1_112), .A2(A[4]), .ZN(n_0_39));
   AND2_X1 i_0_1_132 (.A1(n_0_1_112), .A2(A[5]), .ZN(n_0_40));
   AND2_X1 i_0_1_133 (.A1(n_0_1_112), .A2(A[6]), .ZN(n_0_41));
   AND2_X1 i_0_1_134 (.A1(n_0_1_112), .A2(A[7]), .ZN(n_0_42));
   AND2_X1 i_0_1_135 (.A1(n_0_1_112), .A2(A[8]), .ZN(n_0_43));
   AND2_X1 i_0_1_136 (.A1(n_0_1_112), .A2(A[9]), .ZN(n_0_44));
   AND2_X1 i_0_1_137 (.A1(n_0_1_112), .A2(A[10]), .ZN(n_0_45));
   AND2_X1 i_0_1_138 (.A1(n_0_1_112), .A2(A[11]), .ZN(n_0_46));
   AND2_X1 i_0_1_139 (.A1(n_0_1_112), .A2(A[12]), .ZN(n_0_47));
   AND2_X1 i_0_1_140 (.A1(n_0_1_112), .A2(A[13]), .ZN(n_0_48));
   AND2_X1 i_0_1_141 (.A1(n_0_1_112), .A2(A[14]), .ZN(n_0_49));
   AND2_X1 i_0_1_142 (.A1(n_0_1_112), .A2(A[15]), .ZN(n_0_50));
   AND2_X1 i_0_1_143 (.A1(n_0_1_112), .A2(A[16]), .ZN(n_0_51));
   AND2_X1 i_0_1_144 (.A1(n_0_1_112), .A2(A[17]), .ZN(n_0_52));
   AND2_X1 i_0_1_145 (.A1(n_0_1_112), .A2(A[18]), .ZN(n_0_53));
   AND2_X1 i_0_1_146 (.A1(n_0_1_112), .A2(A[19]), .ZN(n_0_54));
   AND2_X1 i_0_1_147 (.A1(n_0_1_112), .A2(A[20]), .ZN(n_0_55));
   AND2_X1 i_0_1_148 (.A1(n_0_1_112), .A2(A[21]), .ZN(n_0_56));
   AND2_X1 i_0_1_149 (.A1(n_0_1_112), .A2(A[22]), .ZN(n_0_57));
   AND2_X1 i_0_1_150 (.A1(n_0_1_112), .A2(A[23]), .ZN(n_0_58));
   AND2_X1 i_0_1_151 (.A1(n_0_1_112), .A2(A[24]), .ZN(n_0_59));
   AND2_X1 i_0_1_152 (.A1(n_0_1_112), .A2(A[25]), .ZN(n_0_60));
   AND2_X1 i_0_1_153 (.A1(n_0_1_112), .A2(A[26]), .ZN(n_0_61));
   AND2_X1 i_0_1_154 (.A1(n_0_1_112), .A2(A[27]), .ZN(n_0_62));
   AND2_X1 i_0_1_155 (.A1(n_0_1_112), .A2(A[28]), .ZN(n_0_63));
   AND2_X1 i_0_1_156 (.A1(n_0_1_112), .A2(A[29]), .ZN(n_0_64));
   AND2_X1 i_0_1_157 (.A1(n_0_1_112), .A2(A[30]), .ZN(n_0_65));
   AND2_X1 i_0_1_158 (.A1(n_0_1_112), .A2(B[0]), .ZN(n_0_66));
   AND2_X1 i_0_1_159 (.A1(n_0_1_112), .A2(B[1]), .ZN(n_0_67));
   AND2_X1 i_0_1_160 (.A1(n_0_1_112), .A2(B[2]), .ZN(n_0_68));
   AND2_X1 i_0_1_161 (.A1(n_0_1_112), .A2(B[3]), .ZN(n_0_69));
   AND2_X1 i_0_1_162 (.A1(n_0_1_112), .A2(B[4]), .ZN(n_0_70));
   AND2_X1 i_0_1_163 (.A1(n_0_1_112), .A2(B[5]), .ZN(n_0_71));
   AND2_X1 i_0_1_164 (.A1(n_0_1_112), .A2(B[6]), .ZN(n_0_72));
   AND2_X1 i_0_1_165 (.A1(n_0_1_112), .A2(B[7]), .ZN(n_0_73));
   AND2_X1 i_0_1_166 (.A1(n_0_1_112), .A2(B[8]), .ZN(n_0_74));
   AND2_X1 i_0_1_167 (.A1(n_0_1_112), .A2(B[9]), .ZN(n_0_75));
   AND2_X1 i_0_1_168 (.A1(n_0_1_112), .A2(B[10]), .ZN(n_0_76));
   AND2_X1 i_0_1_169 (.A1(n_0_1_112), .A2(B[11]), .ZN(n_0_77));
   AND2_X1 i_0_1_170 (.A1(n_0_1_112), .A2(B[12]), .ZN(n_0_78));
   AND2_X1 i_0_1_171 (.A1(n_0_1_112), .A2(B[13]), .ZN(n_0_79));
   AND2_X1 i_0_1_172 (.A1(n_0_1_112), .A2(B[14]), .ZN(n_0_80));
   AND2_X1 i_0_1_173 (.A1(n_0_1_112), .A2(B[15]), .ZN(n_0_81));
   AND2_X1 i_0_1_174 (.A1(n_0_1_112), .A2(B[16]), .ZN(n_0_82));
   AND2_X1 i_0_1_175 (.A1(n_0_1_112), .A2(B[17]), .ZN(n_0_83));
   AND2_X1 i_0_1_176 (.A1(n_0_1_112), .A2(B[18]), .ZN(n_0_84));
   AND2_X1 i_0_1_177 (.A1(n_0_1_112), .A2(B[19]), .ZN(n_0_85));
   AND2_X1 i_0_1_178 (.A1(n_0_1_112), .A2(B[20]), .ZN(n_0_86));
   AND2_X1 i_0_1_179 (.A1(n_0_1_112), .A2(B[21]), .ZN(n_0_87));
   AND2_X1 i_0_1_180 (.A1(n_0_1_112), .A2(B[22]), .ZN(n_0_88));
   AND2_X1 i_0_1_181 (.A1(n_0_1_112), .A2(B[23]), .ZN(n_0_89));
   AND2_X1 i_0_1_182 (.A1(n_0_1_112), .A2(B[24]), .ZN(n_0_90));
   AND2_X1 i_0_1_183 (.A1(n_0_1_112), .A2(B[25]), .ZN(n_0_91));
   AND2_X1 i_0_1_184 (.A1(n_0_1_112), .A2(B[26]), .ZN(n_0_92));
   AND2_X1 i_0_1_185 (.A1(n_0_1_112), .A2(B[27]), .ZN(n_0_93));
   AND2_X1 i_0_1_186 (.A1(n_0_1_112), .A2(B[28]), .ZN(n_0_94));
   AND2_X1 i_0_1_187 (.A1(n_0_1_112), .A2(B[29]), .ZN(n_0_95));
   AND2_X1 i_0_1_188 (.A1(n_0_1_112), .A2(B[30]), .ZN(n_0_96));
   OR2_X1 i_0_1_189 (.A1(clk), .A2(reset), .ZN(n_0_97));
   INV_X1 i_0_1_190 (.A(n_0_1_27), .ZN(n_0_1_105));
   INV_X1 i_0_1_191 (.A(n_0_1_26), .ZN(n_0_1_106));
   INV_X1 i_0_1_192 (.A(n_0_1_25), .ZN(n_0_1_107));
   INV_X1 i_0_1_193 (.A(n_0_1_24), .ZN(n_0_1_108));
   INV_X1 i_0_1_194 (.A(n_0_1_23), .ZN(n_0_1_109));
   INV_X1 i_0_1_195 (.A(n_0_1_22), .ZN(n_0_1_110));
   INV_X1 i_0_1_66 (.A(n_0_1_14), .ZN(n_0_1_111));
   INV_X1 i_0_1_78 (.A(reset), .ZN(n_0_1_112));
   INV_X1 i_0_1_198 (.A(enable), .ZN(n_0_1_28));
   INV_X1 i_0_1_79 (.A(n_24), .ZN(n_0_1_29));
   OAI21_X1 i_0_1_80 (.A(n_0_1_71), .B1(n_0_1_31), .B2(n_0_1_30), .ZN(n_0_0));
   OAI221_X1 i_0_1_81 (.A(n_0_1_69), .B1(n_0_1_100), .B2(n_0_1_81), .C1(n_0_1_97), 
      .C2(n_0_1_73), .ZN(n_0_1_30));
   INV_X1 i_0_1_82 (.A(n_0_1_61), .ZN(n_0_1_31));
   OAI211_X1 i_0_1_83 (.A(n_0_1_100), .B(n_0_1_97), .C1(n_0_1_65), .C2(n_0_1_63), 
      .ZN(n_0_1_61));
   NAND2_X1 i_0_1_84 (.A1(n_0_1_67), .A2(n_0_1_66), .ZN(n_0_1_63));
   AOI22_X1 i_0_1_85 (.A1(n_0_1_103), .A2(n_0), .B1(n_24), .B2(
      M_resultTruncated[0]), .ZN(n_0_1_65));
   OR4_X1 i_0_1_86 (.A1(n_0_1_101), .A2(n_0_1_98), .A3(n_0_1_92), .A4(n_0_1_95), 
      .ZN(n_0_1_66));
   OAI221_X1 i_0_1_87 (.A(n_0_1_68), .B1(EA[6]), .B2(n_0_1_98), .C1(EB[6]), 
      .C2(n_0_1_101), .ZN(n_0_1_67));
   AND2_X1 i_0_1_88 (.A1(EA[7]), .A2(EB[7]), .ZN(n_0_1_68));
   NOR2_X1 i_0_1_89 (.A1(reset), .A2(n_0_1_70), .ZN(n_0_1_69));
   OAI22_X1 i_0_1_90 (.A1(n_0_1_91), .A2(n_0_1_81), .B1(n_0_1_94), .B2(n_0_1_73), 
      .ZN(n_0_1_70));
   INV_X1 i_0_1_91 (.A(n_0_1_72), .ZN(n_0_1_71));
   NOR4_X1 i_0_1_92 (.A1(reset), .A2(n_0_1_73), .A3(n_0_1_81), .A4(n_0_1_89), 
      .ZN(n_0_1_72));
   NAND3_X1 i_0_1_93 (.A1(n_0_1_78), .A2(n_0_1_77), .A3(n_0_1_74), .ZN(n_0_1_73));
   AND4_X1 i_0_1_94 (.A1(n_0_1_80), .A2(n_0_1_79), .A3(n_0_1_76), .A4(n_0_1_75), 
      .ZN(n_0_1_74));
   NOR4_X1 i_0_1_95 (.A1(n_45), .A2(n_47), .A3(n_41), .A4(n_44), .ZN(n_0_1_75));
   NOR4_X1 i_0_1_96 (.A1(n_37), .A2(n_40), .A3(n_34), .A4(n_35), .ZN(n_0_1_76));
   NOR3_X1 i_0_1_97 (.A1(n_42), .A2(n_43), .A3(n_46), .ZN(n_0_1_77));
   NOR4_X1 i_0_1_98 (.A1(n_38), .A2(n_39), .A3(n_33), .A4(n_36), .ZN(n_0_1_78));
   NOR4_X1 i_0_1_99 (.A1(n_25), .A2(n_26), .A3(n_27), .A4(n_28), .ZN(n_0_1_79));
   NOR4_X1 i_0_1_100 (.A1(n_29), .A2(n_30), .A3(n_31), .A4(n_32), .ZN(n_0_1_80));
   NAND3_X1 i_0_1_101 (.A1(n_0_1_86), .A2(n_0_1_85), .A3(n_0_1_82), .ZN(n_0_1_81));
   AND4_X1 i_0_1_102 (.A1(n_0_1_88), .A2(n_0_1_87), .A3(n_0_1_84), .A4(n_0_1_83), 
      .ZN(n_0_1_82));
   NOR4_X1 i_0_1_103 (.A1(n_68), .A2(n_70), .A3(n_64), .A4(n_67), .ZN(n_0_1_83));
   NOR4_X1 i_0_1_104 (.A1(n_60), .A2(n_63), .A3(n_57), .A4(n_58), .ZN(n_0_1_84));
   NOR3_X1 i_0_1_105 (.A1(n_65), .A2(n_66), .A3(n_69), .ZN(n_0_1_85));
   NOR4_X1 i_0_1_106 (.A1(n_61), .A2(n_62), .A3(n_56), .A4(n_59), .ZN(n_0_1_86));
   NOR4_X1 i_0_1_107 (.A1(n_48), .A2(n_49), .A3(n_50), .A4(n_51), .ZN(n_0_1_87));
   NOR4_X1 i_0_1_108 (.A1(n_52), .A2(n_53), .A3(n_54), .A4(n_55), .ZN(n_0_1_88));
   INV_X1 i_0_1_109 (.A(n_0_1_90), .ZN(n_0_1_89));
   OAI22_X1 i_0_1_110 (.A1(n_0_1_100), .A2(n_0_1_94), .B1(n_0_1_97), .B2(
      n_0_1_91), .ZN(n_0_1_90));
   OR4_X1 i_0_1_111 (.A1(n_0_1_93), .A2(n_0_1_92), .A3(EB[5]), .A4(EB[4]), 
      .ZN(n_0_1_91));
   OR2_X1 i_0_1_112 (.A1(EB[7]), .A2(EB[6]), .ZN(n_0_1_92));
   OR4_X1 i_0_1_113 (.A1(EB[3]), .A2(EB[2]), .A3(EB[1]), .A4(EB[0]), .ZN(
      n_0_1_93));
   OR4_X1 i_0_1_114 (.A1(n_0_1_96), .A2(n_0_1_95), .A3(EA[5]), .A4(EA[4]), 
      .ZN(n_0_1_94));
   OR2_X1 i_0_1_115 (.A1(EA[7]), .A2(EA[6]), .ZN(n_0_1_95));
   OR4_X1 i_0_1_116 (.A1(EA[3]), .A2(EA[2]), .A3(EA[1]), .A4(EA[0]), .ZN(
      n_0_1_96));
   NAND3_X1 i_0_1_117 (.A1(EA[7]), .A2(n_0_1_98), .A3(EA[6]), .ZN(n_0_1_97));
   AND3_X1 i_0_1_118 (.A1(EA[2]), .A2(EA[1]), .A3(n_0_1_99), .ZN(n_0_1_98));
   AND4_X1 i_0_1_119 (.A1(EA[5]), .A2(EA[4]), .A3(EA[3]), .A4(EA[0]), .ZN(
      n_0_1_99));
   NAND3_X1 i_0_1_120 (.A1(EB[7]), .A2(n_0_1_101), .A3(EB[6]), .ZN(n_0_1_100));
   AND3_X1 i_0_1_121 (.A1(EB[2]), .A2(EB[1]), .A3(n_0_1_102), .ZN(n_0_1_101));
   AND4_X1 i_0_1_122 (.A1(EB[5]), .A2(EB[4]), .A3(EB[3]), .A4(EB[0]), .ZN(
      n_0_1_102));
   INV_X1 i_0_1_123 (.A(n_24), .ZN(n_0_1_103));
   AOI211_X1 i_0_1_124 (.A(reset), .B(n_0_1_104), .C1(B_reg), .C2(A_reg), 
      .ZN(n_0_31));
   NOR2_X1 i_0_1_196 (.A1(B_reg), .A2(A_reg), .ZN(n_0_1_104));
endmodule
