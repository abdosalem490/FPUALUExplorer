
// 	Thu Dec 22 21:20:39 2022
//	vlsi
//	192.168.126.129

module datapath__0_13 (M_multiplied, p_0, M_resultTruncated);

output [22:0] M_resultTruncated;
input M_multiplied;
input [22:0] p_0;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;


XOR2_X1 i_22 (.Z (M_resultTruncated[22]), .A (p_0[22]), .B (n_21));
HA_X1 i_21 (.CO (n_21), .S (M_resultTruncated[21]), .A (p_0[21]), .B (n_20));
HA_X1 i_20 (.CO (n_20), .S (M_resultTruncated[20]), .A (p_0[20]), .B (n_19));
HA_X1 i_19 (.CO (n_19), .S (M_resultTruncated[19]), .A (p_0[19]), .B (n_18));
HA_X1 i_18 (.CO (n_18), .S (M_resultTruncated[18]), .A (p_0[18]), .B (n_17));
HA_X1 i_17 (.CO (n_17), .S (M_resultTruncated[17]), .A (p_0[17]), .B (n_16));
HA_X1 i_16 (.CO (n_16), .S (M_resultTruncated[16]), .A (p_0[16]), .B (n_15));
HA_X1 i_15 (.CO (n_15), .S (M_resultTruncated[15]), .A (p_0[15]), .B (n_14));
HA_X1 i_14 (.CO (n_14), .S (M_resultTruncated[14]), .A (p_0[14]), .B (n_13));
HA_X1 i_13 (.CO (n_13), .S (M_resultTruncated[13]), .A (p_0[13]), .B (n_12));
HA_X1 i_12 (.CO (n_12), .S (M_resultTruncated[12]), .A (p_0[12]), .B (n_11));
HA_X1 i_11 (.CO (n_11), .S (M_resultTruncated[11]), .A (p_0[11]), .B (n_10));
HA_X1 i_10 (.CO (n_10), .S (M_resultTruncated[10]), .A (p_0[10]), .B (n_9));
HA_X1 i_9 (.CO (n_9), .S (M_resultTruncated[9]), .A (p_0[9]), .B (n_8));
HA_X1 i_8 (.CO (n_8), .S (M_resultTruncated[8]), .A (p_0[8]), .B (n_7));
HA_X1 i_7 (.CO (n_7), .S (M_resultTruncated[7]), .A (p_0[7]), .B (n_6));
HA_X1 i_6 (.CO (n_6), .S (M_resultTruncated[6]), .A (p_0[6]), .B (n_5));
HA_X1 i_5 (.CO (n_5), .S (M_resultTruncated[5]), .A (p_0[5]), .B (n_4));
HA_X1 i_4 (.CO (n_4), .S (M_resultTruncated[4]), .A (p_0[4]), .B (n_3));
HA_X1 i_3 (.CO (n_3), .S (M_resultTruncated[3]), .A (p_0[3]), .B (n_2));
HA_X1 i_2 (.CO (n_2), .S (M_resultTruncated[2]), .A (p_0[2]), .B (n_1));
HA_X1 i_1 (.CO (n_1), .S (M_resultTruncated[1]), .A (p_0[1]), .B (n_0));
HA_X1 i_0 (.CO (n_0), .S (M_resultTruncated[0]), .A (M_multiplied), .B (p_0[0]));

endmodule //datapath__0_13

module datapath__0_2 (B_imm, A_imm, Res_imm);

output [63:0] Res_imm;
input [31:0] A_imm;
input [31:0] B_imm;
wire n_1538;
wire n_1723;
wire n_1;
wire n_0;
wire n_1514;
wire n_1537;
wire n_1560;
wire n_3;
wire n_2;
wire n_1581;
wire n_5;
wire n_4;
wire n_1559;
wire n_1580;
wire n_8;
wire n_6;
wire n_1466;
wire n_1489;
wire n_1512;
wire n_13;
wire n_9;
wire n_1535;
wire n_1558;
wire n_1579;
wire n_15;
wire n_10;
wire n_1442;
wire n_1465;
wire n_1488;
wire n_21;
wire n_12;
wire n_1511;
wire n_1534;
wire n_1557;
wire n_23;
wire n_14;
wire n_1578;
wire n_25;
wire n_20;
wire n_1418;
wire n_1441;
wire n_1464;
wire n_31;
wire n_22;
wire n_1487;
wire n_1510;
wire n_1533;
wire n_33;
wire n_24;
wire n_1556;
wire n_1577;
wire n_35;
wire n_34;
wire n_32;
wire n_30;
wire n_1394;
wire n_1417;
wire n_1440;
wire n_43;
wire n_42;
wire n_1463;
wire n_1486;
wire n_1509;
wire n_45;
wire n_44;
wire n_1532;
wire n_1555;
wire n_1576;
wire n_47;
wire n_46;
wire n_49;
wire n_36;
wire n_48;
wire n_37;
wire n_1370;
wire n_1393;
wire n_1416;
wire n_57;
wire n_56;
wire n_1439;
wire n_1462;
wire n_1485;
wire n_59;
wire n_58;
wire n_1508;
wire n_1531;
wire n_1554;
wire n_61;
wire n_60;
wire n_1575;
wire n_63;
wire n_62;
wire n_65;
wire n_50;
wire n_64;
wire n_51;
wire n_1346;
wire n_1369;
wire n_1392;
wire n_73;
wire n_72;
wire n_1415;
wire n_1438;
wire n_1461;
wire n_75;
wire n_74;
wire n_1484;
wire n_1507;
wire n_1530;
wire n_77;
wire n_76;
wire n_1553;
wire n_1574;
wire n_66;
wire n_78;
wire n_67;
wire n_80;
wire n_81;
wire n_79;
wire n_83;
wire n_82;
wire n_1322;
wire n_1345;
wire n_1368;
wire n_85;
wire n_84;
wire n_1391;
wire n_1414;
wire n_1437;
wire n_91;
wire n_90;
wire n_1460;
wire n_1483;
wire n_1506;
wire n_95;
wire n_92;
wire n_1529;
wire n_1552;
wire n_1573;
wire n_97;
wire n_93;
wire n_96;
wire n_94;
wire n_1298;
wire n_1321;
wire n_1344;
wire n_99;
wire n_98;
wire n_1367;
wire n_1390;
wire n_1413;
wire n_111;
wire n_110;
wire n_1436;
wire n_1459;
wire n_1482;
wire n_113;
wire n_112;
wire n_1505;
wire n_1528;
wire n_1551;
wire n_117;
wire n_114;
wire n_1572;
wire n_116;
wire n_115;
wire n_1274;
wire n_1297;
wire n_1320;
wire n_133;
wire n_118;
wire n_1343;
wire n_1366;
wire n_1389;
wire n_135;
wire n_119;
wire n_1412;
wire n_1435;
wire n_1458;
wire n_137;
wire n_132;
wire n_1481;
wire n_1504;
wire n_1527;
wire n_139;
wire n_134;
wire n_1550;
wire n_1571;
wire n_141;
wire n_136;
wire n_1250;
wire n_1273;
wire n_1296;
wire n_140;
wire n_138;
wire n_1319;
wire n_1342;
wire n_1365;
wire n_156;
wire n_143;
wire n_1388;
wire n_1411;
wire n_1434;
wire n_158;
wire n_157;
wire n_1457;
wire n_1480;
wire n_1503;
wire n_160;
wire n_159;
wire n_1526;
wire n_1549;
wire n_1570;
wire n_162;
wire n_161;
wire n_164;
wire n_163;
wire n_939;
wire n_166;
wire n_165;
wire n_1032;
wire n_1055;
wire n_1078;
wire n_551;
wire n_550;
wire n_1101;
wire n_1124;
wire n_1147;
wire n_553;
wire n_552;
wire n_1170;
wire n_1193;
wire n_1216;
wire n_555;
wire n_554;
wire n_1239;
wire n_1262;
wire n_1285;
wire n_557;
wire n_556;
wire n_1308;
wire n_1331;
wire n_1354;
wire n_559;
wire n_558;
wire n_1377;
wire n_1400;
wire n_1423;
wire n_561;
wire n_560;
wire n_1446;
wire n_1469;
wire n_1492;
wire n_563;
wire n_562;
wire n_1515;
wire n_800;
wire n_801;
wire n_565;
wire n_564;
wire n_788;
wire n_789;
wire n_790;
wire n_567;
wire n_566;
wire n_785;
wire n_786;
wire n_776;
wire n_569;
wire n_568;
wire n_778;
wire n_793;
wire n_571;
wire n_570;
wire n_573;
wire n_572;
wire n_575;
wire n_574;
wire n_829;
wire n_577;
wire n_576;
wire n_791;
wire n_828;
wire n_579;
wire n_578;
wire n_787;
wire n_780;
wire n_581;
wire n_580;
wire n_854;
wire n_583;
wire n_582;
wire n_792;
wire n_585;
wire n_584;
wire n_855;
wire n_783;
wire n_587;
wire n_586;
wire n_878;
wire n_589;
wire n_588;
wire n_879;
wire n_591;
wire n_590;
wire n_1031;
wire n_1054;
wire n_1077;
wire n_593;
wire n_592;
wire n_1100;
wire n_1123;
wire n_1146;
wire n_595;
wire n_594;
wire n_1169;
wire n_1192;
wire n_1215;
wire n_597;
wire n_596;
wire n_1238;
wire n_1261;
wire n_1284;
wire n_599;
wire n_598;
wire n_1307;
wire n_1330;
wire n_1353;
wire n_601;
wire n_600;
wire n_1376;
wire n_1399;
wire n_1422;
wire n_603;
wire n_602;
wire n_1445;
wire n_1468;
wire n_1491;
wire n_605;
wire n_604;
wire n_607;
wire n_606;
wire n_609;
wire n_608;
wire n_611;
wire n_610;
wire n_613;
wire n_612;
wire n_615;
wire n_614;
wire n_617;
wire n_616;
wire n_619;
wire n_618;
wire n_621;
wire n_620;
wire n_623;
wire n_622;
wire n_625;
wire n_624;
wire n_627;
wire n_626;
wire n_167;
wire n_628;
wire n_168;
wire n_630;
wire n_1030;
wire n_1053;
wire n_1076;
wire n_633;
wire n_632;
wire n_1099;
wire n_1122;
wire n_1145;
wire n_635;
wire n_634;
wire n_1168;
wire n_1191;
wire n_1214;
wire n_637;
wire n_636;
wire n_1237;
wire n_1260;
wire n_1283;
wire n_639;
wire n_638;
wire n_1306;
wire n_1329;
wire n_1352;
wire n_641;
wire n_640;
wire n_1375;
wire n_1398;
wire n_1421;
wire n_643;
wire n_642;
wire n_1444;
wire n_1467;
wire n_645;
wire n_644;
wire n_647;
wire n_646;
wire n_649;
wire n_648;
wire n_651;
wire n_650;
wire n_653;
wire n_652;
wire n_655;
wire n_654;
wire n_657;
wire n_656;
wire n_659;
wire n_658;
wire n_661;
wire n_660;
wire n_663;
wire n_662;
wire n_665;
wire n_169;
wire n_504;
wire n_461;
wire n_1029;
wire n_1052;
wire n_1075;
wire n_671;
wire n_670;
wire n_1098;
wire n_1121;
wire n_1144;
wire n_673;
wire n_672;
wire n_1167;
wire n_1190;
wire n_1213;
wire n_675;
wire n_674;
wire n_1236;
wire n_1259;
wire n_1282;
wire n_677;
wire n_676;
wire n_1305;
wire n_1328;
wire n_1351;
wire n_679;
wire n_678;
wire n_1374;
wire n_1397;
wire n_1420;
wire n_681;
wire n_680;
wire n_1443;
wire n_683;
wire n_682;
wire n_685;
wire n_684;
wire n_687;
wire n_686;
wire n_689;
wire n_688;
wire n_691;
wire n_690;
wire n_693;
wire n_692;
wire n_695;
wire n_694;
wire n_697;
wire n_696;
wire n_699;
wire n_698;
wire n_701;
wire n_505;
wire n_509;
wire n_507;
wire n_1028;
wire n_1051;
wire n_1074;
wire n_707;
wire n_706;
wire n_1097;
wire n_1120;
wire n_1143;
wire n_709;
wire n_708;
wire n_1166;
wire n_1189;
wire n_1212;
wire n_711;
wire n_710;
wire n_1235;
wire n_1258;
wire n_1281;
wire n_713;
wire n_712;
wire n_1304;
wire n_1327;
wire n_1350;
wire n_715;
wire n_714;
wire n_1373;
wire n_1396;
wire n_1419;
wire n_717;
wire n_716;
wire n_719;
wire n_718;
wire n_721;
wire n_720;
wire n_723;
wire n_722;
wire n_725;
wire n_724;
wire n_727;
wire n_726;
wire n_511;
wire n_728;
wire n_513;
wire n_730;
wire n_733;
wire n_732;
wire n_735;
wire n_515;
wire n_519;
wire n_517;
wire n_1027;
wire n_1050;
wire n_1073;
wire n_741;
wire n_740;
wire n_1096;
wire n_1119;
wire n_1142;
wire n_743;
wire n_742;
wire n_1165;
wire n_1188;
wire n_1211;
wire n_745;
wire n_744;
wire n_1234;
wire n_1257;
wire n_1280;
wire n_747;
wire n_746;
wire n_1303;
wire n_1326;
wire n_1349;
wire n_749;
wire n_748;
wire n_1372;
wire n_1395;
wire n_751;
wire n_750;
wire n_753;
wire n_752;
wire n_755;
wire n_754;
wire n_757;
wire n_521;
wire n_759;
wire n_523;
wire n_527;
wire n_525;
wire n_531;
wire n_529;
wire n_1700;
wire n_535;
wire n_533;
wire n_1026;
wire n_1049;
wire n_1072;
wire n_537;
wire n_772;
wire n_1095;
wire n_1118;
wire n_1141;
wire n_539;
wire n_774;
wire n_1371;
wire n_541;
wire n_782;
wire n_543;
wire n_784;
wire n_1688;
wire n_547;
wire n_545;
wire n_1690;
wire n_1691;
wire n_549;
wire n_548;
wire n_631;
wire n_629;
wire n_666;
wire n_664;
wire n_1654;
wire n_1639;
wire n_1634;
wire n_1633;
wire n_1632;
wire n_1631;
wire n_1630;
wire n_1629;
wire n_1678;
wire n_1640;
wire n_1677;
wire n_1641;
wire n_1676;
wire n_1642;
wire n_1675;
wire n_1643;
wire n_1674;
wire n_1644;
wire n_1673;
wire n_1645;
wire n_667;
wire n_1672;
wire n_1646;
wire n_668;
wire n_1670;
wire n_1647;
wire n_669;
wire n_1625;
wire n_700;
wire n_1669;
wire n_1648;
wire n_702;
wire n_1628;
wire n_703;
wire n_1668;
wire n_1649;
wire n_704;
wire n_705;
wire n_1667;
wire n_1650;
wire n_729;
wire n_1666;
wire n_1651;
wire n_731;
wire n_1665;
wire n_1652;
wire n_734;
wire n_1664;
wire n_1653;
wire n_736;
wire n_1663;
wire n_1662;
wire n_1661;
wire n_1660;
wire n_1659;
wire n_737;
wire n_1658;
wire n_738;
wire n_1657;
wire n_739;
wire n_1656;
wire n_1655;
wire n_756;
wire n_973;
wire n_1582;
wire n_1763;
wire n_1584;
wire n_1605;
wire n_1593;
wire n_1592;
wire n_1589;
wire n_1590;
wire n_1587;
wire n_1748;
wire n_1751;
wire n_1594;
wire n_1588;
wire n_1747;
wire n_1750;
wire n_1689;
wire n_1591;
wire n_1749;
wire n_764;
wire n_760;
wire n_921;
wire n_769;
wire n_1713;
wire n_1708;
wire n_1604;
wire n_1603;
wire n_1595;
wire n_1599;
wire n_1601;
wire n_1600;
wire n_1597;
wire n_1596;
wire n_1756;
wire n_1744;
wire n_1752;
wire n_1707;
wire n_1704;
wire n_1609;
wire n_1598;
wire n_770;
wire n_1757;
wire n_1602;
wire n_1709;
wire n_1710;
wire n_1775;
wire n_761;
wire n_1745;
wire n_1742;
wire n_1606;
wire n_1740;
wire n_1738;
wire n_1607;
wire n_977;
wire n_1705;
wire n_1701;
wire n_1777;
wire n_1778;
wire n_1729;
wire n_1616;
wire n_1615;
wire n_1612;
wire n_1613;
wire n_1610;
wire n_1759;
wire n_1671;
wire n_1617;
wire n_1611;
wire n_1697;
wire n_1695;
wire n_1758;
wire n_1699;
wire n_1696;
wire n_1754;
wire n_1614;
wire n_1753;
wire n_1755;
wire n_1703;
wire n_1698;
wire n_1761;
wire n_1762;
wire n_1720;
wire n_1624;
wire n_1718;
wire n_1620;
wire n_1716;
wire n_1618;
wire n_1791;
wire n_1770;
wire n_1769;
wire n_1693;
wire n_1686;
wire n_1719;
wire n_1694;
wire n_1692;
wire n_1804;
wire n_1810;
wire n_1627;
wire n_1626;
wire n_1784;
wire n_1796;
wire n_1806;
wire n_1800;
wire n_1811;
wire n_1637;
wire n_1635;
wire n_1765;
wire n_1767;
wire n_1636;
wire n_1638;
wire n_1819;
wire n_1821;
wire n_1815;
wire n_1795;
wire n_1812;
wire n_1760;
wire n_758;
wire n_771;
wire n_1513;
wire n_1702;
wire n_762;
wire n_1569;
wire n_954;
wire n_955;
wire n_1724;
wire n_1721;
wire n_763;
wire n_1722;
wire n_1773;
wire n_1776;
wire n_768;
wire n_1712;
wire n_1711;
wire n_1706;
wire n_1586;
wire n_1583;
wire n_938;
wire n_773;
wire n_1813;
wire n_1451;
wire n_1474;
wire n_1497;
wire n_353;
wire n_352;
wire n_1382;
wire n_1405;
wire n_1428;
wire n_351;
wire n_350;
wire n_1313;
wire n_1336;
wire n_1359;
wire n_349;
wire n_348;
wire n_363;
wire n_362;
wire n_1430;
wire n_1453;
wire n_1476;
wire n_281;
wire n_280;
wire n_1361;
wire n_1384;
wire n_1407;
wire n_279;
wire n_278;
wire n_1292;
wire n_1315;
wire n_1338;
wire n_277;
wire n_276;
wire n_321;
wire n_320;
wire n_1499;
wire n_1522;
wire n_1545;
wire n_283;
wire n_282;
wire n_1544;
wire n_1565;
wire n_319;
wire n_318;
wire n_1520;
wire n_1543;
wire n_1564;
wire n_355;
wire n_354;
wire n_361;
wire n_360;
wire n_1223;
wire n_1246;
wire n_1269;
wire n_275;
wire n_274;
wire n_1154;
wire n_1177;
wire n_1200;
wire n_273;
wire n_272;
wire n_1385;
wire n_1408;
wire n_1431;
wire n_247;
wire n_246;
wire n_1316;
wire n_1339;
wire n_1362;
wire n_245;
wire n_244;
wire n_1247;
wire n_1270;
wire n_1293;
wire n_243;
wire n_242;
wire n_287;
wire n_286;
wire n_323;
wire n_322;
wire n_1268;
wire n_1291;
wire n_1314;
wire n_311;
wire n_310;
wire n_1199;
wire n_1222;
wire n_1245;
wire n_309;
wire n_308;
wire n_1130;
wire n_1153;
wire n_1176;
wire n_307;
wire n_306;
wire n_359;
wire n_358;
wire n_1475;
wire n_1498;
wire n_1521;
wire n_317;
wire n_316;
wire n_1406;
wire n_1429;
wire n_1452;
wire n_315;
wire n_314;
wire n_1337;
wire n_1360;
wire n_1383;
wire n_313;
wire n_312;
wire n_357;
wire n_356;
wire n_367;
wire n_366;
wire n_409;
wire n_408;
wire n_1427;
wire n_1450;
wire n_1473;
wire n_391;
wire n_390;
wire n_1358;
wire n_1381;
wire n_1404;
wire n_389;
wire n_388;
wire n_1289;
wire n_1312;
wire n_1335;
wire n_387;
wire n_386;
wire n_437;
wire n_436;
wire n_1220;
wire n_1243;
wire n_1266;
wire n_385;
wire n_384;
wire n_403;
wire n_402;
wire n_1496;
wire n_1519;
wire n_1542;
wire n_393;
wire n_392;
wire n_401;
wire n_400;
wire n_449;
wire n_448;
wire n_1151;
wire n_1174;
wire n_1197;
wire n_383;
wire n_382;
wire n_1082;
wire n_1105;
wire n_1128;
wire n_381;
wire n_380;
wire n_1175;
wire n_1198;
wire n_1221;
wire n_345;
wire n_344;
wire n_1106;
wire n_1129;
wire n_1152;
wire n_343;
wire n_342;
wire n_399;
wire n_398;
wire n_405;
wire n_404;
wire n_411;
wire n_410;
wire n_455;
wire n_454;
wire n_291;
wire n_290;
wire n_1178;
wire n_1201;
wire n_1224;
wire n_241;
wire n_240;
wire n_1478;
wire n_1501;
wire n_1524;
wire n_219;
wire n_218;
wire n_1409;
wire n_1432;
wire n_1455;
wire n_217;
wire n_216;
wire n_1340;
wire n_1363;
wire n_1386;
wire n_215;
wire n_214;
wire n_253;
wire n_252;
wire n_289;
wire n_288;
wire n_331;
wire n_330;
wire n_329;
wire n_328;
wire n_1244;
wire n_1267;
wire n_1290;
wire n_347;
wire n_346;
wire n_365;
wire n_364;
wire n_371;
wire n_370;
wire n_327;
wire n_326;
wire n_1523;
wire n_1546;
wire n_1567;
wire n_251;
wire n_250;
wire n_1454;
wire n_1477;
wire n_1500;
wire n_249;
wire n_248;
wire n_1566;
wire n_285;
wire n_284;
wire n_325;
wire n_324;
wire n_369;
wire n_368;
wire n_373;
wire n_372;
wire n_415;
wire n_414;
wire n_397;
wire n_396;
wire n_1563;
wire n_395;
wire n_394;
wire n_1541;
wire n_1562;
wire n_435;
wire n_434;
wire n_441;
wire n_440;
wire n_407;
wire n_406;
wire n_451;
wire n_450;
wire n_413;
wire n_412;
wire n_1265;
wire n_1288;
wire n_1311;
wire n_427;
wire n_426;
wire n_1196;
wire n_1219;
wire n_1242;
wire n_425;
wire n_424;
wire n_1127;
wire n_1150;
wire n_1173;
wire n_423;
wire n_422;
wire n_445;
wire n_444;
wire n_1472;
wire n_1495;
wire n_1518;
wire n_433;
wire n_432;
wire n_1403;
wire n_1426;
wire n_1449;
wire n_431;
wire n_430;
wire n_1334;
wire n_1357;
wire n_1380;
wire n_429;
wire n_428;
wire n_443;
wire n_442;
wire n_1058;
wire n_1081;
wire n_1104;
wire n_421;
wire n_420;
wire n_439;
wire n_438;
wire n_447;
wire n_446;
wire n_453;
wire n_452;
wire n_457;
wire n_456;
wire n_459;
wire n_458;
wire n_483;
wire n_482;
wire n_493;
wire n_492;
wire n_481;
wire n_480;
wire n_479;
wire n_478;
wire n_491;
wire n_490;
wire n_499;
wire n_498;
wire n_1172;
wire n_1195;
wire n_1218;
wire n_467;
wire n_466;
wire n_1103;
wire n_1126;
wire n_1149;
wire n_465;
wire n_464;
wire n_1034;
wire n_1057;
wire n_1080;
wire n_463;
wire n_462;
wire n_489;
wire n_488;
wire n_495;
wire n_494;
wire n_1379;
wire n_1402;
wire n_1425;
wire n_473;
wire n_472;
wire n_1310;
wire n_1333;
wire n_1356;
wire n_471;
wire n_470;
wire n_1241;
wire n_1264;
wire n_1287;
wire n_469;
wire n_468;
wire n_487;
wire n_486;
wire n_1517;
wire n_1540;
wire n_1561;
wire n_477;
wire n_476;
wire n_1448;
wire n_1471;
wire n_1494;
wire n_475;
wire n_474;
wire n_485;
wire n_484;
wire n_497;
wire n_496;
wire n_501;
wire n_500;
wire n_503;
wire n_502;
wire n_775;
wire n_524;
wire n_522;
wire n_534;
wire n_542;
wire n_1102;
wire n_1125;
wire n_1148;
wire n_508;
wire n_1033;
wire n_1056;
wire n_1079;
wire n_506;
wire n_532;
wire n_1309;
wire n_1332;
wire n_1355;
wire n_514;
wire n_1240;
wire n_1263;
wire n_1286;
wire n_512;
wire n_1171;
wire n_1194;
wire n_1217;
wire n_510;
wire n_530;
wire n_538;
wire n_1516;
wire n_1539;
wire n_520;
wire n_1447;
wire n_1470;
wire n_1493;
wire n_518;
wire n_1378;
wire n_1401;
wire n_1424;
wire n_516;
wire n_528;
wire n_526;
wire n_536;
wire n_540;
wire n_544;
wire n_546;
wire n_900;
wire n_1271;
wire n_1294;
wire n_1317;
wire n_213;
wire n_212;
wire n_1202;
wire n_1225;
wire n_1248;
wire n_211;
wire n_210;
wire n_1433;
wire n_1456;
wire n_1479;
wire n_189;
wire n_188;
wire n_1364;
wire n_1387;
wire n_1410;
wire n_187;
wire n_186;
wire n_1295;
wire n_1318;
wire n_1341;
wire n_185;
wire n_184;
wire n_223;
wire n_222;
wire n_255;
wire n_254;
wire n_293;
wire n_292;
wire n_259;
wire n_258;
wire n_295;
wire n_294;
wire n_333;
wire n_332;
wire n_1502;
wire n_1525;
wire n_1548;
wire n_191;
wire n_190;
wire n_1547;
wire n_1568;
wire n_221;
wire n_220;
wire n_257;
wire n_256;
wire n_229;
wire n_228;
wire n_227;
wire n_226;
wire n_263;
wire n_262;
wire n_297;
wire n_296;
wire n_335;
wire n_334;
wire n_375;
wire n_374;
wire n_417;
wire n_416;
wire n_460;
wire n_183;
wire n_182;
wire n_195;
wire n_194;
wire n_193;
wire n_192;
wire n_225;
wire n_224;
wire n_261;
wire n_260;
wire n_299;
wire n_298;
wire n_337;
wire n_336;
wire n_377;
wire n_376;
wire n_419;
wire n_418;
wire n_199;
wire n_197;
wire n_231;
wire n_230;
wire n_265;
wire n_264;
wire n_301;
wire n_300;
wire n_339;
wire n_338;
wire n_201;
wire n_233;
wire n_232;
wire n_267;
wire n_266;
wire n_303;
wire n_302;
wire n_341;
wire n_340;
wire n_379;
wire n_378;
wire n_203;
wire n_235;
wire n_234;
wire n_269;
wire n_268;
wire n_305;
wire n_304;
wire n_196;
wire n_175;
wire n_200;
wire n_205;
wire n_204;
wire n_237;
wire n_236;
wire n_177;
wire n_202;
wire n_207;
wire n_206;
wire n_179;
wire n_181;
wire n_209;
wire n_208;
wire n_239;
wire n_238;
wire n_271;
wire n_270;
wire n_121;
wire n_142;
wire n_123;
wire n_149;
wire n_148;
wire n_173;
wire n_172;
wire n_171;
wire n_170;
wire n_176;
wire n_198;
wire n_147;
wire n_145;
wire n_174;
wire n_125;
wire n_146;
wire n_144;
wire n_151;
wire n_150;
wire n_178;
wire n_127;
wire n_129;
wire n_153;
wire n_152;
wire n_131;
wire n_155;
wire n_154;
wire n_180;
wire n_120;
wire n_122;
wire n_101;
wire n_100;
wire n_103;
wire n_102;
wire n_126;
wire n_105;
wire n_104;
wire n_124;
wire n_128;
wire n_107;
wire n_106;
wire n_89;
wire n_87;
wire n_109;
wire n_108;
wire n_130;
wire n_86;
wire n_71;
wire n_69;
wire n_88;
wire n_68;
wire n_55;
wire n_53;
wire n_70;
wire n_29;
wire n_39;
wire n_38;
wire n_27;
wire n_41;
wire n_40;
wire n_52;
wire n_54;
wire n_26;
wire n_19;
wire n_17;
wire n_28;
wire n_7;
wire n_16;
wire n_11;
wire n_18;
wire n_971;
wire n_968;
wire n_975;
wire n_1536;
wire n_987;
wire n_979;
wire n_981;
wire n_989;
wire n_983;
wire n_1621;
wire n_990;
wire n_1608;
wire n_985;
wire n_998;
wire n_991;
wire n_1008;
wire n_1010;
wire n_1007;
wire n_1011;
wire n_1005;
wire n_1009;
wire n_1164;
wire n_1210;
wire n_1187;
wire n_1256;
wire n_1226;
wire n_1233;
wire n_1249;
wire n_1490;
wire n_1272;
wire n_1279;
wire n_1348;
wire n_1325;
wire n_1302;
wire n_1623;
wire n_1622;
wire n_1619;
wire n_1585;
wire n_1157;
wire n_1180;
wire n_1203;
wire n_945;
wire n_944;
wire n_1156;
wire n_1179;
wire n_961;
wire n_960;
wire n_1087;
wire n_1110;
wire n_1133;
wire n_959;
wire n_958;
wire n_1018;
wire n_1041;
wire n_1064;
wire n_957;
wire n_956;
wire n_965;
wire n_964;
wire n_1088;
wire n_1111;
wire n_1134;
wire n_943;
wire n_942;
wire n_1019;
wire n_1042;
wire n_1065;
wire n_941;
wire n_940;
wire n_1158;
wire n_1181;
wire n_1204;
wire n_927;
wire n_926;
wire n_1089;
wire n_1112;
wire n_1135;
wire n_925;
wire n_924;
wire n_1020;
wire n_1043;
wire n_1066;
wire n_923;
wire n_922;
wire n_947;
wire n_946;
wire n_963;
wire n_962;
wire n_1159;
wire n_1182;
wire n_1205;
wire n_907;
wire n_906;
wire n_1090;
wire n_1113;
wire n_1136;
wire n_905;
wire n_904;
wire n_1227;
wire n_929;
wire n_928;
wire n_949;
wire n_948;
wire n_1021;
wire n_1044;
wire n_1067;
wire n_903;
wire n_902;
wire n_1160;
wire n_1183;
wire n_1206;
wire n_885;
wire n_884;
wire n_1091;
wire n_1114;
wire n_1137;
wire n_883;
wire n_882;
wire n_1022;
wire n_1045;
wire n_1068;
wire n_881;
wire n_880;
wire n_911;
wire n_910;
wire n_1229;
wire n_1252;
wire n_1275;
wire n_887;
wire n_886;
wire n_1228;
wire n_1251;
wire n_909;
wire n_908;
wire n_931;
wire n_930;
wire n_951;
wire n_950;
wire n_967;
wire n_966;
wire n_933;
wire n_932;
wire n_953;
wire n_952;
wire n_969;
wire n_1679;
wire n_1086;
wire n_1109;
wire n_1132;
wire n_1680;
wire n_972;
wire n_1017;
wire n_1040;
wire n_1063;
wire n_1681;
wire n_970;
wire n_1682;
wire n_976;
wire n_1155;
wire n_1683;
wire n_974;
wire n_1684;
wire n_978;
wire n_1685;
wire n_980;
wire n_1230;
wire n_1253;
wire n_1276;
wire n_863;
wire n_862;
wire n_1161;
wire n_1184;
wire n_1207;
wire n_861;
wire n_860;
wire n_1092;
wire n_1115;
wire n_1138;
wire n_859;
wire n_858;
wire n_889;
wire n_888;
wire n_913;
wire n_912;
wire n_935;
wire n_934;
wire n_915;
wire n_914;
wire n_893;
wire n_892;
wire n_1023;
wire n_1046;
wire n_1069;
wire n_857;
wire n_856;
wire n_1231;
wire n_1254;
wire n_1277;
wire n_837;
wire n_836;
wire n_1162;
wire n_1185;
wire n_1208;
wire n_835;
wire n_834;
wire n_1299;
wire n_865;
wire n_864;
wire n_891;
wire n_890;
wire n_1093;
wire n_1116;
wire n_1139;
wire n_833;
wire n_832;
wire n_1024;
wire n_1047;
wire n_1070;
wire n_831;
wire n_830;
wire n_1232;
wire n_1255;
wire n_1278;
wire n_809;
wire n_808;
wire n_1163;
wire n_1186;
wire n_1209;
wire n_807;
wire n_806;
wire n_1094;
wire n_1117;
wire n_1140;
wire n_805;
wire n_804;
wire n_841;
wire n_840;
wire n_867;
wire n_866;
wire n_1301;
wire n_1324;
wire n_1347;
wire n_811;
wire n_810;
wire n_1300;
wire n_1323;
wire n_839;
wire n_838;
wire n_869;
wire n_868;
wire n_895;
wire n_894;
wire n_917;
wire n_916;
wire n_937;
wire n_936;
wire n_1687;
wire n_845;
wire n_844;
wire n_1025;
wire n_1048;
wire n_1071;
wire n_803;
wire n_802;
wire n_781;
wire n_779;
wire n_777;
wire n_813;
wire n_812;
wire n_843;
wire n_842;
wire n_873;
wire n_872;
wire n_871;
wire n_870;
wire n_897;
wire n_896;
wire n_919;
wire n_918;
wire n_815;
wire n_814;
wire n_847;
wire n_846;
wire n_875;
wire n_874;
wire n_899;
wire n_898;
wire n_920;
wire n_819;
wire n_818;
wire n_817;
wire n_816;
wire n_849;
wire n_848;
wire n_821;
wire n_820;
wire n_851;
wire n_850;
wire n_877;
wire n_876;
wire n_901;
wire n_823;
wire n_822;
wire n_795;
wire n_825;
wire n_824;
wire n_853;
wire n_852;
wire n_797;
wire n_827;
wire n_826;
wire n_794;
wire n_765;
wire n_767;
wire n_766;
wire n_799;
wire n_798;
wire n_796;
wire n_1715;
wire n_1714;
wire n_1774;
wire n_1772;
wire n_1768;
wire n_1717;
wire n_1766;
wire n_1725;
wire n_1730;
wire n_1727;
wire n_1764;
wire n_1728;
wire n_1726;
wire n_1731;
wire n_1737;
wire n_1732;
wire n_1733;
wire n_1736;
wire n_1734;
wire n_1743;
wire n_1739;
wire n_1735;
wire n_1741;
wire n_1746;
wire n_1771;
wire n_1085;
wire n_1108;
wire n_1131;
wire n_1779;
wire n_984;
wire n_1016;
wire n_1039;
wire n_1062;
wire n_1780;
wire n_982;
wire n_1781;
wire n_986;
wire n_1782;
wire n_988;
wire n_1783;
wire n_1787;
wire n_1785;
wire n_1786;
wire n_1790;
wire n_1789;
wire n_1788;
wire n_1014;
wire n_1037;
wire n_1060;
wire n_1001;
wire n_1000;
wire n_1015;
wire n_1038;
wire n_1061;
wire n_993;
wire n_992;
wire n_1084;
wire n_1107;
wire n_995;
wire n_994;
wire n_1083;
wire n_1003;
wire n_1002;
wire n_997;
wire n_996;
wire n_1792;
wire n_1004;
wire n_1013;
wire n_1036;
wire n_1059;
wire n_1793;
wire n_1006;
wire n_1794;
wire n_999;
wire n_1797;
wire n_1798;
wire n_1799;
wire n_1801;
wire n_1802;
wire n_1803;
wire n_1805;
wire n_1807;
wire n_1808;
wire n_1809;
wire n_1012;
wire n_1035;
wire n_1814;
wire n_1820;
wire n_1818;
wire n_1816;
wire n_1817;
wire hfn_ipo_n6;


INV_X1 i_1340 (.ZN (n_1821), .A (n_1812));
INV_X1 i_1339 (.ZN (n_1820), .A (n_1798));
INV_X1 i_1338 (.ZN (n_1819), .A (n_1795));
OAI21_X1 i_1337 (.ZN (n_1818), .A (n_1802), .B1 (n_1792), .B2 (n_1794));
OAI211_X1 i_1336 (.ZN (n_1817), .A (n_1786), .B (n_1805), .C1 (n_1803), .C2 (n_1787));
INV_X1 i_1335 (.ZN (n_1816), .A (n_1817));
OAI221_X1 i_1334 (.ZN (n_1815), .A (n_1820), .B1 (n_1797), .B2 (n_1799), .C1 (n_1818), .C2 (n_1816));
AOI22_X1 i_1333 (.ZN (n_1814), .A1 (n_1812), .A2 (n_1819), .B1 (n_1821), .B2 (n_1795));
XNOR2_X1 i_1332 (.ZN (Res_imm[45]), .A (n_1815), .B (n_1814));
NOR2_X1 i_1331 (.ZN (n_1012), .A1 (hfn_ipo_n6), .A2 (n_1653));
NOR2_X1 i_1330 (.ZN (n_1035), .A1 (hfn_ipo_n6), .A2 (n_1678));
FA_X1 i_1329 (.CO (n_1813), .S (n_1812), .A (n_1012), .B (n_1035), .CI (n_1793));
INV_X1 i_1328 (.ZN (n_1811), .A (n_1799));
NOR2_X1 i_1327 (.ZN (n_1810), .A1 (n_1806), .A2 (n_1801));
XOR2_X1 i_1326 (.Z (Res_imm[44]), .A (n_1808), .B (n_1809));
NOR2_X1 i_1325 (.ZN (n_1809), .A1 (n_1798), .A2 (n_1797));
NAND2_X1 i_1324 (.ZN (n_1808), .A1 (n_1807), .A2 (n_1799));
OAI21_X1 i_1323 (.ZN (n_1807), .A (n_1802), .B1 (n_1804), .B2 (n_1806));
INV_X1 i_1322 (.ZN (n_1806), .A (n_1805));
NAND2_X1 i_1321 (.ZN (n_1805), .A1 (n_1796), .A2 (n_1784));
AOI21_X1 i_1320 (.ZN (n_1804), .A (n_1803), .B1 (n_1787), .B2 (n_1786));
NOR2_X1 i_1319 (.ZN (n_1803), .A1 (n_1685), .A2 (n_1783));
NOR2_X1 i_1318 (.ZN (n_1802), .A1 (n_1801), .A2 (n_1800));
NOR2_X1 i_1317 (.ZN (n_1801), .A1 (n_1796), .A2 (n_1784));
NOR2_X1 i_1316 (.ZN (n_1800), .A1 (n_1004), .A2 (n_999));
NAND2_X1 i_1315 (.ZN (n_1799), .A1 (n_1004), .A2 (n_999));
AND2_X1 i_1314 (.ZN (n_1798), .A1 (n_1792), .A2 (n_1794));
NOR2_X1 i_1313 (.ZN (n_1797), .A1 (n_1792), .A2 (n_1794));
NOR2_X1 i_1312 (.ZN (n_1014), .A1 (hfn_ipo_n6), .A2 (n_1651));
NOR2_X1 i_1311 (.ZN (n_1037), .A1 (n_1678), .A2 (n_1652));
NOR2_X1 i_1310 (.ZN (n_1060), .A1 (n_1677), .A2 (n_1653));
NOR2_X1 i_1309 (.ZN (n_1083), .A1 (n_1676), .A2 (hfn_ipo_n6));
NOR2_X1 i_1308 (.ZN (n_1015), .A1 (n_1650), .A2 (hfn_ipo_n6));
NOR2_X1 i_1307 (.ZN (n_1038), .A1 (n_1678), .A2 (n_1651));
NOR2_X1 i_1306 (.ZN (n_1061), .A1 (n_1677), .A2 (n_1652));
NOR2_X1 i_1305 (.ZN (n_1084), .A1 (n_1676), .A2 (n_1653));
NOR2_X1 i_1304 (.ZN (n_1107), .A1 (n_1675), .A2 (hfn_ipo_n6));
NOR2_X1 i_1303 (.ZN (n_1013), .A1 (n_1652), .A2 (hfn_ipo_n6));
NOR2_X1 i_1302 (.ZN (n_1036), .A1 (n_1653), .A2 (n_1678));
NOR2_X1 i_1301 (.ZN (n_1059), .A1 (n_1677), .A2 (hfn_ipo_n6));
FA_X1 i_1300 (.CO (n_999), .S (n_1796), .A (n_1781), .B (n_1782), .CI (n_996));
FA_X1 i_1299 (.CO (n_1795), .S (n_1794), .A (n_1001), .B (n_1006), .CI (n_1003));
FA_X1 i_1298 (.CO (n_1793), .S (n_1006), .A (n_1013), .B (n_1036), .CI (n_1059));
FA_X1 i_1297 (.CO (n_1792), .S (n_1004), .A (n_1000), .B (n_1002), .CI (n_997));
FA_X1 i_1296 (.CO (n_997), .S (n_996), .A (n_1780), .B (n_994), .CI (n_992));
FA_X1 i_1295 (.CO (n_1003), .S (n_1002), .A (n_1083), .B (n_993), .CI (n_995));
FA_X1 i_1294 (.CO (n_995), .S (n_994), .A (n_1084), .B (n_1107), .CI (n_1779));
FA_X1 i_1293 (.CO (n_993), .S (n_992), .A (n_1015), .B (n_1038), .CI (n_1061));
FA_X1 i_1292 (.CO (n_1001), .S (n_1000), .A (n_1014), .B (n_1037), .CI (n_1060));
NOR2_X1 i_1291 (.ZN (n_1791), .A1 (n_1687), .A2 (n_1679));
NOR2_X1 i_1290 (.ZN (n_1790), .A1 (n_1774), .A2 (n_1771));
NOR3_X1 i_1289 (.ZN (n_1789), .A1 (n_1774), .A2 (n_1791), .A3 (n_1769));
OAI211_X2 i_1288 (.ZN (n_1788), .A (n_1719), .B (n_1768), .C1 (n_1766), .C2 (n_1720));
AOI211_X2 i_1287 (.ZN (n_1787), .A (n_1772), .B (n_1790), .C1 (n_1789), .C2 (n_1788));
NAND2_X1 i_1286 (.ZN (n_1786), .A1 (n_1783), .A2 (n_1685));
OAI21_X1 i_1285 (.ZN (n_1785), .A (n_1786), .B1 (n_1783), .B2 (n_1685));
XOR2_X1 i_1284 (.Z (Res_imm[41]), .A (n_1787), .B (n_1785));
NOR2_X1 i_1283 (.ZN (n_1085), .A1 (n_1676), .A2 (n_1652));
NOR2_X1 i_1282 (.ZN (n_1108), .A1 (n_1675), .A2 (n_1653));
NOR2_X1 i_1281 (.ZN (n_1131), .A1 (n_1674), .A2 (hfn_ipo_n6));
NOR2_X1 i_1280 (.ZN (n_1016), .A1 (hfn_ipo_n6), .A2 (n_1649));
NOR2_X1 i_1279 (.ZN (n_1039), .A1 (n_1678), .A2 (n_1650));
NOR2_X1 i_1278 (.ZN (n_1062), .A1 (n_1677), .A2 (n_1651));
FA_X1 i_1277 (.CO (n_1784), .S (n_1783), .A (n_1682), .B (n_1684), .CI (n_988));
FA_X1 i_1276 (.CO (n_1782), .S (n_988), .A (n_984), .B (n_982), .CI (n_986));
FA_X1 i_1275 (.CO (n_1781), .S (n_986), .A (n_1680), .B (n_1681), .CI (n_1683));
FA_X1 i_1274 (.CO (n_1780), .S (n_982), .A (n_1016), .B (n_1039), .CI (n_1062));
FA_X1 i_1273 (.CO (n_1779), .S (n_984), .A (n_1085), .B (n_1108), .CI (n_1131));
INV_X1 i_1272 (.ZN (n_1778), .A (n_1701));
INV_X1 i_1271 (.ZN (n_1777), .A (n_1705));
INV_X1 i_1270 (.ZN (n_1776), .A (n_769));
INV_X1 i_1269 (.ZN (n_1775), .A (n_761));
NOR2_X1 i_1268 (.ZN (n_1774), .A1 (n_969), .A2 (n_980));
AND2_X1 i_1267 (.ZN (n_1772), .A1 (n_969), .A2 (n_980));
NAND2_X1 i_1266 (.ZN (n_1771), .A1 (n_1679), .A2 (n_1687));
INV_X1 i_1265 (.ZN (n_1770), .A (n_1771));
NOR2_X1 i_1264 (.ZN (n_1769), .A1 (n_1686), .A2 (n_1693));
NAND2_X1 i_1263 (.ZN (n_1768), .A1 (n_1686), .A2 (n_1693));
NOR2_X1 i_1262 (.ZN (n_1766), .A1 (n_1692), .A2 (n_1694));
NAND2_X1 i_1261 (.ZN (n_1764), .A1 (n_920), .A2 (n_901));
INV_X1 i_1260 (.ZN (n_1762), .A (n_1764));
NOR2_X1 i_1259 (.ZN (n_1761), .A1 (n_920), .A2 (n_901));
NAND2_X1 i_1258 (.ZN (n_1760), .A1 (n_1695), .A2 (n_1697));
NOR2_X1 i_1257 (.ZN (n_1759), .A1 (n_1695), .A2 (n_1697));
NOR2_X1 i_1256 (.ZN (n_1758), .A1 (n_1696), .A2 (n_1699));
NAND2_X1 i_1255 (.ZN (n_1755), .A1 (n_1698), .A2 (n_1703));
NAND2_X1 i_1254 (.ZN (n_1754), .A1 (n_1696), .A2 (n_1699));
NOR2_X1 i_1253 (.ZN (n_1753), .A1 (n_1698), .A2 (n_1703));
NAND2_X1 i_1252 (.ZN (n_1752), .A1 (n_1704), .A2 (n_1707));
AND2_X1 i_1251 (.ZN (n_1751), .A1 (n_1712), .A2 (n_168));
AOI21_X1 i_1250 (.ZN (n_1746), .A (n_768), .B1 (n_760), .B2 (n_758));
AOI221_X1 i_1249 (.ZN (n_1745), .A (n_1746), .B1 (n_1708), .B2 (n_1713), .C1 (n_1776), .C2 (n_1751));
AND2_X1 i_1248 (.ZN (n_1744), .A1 (n_1706), .A2 (n_1711));
NOR2_X1 i_1247 (.ZN (n_1743), .A1 (n_768), .A2 (n_764));
INV_X1 i_1246 (.ZN (n_1742), .A (n_1743));
OAI21_X1 i_1245 (.ZN (n_1741), .A (n_762), .B1 (n_1586), .B2 (n_1585));
AOI21_X1 i_1244 (.ZN (n_1740), .A (n_1741), .B1 (n_775), .B2 (n_900));
INV_X1 i_1243 (.ZN (n_1739), .A (n_1740));
NAND2_X1 i_1242 (.ZN (n_1738), .A1 (n_1536), .A2 (n_771));
NOR2_X1 i_1241 (.ZN (n_1737), .A1 (n_1701), .A2 (n_1705));
NOR2_X1 i_1240 (.ZN (n_1736), .A1 (n_1709), .A2 (n_1710));
AOI21_X2 i_1239 (.ZN (n_1735), .A (n_1738), .B1 (n_979), .B2 (n_987));
OAI21_X1 i_1238 (.ZN (n_1734), .A (n_1743), .B1 (n_1739), .B2 (n_1735));
AOI21_X1 i_1237 (.ZN (n_1733), .A (n_1736), .B1 (n_1745), .B2 (n_1734));
NOR3_X1 i_1236 (.ZN (n_1732), .A1 (n_1775), .A2 (n_1744), .A3 (n_1733));
OR3_X2 i_1235 (.ZN (n_1731), .A1 (n_770), .A2 (n_1737), .A3 (n_1732));
OAI221_X2 i_1234 (.ZN (n_1730), .A (n_1731), .B1 (n_1778), .B2 (n_1777), .C1 (n_1752), .C2 (n_1737));
INV_X1 i_1233 (.ZN (n_1729), .A (n_1730));
OR3_X1 i_1232 (.ZN (n_1728), .A1 (n_1761), .A2 (n_1758), .A3 (n_1759));
NOR2_X1 i_1231 (.ZN (n_1727), .A1 (n_1753), .A2 (n_1728));
AND2_X1 i_1230 (.ZN (n_1726), .A1 (n_1755), .A2 (n_1754));
OAI221_X1 i_1229 (.ZN (n_1725), .A (n_1764), .B1 (n_1761), .B2 (n_1760), .C1 (n_1728), .C2 (n_1726));
AOI21_X4 i_1228 (.ZN (n_1720), .A (n_1725), .B1 (n_1730), .B2 (n_1727));
NAND2_X1 i_1227 (.ZN (n_1719), .A1 (n_1692), .A2 (n_1694));
AOI21_X1 i_1226 (.ZN (n_1718), .A (n_1766), .B1 (n_1720), .B2 (n_1719));
INV_X1 i_1225 (.ZN (n_1717), .A (n_1718));
AOI21_X1 i_1224 (.ZN (n_1716), .A (n_1769), .B1 (n_1768), .B2 (n_1717));
OR2_X1 i_1223 (.ZN (n_1715), .A1 (n_1774), .A2 (n_1772));
OAI22_X1 i_1222 (.ZN (n_1714), .A1 (n_1679), .A2 (n_1687), .B1 (n_1770), .B2 (n_1716));
XOR2_X2 i_1221 (.Z (Res_imm[40]), .A (n_1715), .B (n_1714));
NOR2_X1 i_1220 (.ZN (n_1156), .A1 (n_1673), .A2 (n_1653));
NOR2_X1 i_1219 (.ZN (n_1179), .A1 (n_1672), .A2 (hfn_ipo_n6));
NOR2_X1 i_1218 (.ZN (n_1157), .A1 (n_1673), .A2 (n_1652));
NOR2_X1 i_1217 (.ZN (n_1180), .A1 (n_1653), .A2 (n_1672));
NOR2_X1 i_1216 (.ZN (n_1203), .A1 (hfn_ipo_n6), .A2 (n_1670));
NOR2_X1 i_1215 (.ZN (n_1087), .A1 (n_1676), .A2 (n_1650));
NOR2_X1 i_1214 (.ZN (n_1110), .A1 (n_1675), .A2 (n_1651));
NOR2_X1 i_1213 (.ZN (n_1133), .A1 (n_1652), .A2 (n_1674));
NOR2_X1 i_1212 (.ZN (n_1018), .A1 (hfn_ipo_n6), .A2 (n_1647));
NOR2_X1 i_1211 (.ZN (n_1041), .A1 (n_1678), .A2 (n_1648));
NOR2_X1 i_1210 (.ZN (n_1064), .A1 (n_1677), .A2 (n_1649));
NOR2_X1 i_1209 (.ZN (n_1088), .A1 (n_1676), .A2 (n_1649));
NOR2_X1 i_1208 (.ZN (n_1111), .A1 (n_1650), .A2 (n_1675));
NOR2_X1 i_1207 (.ZN (n_1134), .A1 (n_1651), .A2 (n_1674));
NOR2_X1 i_1206 (.ZN (n_1019), .A1 (hfn_ipo_n6), .A2 (n_1646));
NOR2_X1 i_1205 (.ZN (n_1042), .A1 (n_1647), .A2 (n_1678));
NOR2_X1 i_1204 (.ZN (n_1065), .A1 (n_1648), .A2 (n_1677));
NOR2_X1 i_1203 (.ZN (n_1158), .A1 (n_1673), .A2 (n_1651));
NOR2_X1 i_1202 (.ZN (n_1181), .A1 (n_1672), .A2 (n_1652));
NOR2_X1 i_1201 (.ZN (n_1204), .A1 (n_1653), .A2 (n_1670));
NOR2_X1 i_1200 (.ZN (n_1089), .A1 (n_1676), .A2 (n_1648));
NOR2_X1 i_1199 (.ZN (n_1112), .A1 (n_1675), .A2 (n_1649));
NOR2_X1 i_1198 (.ZN (n_1135), .A1 (n_1650), .A2 (n_1674));
NOR2_X1 i_1197 (.ZN (n_1020), .A1 (hfn_ipo_n6), .A2 (n_1645));
NOR2_X1 i_1196 (.ZN (n_1043), .A1 (n_1678), .A2 (n_1646));
NOR2_X1 i_1195 (.ZN (n_1066), .A1 (n_1647), .A2 (n_1677));
NOR2_X1 i_1194 (.ZN (n_1227), .A1 (hfn_ipo_n6), .A2 (n_1669));
NOR2_X1 i_1193 (.ZN (n_1159), .A1 (n_1673), .A2 (n_1650));
NOR2_X1 i_1192 (.ZN (n_1182), .A1 (n_1672), .A2 (n_1651));
NOR2_X1 i_1191 (.ZN (n_1205), .A1 (n_1652), .A2 (n_1670));
NOR2_X1 i_1190 (.ZN (n_1090), .A1 (n_1676), .A2 (n_1647));
NOR2_X1 i_1189 (.ZN (n_1113), .A1 (n_1675), .A2 (n_1648));
NOR2_X1 i_1188 (.ZN (n_1136), .A1 (n_1674), .A2 (n_1649));
NOR2_X1 i_1187 (.ZN (n_1021), .A1 (hfn_ipo_n6), .A2 (n_1644));
NOR2_X1 i_1186 (.ZN (n_1044), .A1 (n_1678), .A2 (n_1645));
NOR2_X1 i_1185 (.ZN (n_1067), .A1 (n_1677), .A2 (n_1646));
NOR2_X1 i_1184 (.ZN (n_1160), .A1 (n_1673), .A2 (n_1649));
NOR2_X1 i_1183 (.ZN (n_1183), .A1 (n_1672), .A2 (n_1650));
NOR2_X1 i_1182 (.ZN (n_1206), .A1 (n_1670), .A2 (n_1651));
NOR2_X1 i_1181 (.ZN (n_1091), .A1 (n_1676), .A2 (n_1646));
NOR2_X1 i_1180 (.ZN (n_1114), .A1 (n_1675), .A2 (n_1647));
NOR2_X1 i_1179 (.ZN (n_1137), .A1 (n_1674), .A2 (n_1648));
NOR2_X1 i_1178 (.ZN (n_1022), .A1 (hfn_ipo_n6), .A2 (n_1643));
NOR2_X1 i_1177 (.ZN (n_1045), .A1 (n_1678), .A2 (n_1644));
NOR2_X1 i_1176 (.ZN (n_1068), .A1 (n_1677), .A2 (n_1645));
NOR2_X1 i_1175 (.ZN (n_1228), .A1 (n_1653), .A2 (n_1669));
NOR2_X1 i_1174 (.ZN (n_1251), .A1 (hfn_ipo_n6), .A2 (n_1668));
NOR2_X1 i_1173 (.ZN (n_1229), .A1 (n_1652), .A2 (n_1669));
NOR2_X1 i_1172 (.ZN (n_1252), .A1 (n_1653), .A2 (n_1668));
NOR2_X1 i_1171 (.ZN (n_1275), .A1 (hfn_ipo_n6), .A2 (n_1667));
NOR2_X1 i_1170 (.ZN (n_1086), .A1 (n_1676), .A2 (n_1651));
NOR2_X1 i_1169 (.ZN (n_1109), .A1 (n_1652), .A2 (n_1675));
NOR2_X1 i_1168 (.ZN (n_1132), .A1 (n_1653), .A2 (n_1674));
NOR2_X1 i_1167 (.ZN (n_1017), .A1 (hfn_ipo_n6), .A2 (n_1648));
NOR2_X1 i_1166 (.ZN (n_1040), .A1 (n_1678), .A2 (n_1649));
NOR2_X1 i_1165 (.ZN (n_1063), .A1 (n_1650), .A2 (n_1677));
NOR2_X1 i_1164 (.ZN (n_1155), .A1 (n_1673), .A2 (hfn_ipo_n6));
NOR2_X1 i_1163 (.ZN (n_1230), .A1 (n_1651), .A2 (n_1669));
NOR2_X1 i_1162 (.ZN (n_1253), .A1 (n_1652), .A2 (n_1668));
NOR2_X1 i_1161 (.ZN (n_1276), .A1 (n_1653), .A2 (n_1667));
NOR2_X1 i_1160 (.ZN (n_1161), .A1 (n_1673), .A2 (n_1648));
NOR2_X1 i_1159 (.ZN (n_1184), .A1 (n_1672), .A2 (n_1649));
NOR2_X1 i_1158 (.ZN (n_1207), .A1 (n_1670), .A2 (n_1650));
NOR2_X1 i_1157 (.ZN (n_1092), .A1 (n_1676), .A2 (n_1645));
NOR2_X1 i_1156 (.ZN (n_1115), .A1 (n_1675), .A2 (n_1646));
NOR2_X1 i_1155 (.ZN (n_1138), .A1 (n_1674), .A2 (n_1647));
NOR2_X1 i_1154 (.ZN (n_1023), .A1 (hfn_ipo_n6), .A2 (n_1642));
NOR2_X1 i_1153 (.ZN (n_1046), .A1 (n_1678), .A2 (n_1643));
NOR2_X1 i_1152 (.ZN (n_1069), .A1 (n_1677), .A2 (n_1644));
NOR2_X1 i_1151 (.ZN (n_1299), .A1 (hfn_ipo_n6), .A2 (n_1666));
NOR2_X1 i_1150 (.ZN (n_1231), .A1 (n_1650), .A2 (n_1669));
NOR2_X1 i_1149 (.ZN (n_1254), .A1 (n_1651), .A2 (n_1668));
NOR2_X1 i_1148 (.ZN (n_1277), .A1 (n_1652), .A2 (n_1667));
NOR2_X1 i_1147 (.ZN (n_1162), .A1 (n_1673), .A2 (n_1647));
NOR2_X1 i_1146 (.ZN (n_1185), .A1 (n_1672), .A2 (n_1648));
NOR2_X1 i_1145 (.ZN (n_1208), .A1 (n_1670), .A2 (n_1649));
NOR2_X1 i_1144 (.ZN (n_1093), .A1 (n_1676), .A2 (n_1644));
NOR2_X1 i_1143 (.ZN (n_1116), .A1 (n_1675), .A2 (n_1645));
NOR2_X1 i_1142 (.ZN (n_1139), .A1 (n_1674), .A2 (n_1646));
NOR2_X1 i_1141 (.ZN (n_1024), .A1 (hfn_ipo_n6), .A2 (n_1641));
NOR2_X1 i_1140 (.ZN (n_1047), .A1 (n_1678), .A2 (n_1642));
NOR2_X1 i_1139 (.ZN (n_1070), .A1 (n_1677), .A2 (n_1643));
NOR2_X1 i_1138 (.ZN (n_1232), .A1 (n_1649), .A2 (n_1669));
NOR2_X1 i_1137 (.ZN (n_1255), .A1 (n_1650), .A2 (n_1668));
NOR2_X1 i_1136 (.ZN (n_1278), .A1 (n_1651), .A2 (n_1667));
NOR2_X1 i_1135 (.ZN (n_1163), .A1 (n_1673), .A2 (n_1646));
NOR2_X1 i_1134 (.ZN (n_1186), .A1 (n_1672), .A2 (n_1647));
NOR2_X1 i_1133 (.ZN (n_1209), .A1 (n_1670), .A2 (n_1648));
NOR2_X1 i_1132 (.ZN (n_1094), .A1 (n_1676), .A2 (n_1643));
NOR2_X1 i_1131 (.ZN (n_1117), .A1 (n_1675), .A2 (n_1644));
NOR2_X1 i_1130 (.ZN (n_1140), .A1 (n_1674), .A2 (n_1645));
NOR2_X1 i_1129 (.ZN (n_1300), .A1 (n_1653), .A2 (n_1666));
NOR2_X1 i_1128 (.ZN (n_1323), .A1 (hfn_ipo_n6), .A2 (n_1665));
NOR2_X1 i_1127 (.ZN (n_1301), .A1 (n_1652), .A2 (n_1666));
NOR2_X1 i_1126 (.ZN (n_1324), .A1 (n_1653), .A2 (n_1665));
NOR2_X1 i_1125 (.ZN (n_1347), .A1 (n_1654), .A2 (n_1664));
NOR2_X1 i_1124 (.ZN (n_1025), .A1 (hfn_ipo_n6), .A2 (n_1640));
NOR2_X1 i_1123 (.ZN (n_1048), .A1 (n_1678), .A2 (n_1641));
NOR2_X1 i_1122 (.ZN (n_1071), .A1 (n_1677), .A2 (n_1642));
FA_X1 i_1121 (.CO (n_1713), .S (n_1712), .A (n_169), .B (n_167), .CI (n_461));
FA_X1 i_1120 (.CO (n_1711), .S (n_1710), .A (n_515), .B (n_509), .CI (n_517));
FA_X1 i_1119 (.CO (n_1709), .S (n_1708), .A (n_505), .B (n_504), .CI (n_507));
FA_X1 i_1118 (.CO (n_1707), .S (n_1706), .A (n_766), .B (n_519), .CI (n_533));
FA_X1 i_1117 (.CO (n_1705), .S (n_1704), .A (n_796), .B (n_535), .CI (n_798));
FA_X1 i_1116 (.CO (n_1703), .S (n_1701), .A (n_824), .B (n_799), .CI (n_826));
FA_X1 i_1115 (.CO (n_797), .S (n_796), .A (n_548), .B (n_629), .CI (n_664));
FA_X1 i_1114 (.CO (n_799), .S (n_798), .A (n_765), .B (n_794), .CI (n_767));
FA_X1 i_1113 (.CO (n_767), .S (n_766), .A (n_513), .B (n_529), .CI (n_525));
FA_X1 i_1112 (.CO (n_765), .S (n_1700), .A (n_511), .B (n_523), .CI (n_521));
FA_X1 i_1111 (.CO (n_795), .S (n_794), .A (n_545), .B (n_527), .CI (n_531));
FA_X1 i_1110 (.CO (n_1699), .S (n_1698), .A (n_850), .B (n_827), .CI (n_852));
FA_X1 i_1109 (.CO (n_827), .S (n_826), .A (n_820), .B (n_822), .CI (n_797));
FA_X1 i_1108 (.CO (n_1697), .S (n_1696), .A (n_853), .B (n_874), .CI (n_876));
FA_X1 i_1107 (.CO (n_853), .S (n_852), .A (n_823), .B (n_848), .CI (n_825));
FA_X1 i_1106 (.CO (n_825), .S (n_824), .A (n_818), .B (n_816), .CI (n_795));
FA_X1 i_1105 (.CO (n_823), .S (n_822), .A (n_547), .B (n_666), .CI (n_631));
FA_X1 i_1104 (.CO (n_901), .S (n_1695), .A (n_896), .B (n_877), .CI (n_898));
FA_X1 i_1103 (.CO (n_877), .S (n_876), .A (n_849), .B (n_872), .CI (n_851));
FA_X1 i_1102 (.CO (n_851), .S (n_850), .A (n_821), .B (n_844), .CI (n_846));
FA_X1 i_1101 (.CO (n_821), .S (n_820), .A (n_814), .B (n_812), .CI (n_549));
FA_X1 i_1100 (.CO (n_849), .S (n_848), .A (n_819), .B (n_817), .CI (n_842));
FA_X1 i_1099 (.CO (n_817), .S (n_816), .A (n_541), .B (n_810), .CI (n_808));
FA_X1 i_1098 (.CO (n_819), .S (n_818), .A (n_806), .B (n_804), .CI (n_802));
FA_X1 i_1097 (.CO (n_1694), .S (n_920), .A (n_916), .B (n_899), .CI (n_918));
FA_X1 i_1096 (.CO (n_899), .S (n_898), .A (n_892), .B (n_894), .CI (n_875));
FA_X1 i_1095 (.CO (n_875), .S (n_874), .A (n_847), .B (n_870), .CI (n_868));
FA_X1 i_1094 (.CO (n_847), .S (n_846), .A (n_830), .B (n_815), .CI (n_840));
FA_X1 i_1093 (.CO (n_815), .S (n_814), .A (n_539), .B (n_537), .CI (n_543));
FA_X1 i_1092 (.CO (n_1693), .S (n_1692), .A (n_934), .B (n_919), .CI (n_936));
FA_X1 i_1091 (.CO (n_919), .S (n_918), .A (n_914), .B (n_912), .CI (n_897));
FA_X1 i_1090 (.CO (n_897), .S (n_896), .A (n_890), .B (n_873), .CI (n_871));
FA_X1 i_1089 (.CO (n_871), .S (n_870), .A (n_858), .B (n_856), .CI (n_866));
FA_X1 i_1088 (.CO (n_873), .S (n_872), .A (n_864), .B (n_845), .CI (n_843));
FA_X1 i_1087 (.CO (n_843), .S (n_842), .A (n_803), .B (n_813), .CI (n_838));
FA_X1 i_1086 (.CO (n_813), .S (n_812), .A (n_781), .B (n_779), .CI (n_777));
FA_X1 i_1085 (.CO (n_777), .S (n_1691), .A (n_667), .B (n_668), .CI (n_669));
FA_X1 i_1084 (.CO (n_779), .S (n_1690), .A (n_702), .B (n_704), .CI (n_729));
FA_X1 i_1083 (.CO (n_781), .S (n_1688), .A (n_731), .B (n_734), .CI (n_736));
FA_X1 i_1082 (.CO (n_803), .S (n_802), .A (n_1025), .B (n_1048), .CI (n_1071));
FA_X1 i_1081 (.CO (n_845), .S (n_844), .A (n_836), .B (n_834), .CI (n_832));
FA_X1 i_1080 (.CO (n_1687), .S (n_1686), .A (n_935), .B (n_937), .CI (n_952));
FA_X1 i_1079 (.CO (n_937), .S (n_936), .A (n_915), .B (n_932), .CI (n_917));
FA_X1 i_1078 (.CO (n_917), .S (n_916), .A (n_893), .B (n_891), .CI (n_895));
FA_X1 i_1077 (.CO (n_895), .S (n_894), .A (n_867), .B (n_888), .CI (n_869));
FA_X1 i_1076 (.CO (n_869), .S (n_868), .A (n_839), .B (n_862), .CI (n_860));
FA_X1 i_1075 (.CO (n_839), .S (n_838), .A (n_1300), .B (n_1323), .CI (n_811));
FA_X1 i_1074 (.CO (n_811), .S (n_810), .A (n_1301), .B (n_1324), .CI (n_1347));
FA_X1 i_1073 (.CO (n_867), .S (n_866), .A (n_833), .B (n_831), .CI (n_841));
FA_X1 i_1072 (.CO (n_841), .S (n_840), .A (n_809), .B (n_807), .CI (n_805));
FA_X1 i_1071 (.CO (n_805), .S (n_804), .A (n_1094), .B (n_1117), .CI (n_1140));
FA_X1 i_1070 (.CO (n_807), .S (n_806), .A (n_1163), .B (n_1186), .CI (n_1209));
FA_X1 i_1069 (.CO (n_809), .S (n_808), .A (n_1232), .B (n_1255), .CI (n_1278));
FA_X1 i_1068 (.CO (n_831), .S (n_830), .A (n_1024), .B (n_1047), .CI (n_1070));
FA_X1 i_1065 (.CO (n_833), .S (n_832), .A (n_1093), .B (n_1116), .CI (n_1139));
FA_X1 i_1063 (.CO (n_891), .S (n_890), .A (n_857), .B (n_865), .CI (n_886));
FA_X1 i_1062 (.CO (n_865), .S (n_864), .A (n_1299), .B (n_837), .CI (n_835));
FA_X1 i_1061 (.CO (n_835), .S (n_834), .A (n_1162), .B (n_1185), .CI (n_1208));
FA_X1 i_1060 (.CO (n_837), .S (n_836), .A (n_1231), .B (n_1254), .CI (n_1277));
FA_X1 i_1059 (.CO (n_857), .S (n_856), .A (n_1023), .B (n_1046), .CI (n_1069));
FA_X1 i_1058 (.CO (n_893), .S (n_892), .A (n_884), .B (n_882), .CI (n_880));
FA_X1 i_1057 (.CO (n_915), .S (n_914), .A (n_904), .B (n_902), .CI (n_910));
FA_X1 i_1056 (.CO (n_935), .S (n_934), .A (n_928), .B (n_913), .CI (n_930));
FA_X1 i_1055 (.CO (n_913), .S (n_912), .A (n_889), .B (n_908), .CI (n_906));
FA_X1 i_1054 (.CO (n_889), .S (n_888), .A (n_863), .B (n_861), .CI (n_859));
FA_X1 i_1053 (.CO (n_859), .S (n_858), .A (n_1092), .B (n_1115), .CI (n_1138));
FA_X1 i_1052 (.CO (n_861), .S (n_860), .A (n_1161), .B (n_1184), .CI (n_1207));
FA_X1 i_1051 (.CO (n_863), .S (n_862), .A (n_1230), .B (n_1253), .CI (n_1276));
FA_X1 i_1050 (.CO (n_1685), .S (n_980), .A (n_976), .B (n_967), .CI (n_978));
FA_X1 i_1049 (.CO (n_1684), .S (n_978), .A (n_963), .B (n_974), .CI (n_965));
FA_X1 i_1048 (.CO (n_1683), .S (n_974), .A (n_1155), .B (n_959), .CI (n_957));
FA_X1 i_1047 (.CO (n_1682), .S (n_976), .A (n_961), .B (n_972), .CI (n_970));
FA_X1 i_1045 (.CO (n_1681), .S (n_970), .A (n_1017), .B (n_1040), .CI (n_1063));
FA_X1 i_1044 (.CO (n_1680), .S (n_972), .A (n_1086), .B (n_1109), .CI (n_1132));
FA_X1 i_1042 (.CO (n_969), .S (n_1679), .A (n_964), .B (n_966), .CI (n_953));
FA_X1 i_1041 (.CO (n_953), .S (n_952), .A (n_933), .B (n_948), .CI (n_950));
FA_X1 i_1040 (.CO (n_933), .S (n_932), .A (n_926), .B (n_924), .CI (n_922));
FA_X1 i_1039 (.CO (n_967), .S (n_966), .A (n_962), .B (n_949), .CI (n_951));
FA_X1 i_1038 (.CO (n_951), .S (n_950), .A (n_940), .B (n_931), .CI (n_946));
FA_X1 i_1037 (.CO (n_931), .S (n_930), .A (n_903), .B (n_911), .CI (n_909));
FA_X1 i_1036 (.CO (n_909), .S (n_908), .A (n_1228), .B (n_1251), .CI (n_887));
FA_X1 i_1035 (.CO (n_887), .S (n_886), .A (n_1229), .B (n_1252), .CI (n_1275));
FA_X1 i_1034 (.CO (n_911), .S (n_910), .A (n_885), .B (n_883), .CI (n_881));
FA_X1 i_1033 (.CO (n_881), .S (n_880), .A (n_1022), .B (n_1045), .CI (n_1068));
FA_X1 i_1032 (.CO (n_883), .S (n_882), .A (n_1091), .B (n_1114), .CI (n_1137));
FA_X1 i_1031 (.CO (n_885), .S (n_884), .A (n_1160), .B (n_1183), .CI (n_1206));
FA_X1 i_1030 (.CO (n_903), .S (n_902), .A (n_1021), .B (n_1044), .CI (n_1067));
FA_X1 i_1029 (.CO (n_949), .S (n_948), .A (n_929), .B (n_944), .CI (n_942));
FA_X1 i_1028 (.CO (n_929), .S (n_928), .A (n_1227), .B (n_907), .CI (n_905));
FA_X1 i_1027 (.CO (n_905), .S (n_904), .A (n_1090), .B (n_1113), .CI (n_1136));
FA_X1 i_1026 (.CO (n_907), .S (n_906), .A (n_1159), .B (n_1182), .CI (n_1205));
FA_X1 i_1025 (.CO (n_963), .S (n_962), .A (n_943), .B (n_941), .CI (n_947));
FA_X1 i_1024 (.CO (n_947), .S (n_946), .A (n_927), .B (n_925), .CI (n_923));
FA_X1 i_1022 (.CO (n_923), .S (n_922), .A (n_1020), .B (n_1043), .CI (n_1066));
FA_X1 i_1019 (.CO (n_925), .S (n_924), .A (n_1089), .B (n_1112), .CI (n_1135));
FA_X1 i_1018 (.CO (n_927), .S (n_926), .A (n_1158), .B (n_1181), .CI (n_1204));
FA_X1 i_1017 (.CO (n_941), .S (n_940), .A (n_1019), .B (n_1042), .CI (n_1065));
FA_X1 i_1016 (.CO (n_943), .S (n_942), .A (n_1088), .B (n_1111), .CI (n_1134));
FA_X1 i_1015 (.CO (n_965), .S (n_964), .A (n_960), .B (n_958), .CI (n_956));
FA_X1 i_1014 (.CO (n_957), .S (n_956), .A (n_1018), .B (n_1041), .CI (n_1064));
FA_X1 i_1013 (.CO (n_959), .S (n_958), .A (n_1087), .B (n_1110), .CI (n_1133));
FA_X1 i_1012 (.CO (n_961), .S (n_960), .A (n_1156), .B (n_1179), .CI (n_945));
FA_X1 i_1011 (.CO (n_945), .S (n_944), .A (n_1157), .B (n_1180), .CI (n_1203));
INV_X2 i_1010 (.ZN (n_1678), .A (B_imm[22]));
INV_X2 i_1009 (.ZN (n_1677), .A (B_imm[21]));
INV_X2 i_1008 (.ZN (n_1676), .A (B_imm[20]));
INV_X4 i_1007 (.ZN (n_1675), .A (B_imm[19]));
INV_X4 i_1006 (.ZN (n_1674), .A (B_imm[18]));
INV_X4 i_1005 (.ZN (n_1673), .A (B_imm[17]));
INV_X4 i_1004 (.ZN (n_1672), .A (B_imm[16]));
INV_X4 i_1003 (.ZN (n_1670), .A (B_imm[15]));
INV_X4 i_1002 (.ZN (n_1669), .A (B_imm[14]));
INV_X4 i_1001 (.ZN (n_1668), .A (B_imm[13]));
INV_X4 i_999 (.ZN (n_1667), .A (B_imm[12]));
INV_X4 i_996 (.ZN (n_1666), .A (B_imm[11]));
INV_X4 i_995 (.ZN (n_1665), .A (B_imm[10]));
INV_X4 i_994 (.ZN (n_1664), .A (B_imm[9]));
INV_X4 i_993 (.ZN (n_1663), .A (B_imm[8]));
INV_X4 i_992 (.ZN (n_1662), .A (B_imm[7]));
INV_X4 i_991 (.ZN (n_1661), .A (B_imm[6]));
INV_X2 i_990 (.ZN (n_1660), .A (B_imm[5]));
INV_X2 i_989 (.ZN (n_1659), .A (B_imm[4]));
INV_X2 i_988 (.ZN (n_1658), .A (B_imm[3]));
INV_X2 i_987 (.ZN (n_1657), .A (B_imm[2]));
INV_X2 i_986 (.ZN (n_1656), .A (B_imm[1]));
INV_X2 i_985 (.ZN (n_1655), .A (B_imm[0]));
INV_X1 i_984 (.ZN (n_1654), .A (A_imm[23]));
INV_X2 i_983 (.ZN (n_1653), .A (A_imm[22]));
INV_X2 i_982 (.ZN (n_1652), .A (A_imm[21]));
INV_X4 i_981 (.ZN (n_1651), .A (A_imm[20]));
INV_X4 i_980 (.ZN (n_1650), .A (A_imm[19]));
INV_X4 i_979 (.ZN (n_1649), .A (A_imm[18]));
INV_X2 i_978 (.ZN (n_1648), .A (A_imm[17]));
INV_X4 i_973 (.ZN (n_1647), .A (A_imm[16]));
INV_X2 i_972 (.ZN (n_1646), .A (A_imm[15]));
INV_X2 i_971 (.ZN (n_1645), .A (A_imm[14]));
INV_X4 i_970 (.ZN (n_1644), .A (A_imm[13]));
INV_X2 i_969 (.ZN (n_1643), .A (A_imm[12]));
INV_X4 i_968 (.ZN (n_1642), .A (A_imm[11]));
INV_X4 i_967 (.ZN (n_1641), .A (A_imm[10]));
INV_X4 i_966 (.ZN (n_1640), .A (A_imm[9]));
INV_X4 i_965 (.ZN (n_1639), .A (A_imm[8]));
INV_X8 i_964 (.ZN (n_1634), .A (A_imm[7]));
INV_X8 i_963 (.ZN (n_1633), .A (A_imm[6]));
INV_X4 i_962 (.ZN (n_1632), .A (A_imm[5]));
INV_X8 i_961 (.ZN (n_1631), .A (A_imm[4]));
INV_X8 i_960 (.ZN (n_1630), .A (A_imm[3]));
INV_X4 i_959 (.ZN (n_1629), .A (A_imm[2]));
INV_X4 i_958 (.ZN (n_1628), .A (A_imm[1]));
INV_X4 i_957 (.ZN (n_1625), .A (A_imm[0]));
INV_X1 i_956 (.ZN (n_1623), .A (n_763));
INV_X1 i_955 (.ZN (n_1622), .A (n_418));
INV_X1 i_950 (.ZN (n_1621), .A (n_340));
INV_X1 i_949 (.ZN (n_1619), .A (n_379));
INV_X1 i_948 (.ZN (n_1608), .A (n_305));
NOR2_X1 i_947 (.ZN (n_1586), .A1 (n_775), .A2 (n_900));
NAND2_X1 i_946 (.ZN (n_1585), .A1 (n_773), .A2 (n_938));
INV_X1 i_945 (.ZN (n_1584), .A (n_1585));
NOR2_X1 i_944 (.ZN (n_1583), .A1 (n_460), .A2 (n_419));
NAND2_X1 i_943 (.ZN (n_1569), .A1 (n_460), .A2 (n_419));
NAND2_X1 i_942 (.ZN (n_1536), .A1 (n_1622), .A2 (n_1619));
NOR2_X1 i_941 (.ZN (n_1513), .A1 (n_1622), .A2 (n_1619));
AOI22_X1 i_940 (.ZN (n_1490), .A1 (n_52), .A2 (n_54), .B1 (n_38), .B2 (n_40));
AOI22_X1 i_939 (.ZN (n_1348), .A1 (n_16), .A2 (n_18), .B1 (n_26), .B2 (n_28));
AOI21_X1 i_938 (.ZN (n_1325), .A (n_1623), .B1 (n_954), .B2 (n_955));
NOR2_X1 i_937 (.ZN (n_1302), .A1 (n_16), .A2 (n_18));
OAI21_X1 i_936 (.ZN (n_1279), .A (n_1348), .B1 (n_1325), .B2 (n_1302));
OAI221_X1 i_935 (.ZN (n_1272), .A (n_1279), .B1 (n_26), .B2 (n_28), .C1 (n_38), .C2 (n_40));
OAI222_X1 i_934 (.ZN (n_1256), .A1 (n_86), .A2 (n_88), .B1 (n_106), .B2 (n_108), .C1 (n_128), .C2 (n_130));
OAI22_X1 i_933 (.ZN (n_1249), .A1 (n_68), .A2 (n_70), .B1 (n_52), .B2 (n_54));
AOI211_X1 i_932 (.ZN (n_1233), .A (n_1256), .B (n_1249), .C1 (n_1490), .C2 (n_1272));
AOI22_X1 i_927 (.ZN (n_1226), .A1 (n_68), .A2 (n_70), .B1 (n_86), .B2 (n_88));
OAI211_X1 i_926 (.ZN (n_1210), .A (n_106), .B (n_108), .C1 (n_128), .C2 (n_130));
AOI21_X1 i_925 (.ZN (n_1187), .A (n_1233), .B1 (n_128), .B2 (n_130));
OAI211_X1 i_924 (.ZN (n_1164), .A (n_1210), .B (n_1187), .C1 (n_1256), .C2 (n_1226));
NOR2_X1 i_923 (.ZN (n_1011), .A1 (n_236), .A2 (n_238));
OAI222_X1 i_922 (.ZN (n_1010), .A1 (n_178), .A2 (n_180), .B1 (n_206), .B2 (n_208)
    , .C1 (n_236), .C2 (n_238));
INV_X1 i_921 (.ZN (n_1009), .A (n_1010));
OAI211_X1 i_920 (.ZN (n_1008), .A (n_1009), .B (n_1164), .C1 (n_152), .C2 (n_154));
AOI22_X1 i_919 (.ZN (n_1007), .A1 (n_152), .A2 (n_154), .B1 (n_178), .B2 (n_180));
AOI22_X1 i_918 (.ZN (n_1005), .A1 (n_236), .A2 (n_238), .B1 (n_206), .B2 (n_208));
OAI221_X1 i_917 (.ZN (n_998), .A (n_1008), .B1 (n_1010), .B2 (n_1007), .C1 (n_1011), .C2 (n_1005));
NOR2_X1 i_916 (.ZN (n_991), .A1 (n_304), .A2 (n_271));
NOR2_X2 i_915 (.ZN (n_990), .A1 (n_376), .A2 (n_378));
AOI211_X2 i_914 (.ZN (n_989), .A (n_991), .B (n_990), .C1 (n_1621), .C2 (n_1608));
OAI211_X2 i_913 (.ZN (n_987), .A (n_998), .B (n_989), .C1 (n_268), .C2 (n_270));
AOI22_X1 i_912 (.ZN (n_985), .A1 (n_268), .A2 (n_270), .B1 (n_304), .B2 (n_271));
INV_X1 i_911 (.ZN (n_983), .A (n_985));
NOR3_X1 i_910 (.ZN (n_981), .A1 (n_1621), .A2 (n_990), .A3 (n_1608));
AOI221_X2 i_909 (.ZN (n_979), .A (n_981), .B1 (n_989), .B2 (n_983), .C1 (n_376), .C2 (n_378));
NAND2_X1 i_904 (.ZN (n_977), .A1 (n_987), .A2 (n_979));
OAI21_X1 i_903 (.ZN (n_975), .A (n_1536), .B1 (n_1513), .B2 (n_977));
AOI21_X1 i_902 (.ZN (n_973), .A (n_1583), .B1 (n_1569), .B2 (n_975));
AOI21_X1 i_901 (.ZN (n_971), .A (n_1586), .B1 (n_775), .B2 (n_900));
OAI22_X1 i_900 (.ZN (n_968), .A1 (n_773), .A2 (n_938), .B1 (n_1584), .B2 (n_973));
XNOR2_X1 i_899 (.ZN (Res_imm[24]), .A (n_971), .B (n_968));
NOR2_X1 i_898 (.ZN (n_1451), .A1 (n_1660), .A2 (n_1646));
NOR2_X1 i_897 (.ZN (n_1474), .A1 (n_1659), .A2 (n_1647));
NOR2_X1 i_896 (.ZN (n_1497), .A1 (n_1658), .A2 (n_1648));
NOR2_X1 i_895 (.ZN (n_1382), .A1 (n_1663), .A2 (n_1643));
NOR2_X1 i_894 (.ZN (n_1405), .A1 (n_1662), .A2 (n_1644));
NOR2_X1 i_893 (.ZN (n_1428), .A1 (n_1661), .A2 (n_1645));
NOR2_X1 i_892 (.ZN (n_1313), .A1 (n_1666), .A2 (n_1640));
NOR2_X1 i_891 (.ZN (n_1336), .A1 (n_1665), .A2 (n_1641));
NOR2_X1 i_890 (.ZN (n_1359), .A1 (n_1664), .A2 (n_1642));
NOR2_X1 i_889 (.ZN (n_1430), .A1 (n_1661), .A2 (n_1643));
NOR2_X1 i_888 (.ZN (n_1453), .A1 (n_1660), .A2 (n_1644));
NOR2_X1 i_887 (.ZN (n_1476), .A1 (n_1659), .A2 (n_1645));
NOR2_X1 i_886 (.ZN (n_1361), .A1 (n_1664), .A2 (n_1640));
NOR2_X1 i_881 (.ZN (n_1384), .A1 (n_1663), .A2 (n_1641));
NOR2_X1 i_880 (.ZN (n_1407), .A1 (n_1662), .A2 (n_1642));
NOR2_X1 i_879 (.ZN (n_1292), .A1 (n_1667), .A2 (n_1633));
NOR2_X1 i_878 (.ZN (n_1315), .A1 (n_1666), .A2 (n_1634));
NOR2_X1 i_877 (.ZN (n_1338), .A1 (n_1665), .A2 (n_1639));
NOR2_X1 i_876 (.ZN (n_1544), .A1 (n_1656), .A2 (n_1649));
NOR2_X1 i_875 (.ZN (n_1565), .A1 (n_1655), .A2 (n_1650));
NOR2_X1 i_874 (.ZN (n_1499), .A1 (n_1658), .A2 (n_1646));
NOR2_X1 i_873 (.ZN (n_1522), .A1 (n_1657), .A2 (n_1647));
NOR2_X1 i_872 (.ZN (n_1545), .A1 (n_1656), .A2 (n_1648));
NOR2_X1 i_871 (.ZN (n_1520), .A1 (n_1657), .A2 (n_1649));
NOR2_X1 i_870 (.ZN (n_1543), .A1 (n_1656), .A2 (n_1650));
NOR2_X1 i_869 (.ZN (n_1564), .A1 (n_1655), .A2 (n_1651));
NOR2_X1 i_868 (.ZN (n_1223), .A1 (n_1670), .A2 (n_1630));
NOR2_X1 i_867 (.ZN (n_1246), .A1 (n_1669), .A2 (n_1631));
NOR2_X1 i_866 (.ZN (n_1269), .A1 (n_1668), .A2 (n_1632));
NOR2_X1 i_865 (.ZN (n_1154), .A1 (n_1674), .A2 (n_1625));
NOR2_X1 i_864 (.ZN (n_1177), .A1 (n_1673), .A2 (n_1628));
NOR2_X1 i_863 (.ZN (n_1200), .A1 (n_1672), .A2 (n_1629));
NOR2_X2 i_858 (.ZN (n_1385), .A1 (n_1663), .A2 (n_1640));
NOR2_X1 i_857 (.ZN (n_1408), .A1 (n_1662), .A2 (n_1641));
NOR2_X1 i_856 (.ZN (n_1431), .A1 (n_1661), .A2 (n_1642));
NOR2_X1 i_855 (.ZN (n_1316), .A1 (n_1666), .A2 (n_1633));
NOR2_X1 i_854 (.ZN (n_1339), .A1 (n_1665), .A2 (n_1634));
NOR2_X1 i_853 (.ZN (n_1362), .A1 (n_1664), .A2 (n_1639));
NOR2_X1 i_852 (.ZN (n_1247), .A1 (n_1669), .A2 (n_1630));
NOR2_X1 i_851 (.ZN (n_1270), .A1 (n_1668), .A2 (n_1631));
NOR2_X1 i_850 (.ZN (n_1293), .A1 (n_1667), .A2 (n_1632));
NOR2_X1 i_849 (.ZN (n_1268), .A1 (n_1668), .A2 (n_1633));
NOR2_X1 i_848 (.ZN (n_1291), .A1 (n_1667), .A2 (n_1634));
NOR2_X1 i_847 (.ZN (n_1314), .A1 (n_1666), .A2 (n_1639));
NOR2_X1 i_846 (.ZN (n_1199), .A1 (n_1672), .A2 (n_1630));
NOR2_X2 i_845 (.ZN (n_1222), .A1 (n_1670), .A2 (n_1631));
NOR2_X1 i_844 (.ZN (n_1245), .A1 (n_1669), .A2 (n_1632));
NOR2_X1 i_843 (.ZN (n_1130), .A1 (n_1675), .A2 (n_1625));
NOR2_X1 i_842 (.ZN (n_1153), .A1 (n_1674), .A2 (n_1628));
NOR2_X1 i_841 (.ZN (n_1176), .A1 (n_1673), .A2 (n_1629));
NOR2_X1 i_840 (.ZN (n_1475), .A1 (n_1659), .A2 (n_1646));
NOR2_X1 i_835 (.ZN (n_1498), .A1 (n_1658), .A2 (n_1647));
NOR2_X1 i_834 (.ZN (n_1521), .A1 (n_1657), .A2 (n_1648));
NOR2_X1 i_833 (.ZN (n_1406), .A1 (n_1662), .A2 (n_1643));
NOR2_X1 i_832 (.ZN (n_1429), .A1 (n_1661), .A2 (n_1644));
NOR2_X1 i_831 (.ZN (n_1452), .A1 (n_1660), .A2 (n_1645));
NOR2_X1 i_830 (.ZN (n_1337), .A1 (n_1665), .A2 (n_1640));
NOR2_X1 i_829 (.ZN (n_1360), .A1 (n_1664), .A2 (n_1641));
NOR2_X1 i_828 (.ZN (n_1383), .A1 (n_1663), .A2 (n_1642));
NOR2_X1 i_827 (.ZN (n_1427), .A1 (n_1661), .A2 (n_1646));
NOR2_X1 i_826 (.ZN (n_1450), .A1 (n_1660), .A2 (n_1647));
NOR2_X1 i_825 (.ZN (n_1473), .A1 (n_1659), .A2 (n_1648));
NOR2_X1 i_824 (.ZN (n_1358), .A1 (n_1664), .A2 (n_1643));
NOR2_X1 i_823 (.ZN (n_1381), .A1 (n_1663), .A2 (n_1644));
NOR2_X1 i_822 (.ZN (n_1404), .A1 (n_1662), .A2 (n_1645));
NOR2_X1 i_821 (.ZN (n_1289), .A1 (n_1667), .A2 (n_1640));
NOR2_X1 i_820 (.ZN (n_1312), .A1 (n_1666), .A2 (n_1641));
NOR2_X1 i_819 (.ZN (n_1335), .A1 (n_1665), .A2 (n_1642));
NOR2_X1 i_818 (.ZN (n_1220), .A1 (n_1670), .A2 (n_1633));
NOR2_X1 i_817 (.ZN (n_1243), .A1 (n_1669), .A2 (n_1634));
NOR2_X1 i_814 (.ZN (n_1266), .A1 (n_1668), .A2 (n_1639));
NOR2_X1 i_812 (.ZN (n_1496), .A1 (n_1658), .A2 (n_1649));
NOR2_X1 i_811 (.ZN (n_1519), .A1 (n_1657), .A2 (n_1650));
NOR2_X1 i_810 (.ZN (n_1542), .A1 (n_1656), .A2 (n_1651));
NOR2_X1 i_809 (.ZN (n_1151), .A1 (n_1674), .A2 (n_1630));
NOR2_X1 i_808 (.ZN (n_1174), .A1 (n_1673), .A2 (n_1631));
NOR2_X1 i_807 (.ZN (n_1197), .A1 (n_1672), .A2 (n_1632));
NOR2_X1 i_806 (.ZN (n_1082), .A1 (n_1677), .A2 (n_1625));
NOR2_X1 i_805 (.ZN (n_1105), .A1 (n_1676), .A2 (n_1628));
NOR2_X1 i_804 (.ZN (n_1128), .A1 (n_1675), .A2 (n_1629));
NOR2_X1 i_803 (.ZN (n_1175), .A1 (n_1673), .A2 (n_1630));
NOR2_X1 i_802 (.ZN (n_1198), .A1 (n_1672), .A2 (n_1631));
NOR2_X1 i_801 (.ZN (n_1221), .A1 (n_1670), .A2 (n_1632));
NOR2_X1 i_800 (.ZN (n_1106), .A1 (n_1676), .A2 (n_1625));
NOR2_X1 i_799 (.ZN (n_1129), .A1 (n_1675), .A2 (n_1628));
NOR2_X1 i_798 (.ZN (n_1152), .A1 (n_1674), .A2 (n_1629));
NOR2_X1 i_797 (.ZN (n_1178), .A1 (n_1673), .A2 (n_1625));
NOR2_X1 i_796 (.ZN (n_1201), .A1 (n_1672), .A2 (n_1628));
NOR2_X1 i_795 (.ZN (n_1224), .A1 (n_1670), .A2 (n_1629));
NOR2_X1 i_794 (.ZN (n_1478), .A1 (n_1659), .A2 (n_1643));
NOR2_X1 i_793 (.ZN (n_1501), .A1 (n_1658), .A2 (n_1644));
NOR2_X1 i_791 (.ZN (n_1524), .A1 (n_1657), .A2 (n_1645));
NOR2_X1 i_789 (.ZN (n_1409), .A1 (n_1662), .A2 (n_1640));
NOR2_X1 i_788 (.ZN (n_1432), .A1 (n_1661), .A2 (n_1641));
NOR2_X1 i_787 (.ZN (n_1455), .A1 (n_1660), .A2 (n_1642));
NOR2_X1 i_786 (.ZN (n_1340), .A1 (n_1665), .A2 (n_1633));
NOR2_X1 i_785 (.ZN (n_1363), .A1 (n_1664), .A2 (n_1634));
NOR2_X1 i_784 (.ZN (n_1386), .A1 (n_1663), .A2 (n_1639));
NOR2_X1 i_783 (.ZN (n_1244), .A1 (n_1669), .A2 (n_1633));
NOR2_X1 i_782 (.ZN (n_1267), .A1 (n_1668), .A2 (n_1634));
NOR2_X1 i_781 (.ZN (n_1290), .A1 (n_1667), .A2 (n_1639));
NOR2_X1 i_780 (.ZN (n_1566), .A1 (n_1655), .A2 (n_1649));
NOR2_X1 i_779 (.ZN (n_1523), .A1 (n_1657), .A2 (n_1646));
NOR2_X1 i_778 (.ZN (n_1546), .A1 (n_1656), .A2 (n_1647));
NOR2_X1 i_777 (.ZN (n_1567), .A1 (n_1655), .A2 (n_1648));
NOR2_X1 i_776 (.ZN (n_1454), .A1 (n_1660), .A2 (n_1643));
NOR2_X1 i_775 (.ZN (n_1477), .A1 (n_1659), .A2 (n_1644));
NOR2_X1 i_774 (.ZN (n_1500), .A1 (n_1658), .A2 (n_1645));
NOR2_X1 i_773 (.ZN (n_1563), .A1 (n_1655), .A2 (n_1652));
NOR2_X1 i_772 (.ZN (n_1541), .A1 (n_1656), .A2 (n_1652));
NOR2_X1 i_771 (.ZN (n_1562), .A1 (n_1655), .A2 (n_1653));
NOR2_X1 i_770 (.ZN (n_1265), .A1 (n_1668), .A2 (n_1640));
NOR2_X1 i_769 (.ZN (n_1288), .A1 (n_1667), .A2 (n_1641));
NOR2_X1 i_768 (.ZN (n_1311), .A1 (n_1666), .A2 (n_1642));
NOR2_X1 i_766 (.ZN (n_1196), .A1 (n_1672), .A2 (n_1633));
NOR2_X1 i_765 (.ZN (n_1219), .A1 (n_1670), .A2 (n_1634));
NOR2_X1 i_764 (.ZN (n_1242), .A1 (n_1669), .A2 (n_1639));
NOR2_X1 i_763 (.ZN (n_1127), .A1 (n_1675), .A2 (n_1630));
NOR2_X1 i_762 (.ZN (n_1150), .A1 (n_1674), .A2 (n_1631));
NOR2_X1 i_761 (.ZN (n_1173), .A1 (n_1673), .A2 (n_1632));
NOR2_X1 i_760 (.ZN (n_1472), .A1 (n_1659), .A2 (n_1649));
NOR2_X1 i_759 (.ZN (n_1495), .A1 (n_1658), .A2 (n_1650));
NOR2_X1 i_758 (.ZN (n_1518), .A1 (n_1657), .A2 (n_1651));
NOR2_X1 i_757 (.ZN (n_1403), .A1 (n_1662), .A2 (n_1646));
NOR2_X1 i_756 (.ZN (n_1426), .A1 (n_1661), .A2 (n_1647));
NOR2_X1 i_755 (.ZN (n_1449), .A1 (n_1660), .A2 (n_1648));
NOR2_X1 i_754 (.ZN (n_1334), .A1 (n_1665), .A2 (n_1643));
NOR2_X1 i_753 (.ZN (n_1357), .A1 (n_1664), .A2 (n_1644));
NOR2_X1 i_752 (.ZN (n_1380), .A1 (n_1663), .A2 (n_1645));
NOR2_X1 i_751 (.ZN (n_1058), .A1 (n_1678), .A2 (n_1625));
NOR2_X1 i_750 (.ZN (n_1081), .A1 (n_1677), .A2 (n_1628));
NOR2_X1 i_749 (.ZN (n_1104), .A1 (n_1676), .A2 (n_1629));
NOR2_X1 i_748 (.ZN (n_1172), .A1 (n_1673), .A2 (n_1633));
NOR2_X1 i_747 (.ZN (n_1195), .A1 (n_1672), .A2 (n_1634));
NOR2_X1 i_746 (.ZN (n_1218), .A1 (n_1670), .A2 (n_1639));
NOR2_X1 i_745 (.ZN (n_1103), .A1 (n_1676), .A2 (n_1630));
NOR2_X1 i_743 (.ZN (n_1126), .A1 (n_1675), .A2 (n_1631));
NOR2_X1 i_742 (.ZN (n_1149), .A1 (n_1674), .A2 (n_1632));
NOR2_X1 i_741 (.ZN (n_1034), .A1 (n_1654), .A2 (n_1625));
NOR2_X1 i_740 (.ZN (n_1057), .A1 (n_1678), .A2 (n_1628));
NOR2_X1 i_739 (.ZN (n_1080), .A1 (n_1677), .A2 (n_1629));
NOR2_X1 i_738 (.ZN (n_1379), .A1 (n_1663), .A2 (n_1646));
NOR2_X1 i_737 (.ZN (n_1402), .A1 (n_1662), .A2 (n_1647));
NOR2_X1 i_736 (.ZN (n_1425), .A1 (n_1661), .A2 (n_1648));
NOR2_X1 i_735 (.ZN (n_1310), .A1 (n_1666), .A2 (n_1643));
NOR2_X1 i_734 (.ZN (n_1333), .A1 (n_1665), .A2 (n_1644));
NOR2_X1 i_733 (.ZN (n_1356), .A1 (n_1664), .A2 (n_1645));
NOR2_X1 i_732 (.ZN (n_1241), .A1 (n_1669), .A2 (n_1640));
NOR2_X1 i_731 (.ZN (n_1264), .A1 (n_1668), .A2 (n_1641));
NOR2_X1 i_730 (.ZN (n_1287), .A1 (n_1667), .A2 (n_1642));
NOR2_X1 i_729 (.ZN (n_1517), .A1 (n_1657), .A2 (n_1652));
NOR2_X1 i_728 (.ZN (n_1540), .A1 (n_1656), .A2 (n_1653));
NOR2_X1 i_727 (.ZN (n_1561), .A1 (n_1655), .A2 (n_1654));
NOR2_X1 i_726 (.ZN (n_1448), .A1 (n_1660), .A2 (n_1649));
NOR2_X1 i_725 (.ZN (n_1471), .A1 (n_1659), .A2 (n_1650));
NOR2_X1 i_724 (.ZN (n_1494), .A1 (n_1658), .A2 (n_1651));
NOR2_X1 i_723 (.ZN (n_1102), .A1 (n_1676), .A2 (n_1631));
NOR2_X1 i_722 (.ZN (n_1125), .A1 (n_1675), .A2 (n_1632));
NOR2_X1 i_721 (.ZN (n_1148), .A1 (n_1674), .A2 (n_1633));
NOR2_X1 i_720 (.ZN (n_1033), .A1 (n_1654), .A2 (n_1628));
NOR2_X1 i_719 (.ZN (n_1056), .A1 (n_1678), .A2 (n_1629));
NOR2_X1 i_718 (.ZN (n_1079), .A1 (n_1677), .A2 (n_1630));
NOR2_X1 i_717 (.ZN (n_1309), .A1 (n_1666), .A2 (n_1644));
NOR2_X1 i_716 (.ZN (n_1332), .A1 (n_1665), .A2 (n_1645));
NOR2_X1 i_715 (.ZN (n_1355), .A1 (n_1664), .A2 (n_1646));
NOR2_X1 i_714 (.ZN (n_1240), .A1 (n_1669), .A2 (n_1641));
NOR2_X1 i_713 (.ZN (n_1263), .A1 (n_1668), .A2 (n_1642));
NOR2_X1 i_712 (.ZN (n_1286), .A1 (n_1667), .A2 (n_1643));
NOR2_X1 i_711 (.ZN (n_1171), .A1 (n_1673), .A2 (n_1634));
NOR2_X1 i_710 (.ZN (n_1194), .A1 (n_1672), .A2 (n_1639));
NOR2_X1 i_709 (.ZN (n_1217), .A1 (n_1670), .A2 (n_1640));
NOR2_X1 i_708 (.ZN (n_1516), .A1 (n_1657), .A2 (n_1653));
NOR2_X1 i_707 (.ZN (n_1539), .A1 (n_1656), .A2 (n_1654));
NOR2_X1 i_706 (.ZN (n_1447), .A1 (n_1660), .A2 (n_1650));
NOR2_X1 i_705 (.ZN (n_1470), .A1 (n_1659), .A2 (n_1651));
NOR2_X1 i_704 (.ZN (n_1493), .A1 (n_1658), .A2 (n_1652));
NOR2_X1 i_703 (.ZN (n_1378), .A1 (n_1663), .A2 (n_1647));
NOR2_X1 i_702 (.ZN (n_1401), .A1 (n_1662), .A2 (n_1648));
NOR2_X1 i_701 (.ZN (n_1424), .A1 (n_1661), .A2 (n_1649));
NOR2_X1 i_700 (.ZN (n_1271), .A1 (n_1668), .A2 (n_1630));
NOR2_X1 i_699 (.ZN (n_1294), .A1 (n_1667), .A2 (n_1631));
NOR2_X1 i_698 (.ZN (n_1317), .A1 (n_1666), .A2 (n_1632));
NOR2_X1 i_697 (.ZN (n_1202), .A1 (n_1672), .A2 (n_1625));
NOR2_X1 i_696 (.ZN (n_1225), .A1 (n_1670), .A2 (n_1628));
NOR2_X1 i_695 (.ZN (n_1248), .A1 (n_1669), .A2 (n_1629));
NOR2_X1 i_694 (.ZN (n_1433), .A1 (n_1661), .A2 (n_1640));
NOR2_X1 i_693 (.ZN (n_1456), .A1 (n_1660), .A2 (n_1641));
NOR2_X1 i_692 (.ZN (n_1479), .A1 (n_1659), .A2 (n_1642));
NOR2_X1 i_691 (.ZN (n_1364), .A1 (n_1664), .A2 (n_1633));
NOR2_X1 i_690 (.ZN (n_1387), .A1 (n_1663), .A2 (n_1634));
NOR2_X1 i_689 (.ZN (n_1410), .A1 (n_1662), .A2 (n_1639));
NOR2_X1 i_688 (.ZN (n_1295), .A1 (n_1667), .A2 (n_1630));
NOR2_X1 i_687 (.ZN (n_1318), .A1 (n_1666), .A2 (n_1631));
NOR2_X1 i_686 (.ZN (n_1341), .A1 (n_1665), .A2 (n_1632));
NOR2_X1 i_685 (.ZN (n_1547), .A1 (n_1656), .A2 (n_1646));
NOR2_X1 i_684 (.ZN (n_1568), .A1 (n_1655), .A2 (n_1647));
NOR2_X1 i_683 (.ZN (n_1502), .A1 (n_1658), .A2 (n_1643));
NOR2_X1 i_682 (.ZN (n_1525), .A1 (n_1657), .A2 (n_1644));
NOR2_X1 i_681 (.ZN (n_1548), .A1 (n_1656), .A2 (n_1645));
HA_X1 i_680 (.CO (n_11), .S (n_955), .A (n_3), .B (n_6));
FA_X1 i_679 (.CO (n_7), .S (n_954), .A (n_737), .B (n_738), .CI (n_739));
HA_X1 i_678 (.CO (n_19), .S (n_18), .A (n_9), .B (n_11));
FA_X1 i_677 (.CO (n_17), .S (n_16), .A (n_7), .B (n_8), .CI (n_10));
HA_X1 i_676 (.CO (n_29), .S (n_28), .A (n_19), .B (n_17));
FA_X1 i_675 (.CO (n_27), .S (n_26), .A (n_14), .B (n_12), .CI (n_20));
HA_X1 i_674 (.CO (n_55), .S (n_54), .A (n_39), .B (n_37));
FA_X1 i_673 (.CO (n_53), .S (n_52), .A (n_36), .B (n_32), .CI (n_41));
HA_X1 i_672 (.CO (n_41), .S (n_40), .A (n_30), .B (n_27));
FA_X1 i_671 (.CO (n_39), .S (n_38), .A (n_24), .B (n_22), .CI (n_29));
HA_X1 i_670 (.CO (n_71), .S (n_70), .A (n_55), .B (n_53));
FA_X1 i_669 (.CO (n_69), .S (n_68), .A (n_48), .B (n_50), .CI (n_51));
HA_X1 i_668 (.CO (n_89), .S (n_88), .A (n_71), .B (n_69));
FA_X1 i_667 (.CO (n_87), .S (n_86), .A (n_64), .B (n_79), .CI (n_82));
HA_X1 i_666 (.CO (n_131), .S (n_130), .A (n_107), .B (n_109));
HA_X1 i_665 (.CO (n_109), .S (n_108), .A (n_89), .B (n_87));
FA_X1 i_664 (.CO (n_107), .S (n_106), .A (n_102), .B (n_100), .CI (n_104));
FA_X1 i_663 (.CO (n_145), .S (n_144), .A (n_116), .B (n_136), .CI (n_134));
FA_X1 i_662 (.CO (n_147), .S (n_146), .A (n_132), .B (n_119), .CI (n_118));
FA_X1 i_661 (.CO (n_129), .S (n_128), .A (n_105), .B (n_124), .CI (n_126));
FA_X1 i_660 (.CO (n_125), .S (n_124), .A (n_98), .B (n_120), .CI (n_115));
FA_X1 i_659 (.CO (n_105), .S (n_104), .A (n_94), .B (n_81), .CI (n_83));
FA_X1 i_658 (.CO (n_127), .S (n_126), .A (n_101), .B (n_103), .CI (n_122));
FA_X1 i_657 (.CO (n_103), .S (n_102), .A (n_90), .B (n_84), .CI (n_67));
FA_X1 i_656 (.CO (n_101), .S (n_100), .A (n_66), .B (n_93), .CI (n_92));
FA_X1 i_655 (.CO (n_123), .S (n_122), .A (n_114), .B (n_112), .CI (n_110));
FA_X1 i_654 (.CO (n_939), .S (n_142), .A (n_113), .B (n_111), .CI (n_99));
FA_X1 i_653 (.CO (n_121), .S (n_120), .A (n_91), .B (n_85), .CI (n_96));
HA_X1 i_652 (.CO (n_181), .S (n_180), .A (n_153), .B (n_155));
HA_X1 i_651 (.CO (n_155), .S (n_154), .A (n_150), .B (n_131));
FA_X1 i_650 (.CO (n_153), .S (n_152), .A (n_148), .B (n_127), .CI (n_129));
FA_X1 i_649 (.CO (n_179), .S (n_178), .A (n_174), .B (n_151), .CI (n_176));
FA_X1 i_648 (.CO (n_151), .S (n_150), .A (n_125), .B (n_146), .CI (n_144));
FA_X1 i_647 (.CO (n_201), .S (n_200), .A (n_166), .B (n_194), .CI (n_192));
FA_X1 i_646 (.CO (n_175), .S (n_174), .A (n_147), .B (n_145), .CI (n_165));
FA_X1 i_645 (.CO (n_197), .S (n_196), .A (n_164), .B (n_190), .CI (n_188));
FA_X1 i_644 (.CO (n_203), .S (n_202), .A (n_171), .B (n_173), .CI (n_198));
FA_X1 i_643 (.CO (n_199), .S (n_198), .A (n_186), .B (n_184), .CI (n_182));
FA_X1 i_642 (.CO (n_177), .S (n_176), .A (n_149), .B (n_172), .CI (n_170));
FA_X1 i_641 (.CO (n_171), .S (n_170), .A (n_161), .B (n_159), .CI (n_157));
FA_X1 i_640 (.CO (n_173), .S (n_172), .A (n_143), .B (n_138), .CI (n_163));
FA_X1 i_639 (.CO (n_149), .S (n_148), .A (n_121), .B (n_142), .CI (n_123));
HA_X1 i_638 (.CO (n_271), .S (n_270), .A (n_237), .B (n_239));
HA_X1 i_637 (.CO (n_239), .S (n_238), .A (n_207), .B (n_209));
HA_X1 i_636 (.CO (n_209), .S (n_208), .A (n_179), .B (n_181));
FA_X1 i_635 (.CO (n_207), .S (n_206), .A (n_177), .B (n_202), .CI (n_204));
FA_X1 i_634 (.CO (n_237), .S (n_236), .A (n_232), .B (n_205), .CI (n_234));
FA_X1 i_633 (.CO (n_205), .S (n_204), .A (n_196), .B (n_175), .CI (n_200));
HA_X1 i_632 (.CO (n_305), .S (n_304), .A (n_269), .B (n_302));
FA_X1 i_631 (.CO (n_269), .S (n_268), .A (n_235), .B (n_264), .CI (n_266));
FA_X1 i_630 (.CO (n_235), .S (n_234), .A (n_226), .B (n_230), .CI (n_203));
HA_X1 i_629 (.CO (n_379), .S (n_378), .A (n_339), .B (n_341));
HA_X1 i_628 (.CO (n_341), .S (n_340), .A (n_303), .B (n_338));
FA_X1 i_627 (.CO (n_303), .S (n_302), .A (n_267), .B (n_298), .CI (n_300));
FA_X1 i_626 (.CO (n_267), .S (n_266), .A (n_260), .B (n_262), .CI (n_233));
FA_X1 i_625 (.CO (n_233), .S (n_232), .A (n_224), .B (n_201), .CI (n_228));
FA_X1 i_624 (.CO (n_339), .S (n_338), .A (n_334), .B (n_301), .CI (n_336));
FA_X1 i_623 (.CO (n_301), .S (n_300), .A (n_294), .B (n_265), .CI (n_296));
FA_X1 i_622 (.CO (n_265), .S (n_264), .A (n_231), .B (n_258), .CI (n_256));
FA_X1 i_621 (.CO (n_231), .S (n_230), .A (n_222), .B (n_199), .CI (n_197));
HA_X1 i_620 (.CO (n_419), .S (n_418), .A (n_377), .B (n_416));
FA_X1 i_619 (.CO (n_377), .S (n_376), .A (n_337), .B (n_372), .CI (n_374));
FA_X1 i_618 (.CO (n_337), .S (n_336), .A (n_330), .B (n_299), .CI (n_332));
FA_X1 i_617 (.CO (n_299), .S (n_298), .A (n_261), .B (n_292), .CI (n_290));
FA_X1 i_616 (.CO (n_261), .S (n_260), .A (n_240), .B (n_225), .CI (n_254));
FA_X1 i_615 (.CO (n_225), .S (n_224), .A (n_183), .B (n_195), .CI (n_193));
FA_X1 i_614 (.CO (n_193), .S (n_192), .A (n_756), .B (n_162), .CI (n_160));
FA_X1 i_613 (.CO (n_195), .S (n_194), .A (n_158), .B (n_156), .CI (n_140));
FA_X1 i_612 (.CO (n_183), .S (n_182), .A (n_700), .B (n_703), .CI (n_705));
HA_X1 i_611 (.CO (n_938), .S (n_460), .A (n_417), .B (n_458));
FA_X1 i_610 (.CO (n_417), .S (n_416), .A (n_375), .B (n_412), .CI (n_414));
FA_X1 i_609 (.CO (n_375), .S (n_374), .A (n_333), .B (n_335), .CI (n_370));
FA_X1 i_608 (.CO (n_335), .S (n_334), .A (n_326), .B (n_324), .CI (n_297));
FA_X1 i_607 (.CO (n_297), .S (n_296), .A (n_257), .B (n_288), .CI (n_263));
FA_X1 i_606 (.CO (n_263), .S (n_262), .A (n_252), .B (n_229), .CI (n_227));
FA_X1 i_605 (.CO (n_227), .S (n_226), .A (n_220), .B (n_218), .CI (n_216));
FA_X1 i_604 (.CO (n_229), .S (n_228), .A (n_214), .B (n_212), .CI (n_210));
FA_X1 i_603 (.CO (n_257), .S (n_256), .A (n_221), .B (n_250), .CI (n_248));
FA_X1 i_602 (.CO (n_221), .S (n_220), .A (n_1547), .B (n_1568), .CI (n_191));
FA_X1 i_601 (.CO (n_191), .S (n_190), .A (n_1502), .B (n_1525), .CI (n_1548));
FA_X1 i_600 (.CO (n_333), .S (n_332), .A (n_293), .B (n_295), .CI (n_328));
FA_X1 i_599 (.CO (n_295), .S (n_294), .A (n_286), .B (n_284), .CI (n_259));
FA_X1 i_598 (.CO (n_259), .S (n_258), .A (n_246), .B (n_244), .CI (n_242));
FA_X1 i_597 (.CO (n_293), .S (n_292), .A (n_274), .B (n_272), .CI (n_255));
FA_X1 i_596 (.CO (n_255), .S (n_254), .A (n_213), .B (n_211), .CI (n_223));
FA_X1 i_595 (.CO (n_223), .S (n_222), .A (n_189), .B (n_187), .CI (n_185));
FA_X1 i_594 (.CO (n_185), .S (n_184), .A (n_1295), .B (n_1318), .CI (n_1341));
FA_X1 i_593 (.CO (n_187), .S (n_186), .A (n_1364), .B (n_1387), .CI (n_1410));
FA_X1 i_592 (.CO (n_189), .S (n_188), .A (n_1433), .B (n_1456), .CI (n_1479));
FA_X1 i_591 (.CO (n_211), .S (n_210), .A (n_1202), .B (n_1225), .CI (n_1248));
FA_X1 i_590 (.CO (n_213), .S (n_212), .A (n_1271), .B (n_1294), .CI (n_1317));
HA_X1 i_589 (.CO (n_921), .S (n_900), .A (n_503), .B (n_546));
FA_X1 i_588 (.CO (n_879), .S (n_546), .A (n_542), .B (n_501), .CI (n_544));
FA_X1 i_587 (.CO (n_878), .S (n_544), .A (n_499), .B (n_538), .CI (n_540));
FA_X1 i_586 (.CO (n_855), .S (n_540), .A (n_528), .B (n_493), .CI (n_536));
FA_X1 i_585 (.CO (n_854), .S (n_536), .A (n_487), .B (n_485), .CI (n_526));
FA_X1 i_584 (.CO (n_829), .S (n_526), .A (n_463), .B (n_481), .CI (n_479));
FA_X1 i_583 (.CO (n_828), .S (n_528), .A (n_520), .B (n_518), .CI (n_516));
FA_X1 i_582 (.CO (n_801), .S (n_516), .A (n_1378), .B (n_1401), .CI (n_1424));
FA_X1 i_581 (.CO (n_800), .S (n_518), .A (n_1447), .B (n_1470), .CI (n_1493));
FA_X1 i_580 (.CO (n_793), .S (n_520), .A (n_1516), .B (n_1539), .CI (n_477));
FA_X1 i_579 (.CO (n_792), .S (n_538), .A (n_491), .B (n_532), .CI (n_530));
FA_X1 i_578 (.CO (n_791), .S (n_530), .A (n_514), .B (n_512), .CI (n_510));
FA_X1 i_577 (.CO (n_790), .S (n_510), .A (n_1171), .B (n_1194), .CI (n_1217));
FA_X1 i_576 (.CO (n_789), .S (n_512), .A (n_1240), .B (n_1263), .CI (n_1286));
FA_X1 i_575 (.CO (n_788), .S (n_514), .A (n_1309), .B (n_1332), .CI (n_1355));
FA_X1 i_574 (.CO (n_787), .S (n_532), .A (n_508), .B (n_506), .CI (n_483));
FA_X1 i_573 (.CO (n_786), .S (n_506), .A (n_1033), .B (n_1056), .CI (n_1079));
FA_X1 i_572 (.CO (n_785), .S (n_508), .A (n_1102), .B (n_1125), .CI (n_1148));
FA_X1 i_571 (.CO (n_783), .S (n_542), .A (n_534), .B (n_495), .CI (n_497));
FA_X1 i_570 (.CO (n_780), .S (n_534), .A (n_524), .B (n_522), .CI (n_489));
FA_X1 i_569 (.CO (n_778), .S (n_522), .A (n_475), .B (n_473), .CI (n_471));
FA_X1 i_568 (.CO (n_776), .S (n_524), .A (n_469), .B (n_467), .CI (n_465));
HA_X1 i_567 (.CO (n_775), .S (n_773), .A (n_459), .B (n_502));
FA_X1 i_566 (.CO (n_503), .S (n_502), .A (n_498), .B (n_457), .CI (n_500));
FA_X1 i_565 (.CO (n_501), .S (n_500), .A (n_494), .B (n_455), .CI (n_496));
FA_X1 i_564 (.CO (n_497), .S (n_496), .A (n_486), .B (n_484), .CI (n_451));
FA_X1 i_563 (.CO (n_485), .S (n_484), .A (n_435), .B (n_476), .CI (n_474));
FA_X1 i_562 (.CO (n_475), .S (n_474), .A (n_1448), .B (n_1471), .CI (n_1494));
FA_X1 i_561 (.CO (n_477), .S (n_476), .A (n_1517), .B (n_1540), .CI (n_1561));
FA_X1 i_560 (.CO (n_487), .S (n_486), .A (n_472), .B (n_470), .CI (n_468));
FA_X1 i_559 (.CO (n_469), .S (n_468), .A (n_1241), .B (n_1264), .CI (n_1287));
FA_X1 i_558 (.CO (n_471), .S (n_470), .A (n_1310), .B (n_1333), .CI (n_1356));
FA_X1 i_557 (.CO (n_473), .S (n_472), .A (n_1379), .B (n_1402), .CI (n_1425));
FA_X1 i_556 (.CO (n_495), .S (n_494), .A (n_449), .B (n_447), .CI (n_488));
FA_X1 i_555 (.CO (n_489), .S (n_488), .A (n_466), .B (n_464), .CI (n_462));
FA_X1 i_554 (.CO (n_463), .S (n_462), .A (n_1034), .B (n_1057), .CI (n_1080));
FA_X1 i_553 (.CO (n_465), .S (n_464), .A (n_1103), .B (n_1126), .CI (n_1149));
FA_X1 i_552 (.CO (n_467), .S (n_466), .A (n_1172), .B (n_1195), .CI (n_1218));
FA_X1 i_551 (.CO (n_499), .S (n_498), .A (n_492), .B (n_490), .CI (n_453));
FA_X1 i_550 (.CO (n_491), .S (n_490), .A (n_480), .B (n_478), .CI (n_445));
FA_X1 i_549 (.CO (n_479), .S (n_478), .A (n_433), .B (n_431), .CI (n_429));
FA_X1 i_548 (.CO (n_481), .S (n_480), .A (n_427), .B (n_425), .CI (n_423));
FA_X1 i_547 (.CO (n_493), .S (n_492), .A (n_443), .B (n_441), .CI (n_482));
FA_X1 i_546 (.CO (n_483), .S (n_482), .A (n_421), .B (n_439), .CI (n_437));
FA_X1 i_545 (.CO (n_459), .S (n_458), .A (n_454), .B (n_415), .CI (n_456));
FA_X1 i_544 (.CO (n_457), .S (n_456), .A (n_450), .B (n_413), .CI (n_452));
FA_X1 i_543 (.CO (n_453), .S (n_452), .A (n_444), .B (n_442), .CI (n_446));
FA_X1 i_542 (.CO (n_447), .S (n_446), .A (n_420), .B (n_399), .CI (n_438));
FA_X1 i_541 (.CO (n_439), .S (n_438), .A (n_385), .B (n_383), .CI (n_381));
FA_X1 i_540 (.CO (n_421), .S (n_420), .A (n_1058), .B (n_1081), .CI (n_1104));
FA_X1 i_539 (.CO (n_443), .S (n_442), .A (n_432), .B (n_430), .CI (n_428));
FA_X1 i_538 (.CO (n_429), .S (n_428), .A (n_1334), .B (n_1357), .CI (n_1380));
FA_X1 i_537 (.CO (n_431), .S (n_430), .A (n_1403), .B (n_1426), .CI (n_1449));
FA_X1 i_536 (.CO (n_433), .S (n_432), .A (n_1472), .B (n_1495), .CI (n_1518));
FA_X1 i_535 (.CO (n_445), .S (n_444), .A (n_426), .B (n_424), .CI (n_422));
FA_X1 i_534 (.CO (n_423), .S (n_422), .A (n_1127), .B (n_1150), .CI (n_1173));
FA_X1 i_533 (.CO (n_425), .S (n_424), .A (n_1196), .B (n_1219), .CI (n_1242));
FA_X1 i_532 (.CO (n_427), .S (n_426), .A (n_1265), .B (n_1288), .CI (n_1311));
FA_X1 i_531 (.CO (n_413), .S (n_412), .A (n_369), .B (n_408), .CI (n_406));
FA_X1 i_530 (.CO (n_451), .S (n_450), .A (n_440), .B (n_407), .CI (n_405));
FA_X1 i_529 (.CO (n_407), .S (n_406), .A (n_396), .B (n_394), .CI (n_365));
FA_X1 i_528 (.CO (n_441), .S (n_440), .A (n_397), .B (n_395), .CI (n_434));
FA_X1 i_527 (.CO (n_435), .S (n_434), .A (n_1541), .B (n_1562), .CI (n_393));
FA_X1 i_526 (.CO (n_395), .S (n_394), .A (n_1563), .B (n_355), .CI (n_353));
FA_X1 i_525 (.CO (n_397), .S (n_396), .A (n_351), .B (n_349), .CI (n_347));
FA_X1 i_524 (.CO (n_415), .S (n_414), .A (n_371), .B (n_373), .CI (n_410));
FA_X1 i_523 (.CO (n_373), .S (n_372), .A (n_362), .B (n_368), .CI (n_366));
FA_X1 i_522 (.CO (n_369), .S (n_368), .A (n_327), .B (n_325), .CI (n_360));
FA_X1 i_521 (.CO (n_325), .S (n_324), .A (n_285), .B (n_318), .CI (n_316));
FA_X1 i_520 (.CO (n_285), .S (n_284), .A (n_1566), .B (n_251), .CI (n_249));
FA_X1 i_519 (.CO (n_249), .S (n_248), .A (n_1454), .B (n_1477), .CI (n_1500));
FA_X1 i_518 (.CO (n_251), .S (n_250), .A (n_1523), .B (n_1546), .CI (n_1567));
FA_X1 i_517 (.CO (n_327), .S (n_326), .A (n_314), .B (n_312), .CI (n_310));
FA_X1 i_516 (.CO (n_371), .S (n_370), .A (n_331), .B (n_329), .CI (n_364));
FA_X1 i_515 (.CO (n_365), .S (n_364), .A (n_346), .B (n_344), .CI (n_342));
FA_X1 i_514 (.CO (n_347), .S (n_346), .A (n_1244), .B (n_1267), .CI (n_1290));
FA_X1 i_513 (.CO (n_329), .S (n_328), .A (n_308), .B (n_306), .CI (n_322));
FA_X1 i_512 (.CO (n_331), .S (n_330), .A (n_320), .B (n_291), .CI (n_289));
FA_X1 i_511 (.CO (n_289), .S (n_288), .A (n_241), .B (n_253), .CI (n_282));
FA_X1 i_510 (.CO (n_253), .S (n_252), .A (n_219), .B (n_217), .CI (n_215));
FA_X1 i_509 (.CO (n_215), .S (n_214), .A (n_1340), .B (n_1363), .CI (n_1386));
FA_X1 i_508 (.CO (n_217), .S (n_216), .A (n_1409), .B (n_1432), .CI (n_1455));
FA_X1 i_507 (.CO (n_219), .S (n_218), .A (n_1478), .B (n_1501), .CI (n_1524));
FA_X1 i_506 (.CO (n_241), .S (n_240), .A (n_1178), .B (n_1201), .CI (n_1224));
FA_X1 i_505 (.CO (n_291), .S (n_290), .A (n_280), .B (n_278), .CI (n_276));
FA_X1 i_504 (.CO (n_455), .S (n_454), .A (n_409), .B (n_448), .CI (n_411));
FA_X1 i_503 (.CO (n_411), .S (n_410), .A (n_404), .B (n_402), .CI (n_400));
FA_X1 i_502 (.CO (n_405), .S (n_404), .A (n_382), .B (n_380), .CI (n_398));
FA_X1 i_501 (.CO (n_399), .S (n_398), .A (n_345), .B (n_343), .CI (n_359));
FA_X1 i_500 (.CO (n_343), .S (n_342), .A (n_1106), .B (n_1129), .CI (n_1152));
FA_X1 i_499 (.CO (n_345), .S (n_344), .A (n_1175), .B (n_1198), .CI (n_1221));
FA_X1 i_498 (.CO (n_381), .S (n_380), .A (n_1082), .B (n_1105), .CI (n_1128));
FA_X1 i_497 (.CO (n_383), .S (n_382), .A (n_1151), .B (n_1174), .CI (n_1197));
FA_X1 i_496 (.CO (n_449), .S (n_448), .A (n_436), .B (n_403), .CI (n_401));
FA_X1 i_495 (.CO (n_401), .S (n_400), .A (n_357), .B (n_392), .CI (n_390));
FA_X1 i_494 (.CO (n_393), .S (n_392), .A (n_1496), .B (n_1519), .CI (n_1542));
FA_X1 i_493 (.CO (n_403), .S (n_402), .A (n_388), .B (n_386), .CI (n_384));
FA_X1 i_492 (.CO (n_385), .S (n_384), .A (n_1220), .B (n_1243), .CI (n_1266));
FA_X1 i_491 (.CO (n_437), .S (n_436), .A (n_391), .B (n_389), .CI (n_387));
FA_X1 i_490 (.CO (n_387), .S (n_386), .A (n_1289), .B (n_1312), .CI (n_1335));
FA_X1 i_489 (.CO (n_389), .S (n_388), .A (n_1358), .B (n_1381), .CI (n_1404));
FA_X1 i_488 (.CO (n_391), .S (n_390), .A (n_1427), .B (n_1450), .CI (n_1473));
FA_X1 i_487 (.CO (n_409), .S (n_408), .A (n_363), .B (n_361), .CI (n_367));
FA_X1 i_486 (.CO (n_367), .S (n_366), .A (n_323), .B (n_358), .CI (n_356));
FA_X1 i_485 (.CO (n_357), .S (n_356), .A (n_317), .B (n_315), .CI (n_313));
FA_X1 i_484 (.CO (n_313), .S (n_312), .A (n_1337), .B (n_1360), .CI (n_1383));
FA_X1 i_483 (.CO (n_315), .S (n_314), .A (n_1406), .B (n_1429), .CI (n_1452));
FA_X1 i_482 (.CO (n_317), .S (n_316), .A (n_1475), .B (n_1498), .CI (n_1521));
FA_X1 i_481 (.CO (n_359), .S (n_358), .A (n_311), .B (n_309), .CI (n_307));
FA_X1 i_480 (.CO (n_307), .S (n_306), .A (n_1130), .B (n_1153), .CI (n_1176));
FA_X1 i_479 (.CO (n_309), .S (n_308), .A (n_1199), .B (n_1222), .CI (n_1245));
FA_X1 i_478 (.CO (n_311), .S (n_310), .A (n_1268), .B (n_1291), .CI (n_1314));
FA_X1 i_477 (.CO (n_323), .S (n_322), .A (n_275), .B (n_273), .CI (n_287));
FA_X1 i_476 (.CO (n_287), .S (n_286), .A (n_247), .B (n_245), .CI (n_243));
FA_X1 i_475 (.CO (n_243), .S (n_242), .A (n_1247), .B (n_1270), .CI (n_1293));
FA_X1 i_474 (.CO (n_245), .S (n_244), .A (n_1316), .B (n_1339), .CI (n_1362));
FA_X1 i_473 (.CO (n_247), .S (n_246), .A (n_1385), .B (n_1408), .CI (n_1431));
FA_X1 i_472 (.CO (n_273), .S (n_272), .A (n_1154), .B (n_1177), .CI (n_1200));
FA_X1 i_471 (.CO (n_275), .S (n_274), .A (n_1223), .B (n_1246), .CI (n_1269));
FA_X1 i_470 (.CO (n_361), .S (n_360), .A (n_321), .B (n_319), .CI (n_354));
FA_X1 i_469 (.CO (n_355), .S (n_354), .A (n_1520), .B (n_1543), .CI (n_1564));
FA_X1 i_468 (.CO (n_319), .S (n_318), .A (n_1544), .B (n_1565), .CI (n_283));
FA_X1 i_467 (.CO (n_283), .S (n_282), .A (n_1499), .B (n_1522), .CI (n_1545));
FA_X1 i_466 (.CO (n_321), .S (n_320), .A (n_281), .B (n_279), .CI (n_277));
FA_X1 i_465 (.CO (n_277), .S (n_276), .A (n_1292), .B (n_1315), .CI (n_1338));
FA_X1 i_464 (.CO (n_279), .S (n_278), .A (n_1361), .B (n_1384), .CI (n_1407));
FA_X1 i_463 (.CO (n_281), .S (n_280), .A (n_1430), .B (n_1453), .CI (n_1476));
FA_X1 i_462 (.CO (n_363), .S (n_362), .A (n_352), .B (n_350), .CI (n_348));
FA_X1 i_461 (.CO (n_349), .S (n_348), .A (n_1313), .B (n_1336), .CI (n_1359));
FA_X1 i_460 (.CO (n_351), .S (n_350), .A (n_1382), .B (n_1405), .CI (n_1428));
FA_X1 i_459 (.CO (n_353), .S (n_352), .A (n_1451), .B (n_1474), .CI (n_1497));
INV_X1 i_458 (.ZN (n_1773), .A (n_0));
INV_X1 i_457 (.ZN (n_1767), .A (n_1813));
NAND2_X1 i_456 (.ZN (n_1765), .A1 (hfn_ipo_n6), .A2 (n_1767));
NOR2_X2 i_455 (.ZN (n_1763), .A1 (n_938), .A2 (n_773));
NOR3_X1 i_454 (.ZN (n_771), .A1 (n_1763), .A2 (n_1586), .A3 (n_1583));
NOR2_X1 i_453 (.ZN (n_1757), .A1 (n_1711), .A2 (n_1706));
INV_X1 i_452 (.ZN (n_1756), .A (n_1757));
OAI21_X1 i_451 (.ZN (n_770), .A (n_1756), .B1 (n_1707), .B2 (n_1704));
NOR2_X1 i_450 (.ZN (n_769), .A1 (n_1713), .A2 (n_1708));
NOR2_X2 i_449 (.ZN (n_1750), .A1 (n_591), .A2 (n_630));
INV_X1 i_448 (.ZN (n_1749), .A (n_1750));
NOR2_X1 i_447 (.ZN (n_1748), .A1 (n_168), .A2 (n_1712));
INV_X1 i_446 (.ZN (n_1747), .A (n_1748));
NAND3_X1 i_445 (.ZN (n_768), .A1 (n_1776), .A2 (n_1747), .A3 (n_1749));
NOR2_X1 i_444 (.ZN (n_764), .A1 (n_921), .A2 (n_590));
AND2_X1 i_443 (.ZN (n_1724), .A1 (n_2), .A2 (n_4));
NOR2_X1 i_442 (.ZN (n_1723), .A1 (n_1656), .A2 (n_1628));
AOI22_X1 i_441 (.ZN (n_1722), .A1 (A_imm[2]), .A2 (n_0), .B1 (A_imm[0]), .B2 (n_1723));
AOI211_X1 i_440 (.ZN (n_1721), .A (n_1655), .B (n_1722), .C1 (n_1629), .C2 (n_1773));
OAI222_X1 i_439 (.ZN (n_763), .A1 (n_954), .A2 (n_955), .B1 (n_2), .B2 (n_4), .C1 (n_1724), .C2 (n_1721));
INV_X1 i_438 (.ZN (n_1702), .A (n_1569));
OAI21_X1 i_437 (.ZN (n_762), .A (n_771), .B1 (n_1513), .B2 (n_1702));
NAND2_X1 i_436 (.ZN (n_761), .A1 (n_1709), .A2 (n_1710));
NAND2_X1 i_435 (.ZN (n_760), .A1 (n_921), .A2 (n_590));
NAND2_X1 i_434 (.ZN (n_758), .A1 (n_591), .A2 (n_630));
INV_X1 i_433 (.ZN (n_1689), .A (n_758));
INV_X1 i_432 (.ZN (n_1671), .A (n_1760));
AOI21_X1 i_431 (.ZN (n_1638), .A (n_1815), .B1 (n_1795), .B2 (n_1812));
AOI21_X1 i_430 (.ZN (n_1637), .A (n_1638), .B1 (n_1819), .B2 (n_1821));
NAND2_X1 i_429 (.ZN (n_1636), .A1 (n_1765), .A2 (n_1637));
OAI21_X1 i_428 (.ZN (Res_imm[47]), .A (n_1636), .B1 (hfn_ipo_n6), .B2 (n_1767));
OAI21_X1 i_427 (.ZN (n_1635), .A (n_1765), .B1 (hfn_ipo_n6), .B2 (n_1767));
XNOR2_X1 i_426 (.ZN (Res_imm[46]), .A (n_1637), .B (n_1635));
NOR2_X1 i_425 (.ZN (n_1627), .A1 (n_1800), .A2 (n_1811));
OAI22_X1 i_424 (.ZN (n_1626), .A1 (n_1784), .A2 (n_1796), .B1 (n_1806), .B2 (n_1804));
XNOR2_X1 i_423 (.ZN (Res_imm[43]), .A (n_1627), .B (n_1626));
XOR2_X1 i_422 (.Z (Res_imm[42]), .A (n_1804), .B (n_1810));
OAI21_X1 i_421 (.ZN (n_1624), .A (n_1719), .B1 (n_1694), .B2 (n_1692));
AOI21_X1 i_420 (.ZN (n_1620), .A (n_1769), .B1 (n_1693), .B2 (n_1686));
NOR2_X1 i_419 (.ZN (n_1618), .A1 (n_1791), .A2 (n_1770));
XOR2_X1 i_418 (.Z (Res_imm[39]), .A (n_1716), .B (n_1618));
XOR2_X1 i_417 (.Z (Res_imm[38]), .A (n_1718), .B (n_1620));
XOR2_X1 i_416 (.Z (Res_imm[37]), .A (n_1720), .B (n_1624));
NOR2_X1 i_415 (.ZN (n_1617), .A1 (n_1761), .A2 (n_1762));
OAI21_X1 i_414 (.ZN (n_1616), .A (n_1755), .B1 (n_1703), .B2 (n_1698));
AOI21_X2 i_413 (.ZN (n_1615), .A (n_1753), .B1 (n_1729), .B2 (n_1755));
INV_X1 i_412 (.ZN (n_1614), .A (n_1615));
AOI21_X1 i_411 (.ZN (n_1613), .A (n_1758), .B1 (n_1754), .B2 (n_1614));
AOI21_X1 i_410 (.ZN (n_1612), .A (n_1758), .B1 (n_1699), .B2 (n_1696));
OAI22_X1 i_409 (.ZN (n_1611), .A1 (n_1697), .A2 (n_1695), .B1 (n_1671), .B2 (n_1613));
XNOR2_X1 i_408 (.ZN (Res_imm[36]), .A (n_1617), .B (n_1611));
NOR2_X1 i_407 (.ZN (n_1610), .A1 (n_1759), .A2 (n_1671));
XOR2_X1 i_406 (.Z (Res_imm[35]), .A (n_1613), .B (n_1610));
XOR2_X2 i_405 (.Z (Res_imm[34]), .A (n_1615), .B (n_1612));
XOR2_X1 i_404 (.Z (Res_imm[33]), .A (n_1729), .B (n_1616));
OAI22_X1 i_403 (.ZN (n_1609), .A1 (n_1705), .A2 (n_1701), .B1 (n_1777), .B2 (n_1778));
INV_X1 i_402 (.ZN (n_1607), .A (n_977));
OAI21_X1 i_401 (.ZN (n_1606), .A (n_1740), .B1 (n_1738), .B2 (n_1607));
INV_X2 i_400 (.ZN (n_1605), .A (n_1606));
OAI21_X1 i_399 (.ZN (n_1604), .A (n_1745), .B1 (n_1742), .B2 (n_1605));
OAI21_X1 i_398 (.ZN (n_1603), .A (n_761), .B1 (n_1709), .B2 (n_1710));
OAI22_X1 i_397 (.ZN (n_1602), .A1 (n_1709), .A2 (n_1710), .B1 (n_1775), .B2 (n_1604));
INV_X1 i_396 (.ZN (n_1601), .A (n_1602));
OR2_X1 i_395 (.ZN (n_1600), .A1 (n_1757), .A2 (n_1744));
NOR2_X1 i_394 (.ZN (n_1599), .A1 (n_1601), .A2 (n_1600));
OAI21_X1 i_393 (.ZN (n_1598), .A (n_1752), .B1 (n_770), .B2 (n_1599));
XNOR2_X1 i_392 (.ZN (Res_imm[32]), .A (n_1609), .B (n_1598));
OAI21_X1 i_391 (.ZN (n_1597), .A (n_1752), .B1 (n_1707), .B2 (n_1704));
OAI21_X1 i_390 (.ZN (n_1596), .A (n_1756), .B1 (n_1744), .B2 (n_1601));
XOR2_X1 i_389 (.Z (Res_imm[31]), .A (n_1597), .B (n_1596));
AOI21_X1 i_388 (.ZN (n_1595), .A (n_1599), .B1 (n_1601), .B2 (n_1600));
INV_X1 i_387 (.ZN (Res_imm[30]), .A (n_1595));
XNOR2_X1 i_386 (.ZN (Res_imm[29]), .A (n_1604), .B (n_1603));
AOI21_X1 i_385 (.ZN (n_1594), .A (n_769), .B1 (n_1713), .B2 (n_1708));
OAI21_X1 i_384 (.ZN (n_1593), .A (n_760), .B1 (n_921), .B2 (n_590));
AOI21_X2 i_383 (.ZN (n_1592), .A (n_764), .B1 (n_760), .B2 (n_1605));
OAI21_X1 i_382 (.ZN (n_1591), .A (n_1749), .B1 (n_1689), .B2 (n_1592));
INV_X1 i_381 (.ZN (n_1590), .A (n_1591));
NOR2_X1 i_380 (.ZN (n_1589), .A1 (n_1750), .A2 (n_1689));
OAI21_X1 i_379 (.ZN (n_1588), .A (n_1747), .B1 (n_1751), .B2 (n_1590));
XNOR2_X1 i_378 (.ZN (Res_imm[28]), .A (n_1594), .B (n_1588));
NOR2_X1 i_377 (.ZN (n_1587), .A1 (n_1748), .A2 (n_1751));
XOR2_X2 i_376 (.Z (Res_imm[27]), .A (n_1590), .B (n_1587));
XOR2_X2 i_375 (.Z (Res_imm[26]), .A (n_1592), .B (n_1589));
XOR2_X1 i_374 (.Z (Res_imm[25]), .A (n_1605), .B (n_1593));
NOR2_X1 i_373 (.ZN (n_1582), .A1 (n_1763), .A2 (n_1584));
XOR2_X2 i_372 (.Z (Res_imm[23]), .A (n_973), .B (n_1582));
NOR2_X1 i_371 (.ZN (n_1581), .A1 (n_1655), .A2 (n_1630));
NOR2_X1 i_370 (.ZN (n_1580), .A1 (n_1655), .A2 (n_1631));
NOR2_X1 i_369 (.ZN (n_1579), .A1 (n_1655), .A2 (n_1632));
NOR2_X1 i_368 (.ZN (n_1578), .A1 (n_1655), .A2 (n_1633));
NOR2_X1 i_367 (.ZN (n_1577), .A1 (n_1655), .A2 (n_1634));
NOR2_X1 i_366 (.ZN (n_1576), .A1 (n_1655), .A2 (n_1639));
NOR2_X1 i_365 (.ZN (n_1575), .A1 (n_1655), .A2 (n_1640));
NOR2_X1 i_364 (.ZN (n_1574), .A1 (n_1655), .A2 (n_1641));
NOR2_X1 i_1067 (.ZN (n_1573), .A1 (n_1655), .A2 (n_1642));
NOR2_X1 i_1066 (.ZN (n_1572), .A1 (n_1655), .A2 (n_1643));
NOR2_X1 i_363 (.ZN (n_1571), .A1 (n_1655), .A2 (n_1644));
NOR2_X1 i_1064 (.ZN (n_1570), .A1 (n_1655), .A2 (n_1645));
NOR2_X1 i_362 (.ZN (n_756), .A1 (n_1655), .A2 (n_1646));
NOR2_X1 i_361 (.ZN (n_1560), .A1 (n_1656), .A2 (n_1629));
NOR2_X1 i_360 (.ZN (n_1559), .A1 (n_1656), .A2 (n_1630));
NOR2_X1 i_359 (.ZN (n_1558), .A1 (n_1656), .A2 (n_1631));
NOR2_X1 i_358 (.ZN (n_1557), .A1 (n_1656), .A2 (n_1632));
NOR2_X1 i_357 (.ZN (n_1556), .A1 (n_1656), .A2 (n_1633));
NOR2_X1 i_356 (.ZN (n_1555), .A1 (n_1656), .A2 (n_1634));
NOR2_X1 i_355 (.ZN (n_1554), .A1 (n_1656), .A2 (n_1639));
NOR2_X1 i_354 (.ZN (n_1553), .A1 (n_1656), .A2 (n_1640));
NOR2_X1 i_1046 (.ZN (n_1552), .A1 (n_1656), .A2 (n_1641));
NOR2_X1 i_353 (.ZN (n_1551), .A1 (n_1656), .A2 (n_1642));
NOR2_X1 i_352 (.ZN (n_1550), .A1 (n_1656), .A2 (n_1643));
NOR2_X1 i_1043 (.ZN (n_1549), .A1 (n_1656), .A2 (n_1644));
NOR2_X1 i_351 (.ZN (n_1538), .A1 (n_1657), .A2 (n_1625));
NOR2_X1 i_350 (.ZN (n_1537), .A1 (n_1657), .A2 (n_1628));
NOR2_X1 i_349 (.ZN (n_739), .A1 (n_1657), .A2 (n_1629));
NOR2_X1 i_348 (.ZN (n_1535), .A1 (n_1657), .A2 (n_1630));
NOR2_X1 i_347 (.ZN (n_1534), .A1 (n_1657), .A2 (n_1631));
NOR2_X1 i_346 (.ZN (n_1533), .A1 (n_1657), .A2 (n_1632));
NOR2_X1 i_345 (.ZN (n_1532), .A1 (n_1657), .A2 (n_1633));
NOR2_X1 i_344 (.ZN (n_1531), .A1 (n_1657), .A2 (n_1634));
NOR2_X1 i_343 (.ZN (n_1530), .A1 (n_1657), .A2 (n_1639));
NOR2_X1 i_1023 (.ZN (n_1529), .A1 (n_1657), .A2 (n_1640));
NOR2_X1 i_342 (.ZN (n_1528), .A1 (n_1657), .A2 (n_1641));
NOR2_X1 i_1021 (.ZN (n_1527), .A1 (n_1657), .A2 (n_1642));
NOR2_X1 i_1020 (.ZN (n_1526), .A1 (n_1657), .A2 (n_1643));
NOR2_X1 i_341 (.ZN (n_1515), .A1 (n_1657), .A2 (n_1654));
NOR2_X1 i_340 (.ZN (n_1514), .A1 (n_1658), .A2 (n_1625));
NOR2_X1 i_339 (.ZN (n_738), .A1 (n_1658), .A2 (n_1628));
NOR2_X1 i_338 (.ZN (n_1512), .A1 (n_1658), .A2 (n_1629));
NOR2_X1 i_337 (.ZN (n_1511), .A1 (n_1658), .A2 (n_1630));
NOR2_X1 i_336 (.ZN (n_1510), .A1 (n_1658), .A2 (n_1631));
NOR2_X1 i_335 (.ZN (n_1509), .A1 (n_1658), .A2 (n_1632));
NOR2_X1 i_334 (.ZN (n_1508), .A1 (n_1658), .A2 (n_1633));
NOR2_X1 i_333 (.ZN (n_1507), .A1 (n_1658), .A2 (n_1634));
NOR2_X1 i_1000 (.ZN (n_1506), .A1 (n_1658), .A2 (n_1639));
NOR2_X1 i_332 (.ZN (n_1505), .A1 (n_1658), .A2 (n_1640));
NOR2_X1 i_998 (.ZN (n_1504), .A1 (n_1658), .A2 (n_1641));
NOR2_X1 i_997 (.ZN (n_1503), .A1 (n_1658), .A2 (n_1642));
NOR2_X1 i_331 (.ZN (n_1492), .A1 (n_1658), .A2 (n_1653));
NOR2_X1 i_330 (.ZN (n_1491), .A1 (n_1658), .A2 (n_1654));
NOR2_X1 i_329 (.ZN (n_737), .A1 (n_1659), .A2 (n_1625));
NOR2_X1 i_328 (.ZN (n_1489), .A1 (n_1659), .A2 (n_1628));
NOR2_X1 i_327 (.ZN (n_1488), .A1 (n_1659), .A2 (n_1629));
NOR2_X1 i_326 (.ZN (n_1487), .A1 (n_1659), .A2 (n_1630));
NOR2_X1 i_325 (.ZN (n_1486), .A1 (n_1659), .A2 (n_1631));
NOR2_X1 i_324 (.ZN (n_1485), .A1 (n_1659), .A2 (n_1632));
NOR2_X1 i_323 (.ZN (n_1484), .A1 (n_1659), .A2 (n_1633));
NOR2_X1 i_977 (.ZN (n_1483), .A1 (n_1659), .A2 (n_1634));
NOR2_X1 i_976 (.ZN (n_1482), .A1 (n_1659), .A2 (n_1639));
NOR2_X1 i_975 (.ZN (n_1481), .A1 (n_1659), .A2 (n_1640));
NOR2_X1 i_974 (.ZN (n_1480), .A1 (n_1659), .A2 (n_1641));
NOR2_X1 i_322 (.ZN (n_1469), .A1 (n_1659), .A2 (n_1652));
NOR2_X1 i_321 (.ZN (n_1468), .A1 (n_1659), .A2 (n_1653));
NOR2_X1 i_320 (.ZN (n_1467), .A1 (n_1659), .A2 (n_1654));
NOR2_X1 i_319 (.ZN (n_1466), .A1 (n_1660), .A2 (n_1625));
NOR2_X1 i_318 (.ZN (n_1465), .A1 (n_1660), .A2 (n_1628));
NOR2_X1 i_317 (.ZN (n_1464), .A1 (n_1660), .A2 (n_1629));
NOR2_X1 i_316 (.ZN (n_1463), .A1 (n_1660), .A2 (n_1630));
NOR2_X1 i_315 (.ZN (n_1462), .A1 (n_1660), .A2 (n_1631));
NOR2_X1 i_314 (.ZN (n_1461), .A1 (n_1660), .A2 (n_1632));
NOR2_X1 i_954 (.ZN (n_1460), .A1 (n_1660), .A2 (n_1633));
NOR2_X1 i_953 (.ZN (n_1459), .A1 (n_1660), .A2 (n_1634));
NOR2_X1 i_952 (.ZN (n_1458), .A1 (n_1660), .A2 (n_1639));
NOR2_X1 i_951 (.ZN (n_1457), .A1 (n_1660), .A2 (n_1640));
NOR2_X1 i_313 (.ZN (n_1446), .A1 (n_1660), .A2 (n_1651));
NOR2_X1 i_312 (.ZN (n_1445), .A1 (n_1660), .A2 (n_1652));
NOR2_X1 i_311 (.ZN (n_1444), .A1 (n_1660), .A2 (n_1653));
NOR2_X1 i_310 (.ZN (n_1443), .A1 (n_1660), .A2 (n_1654));
NOR2_X1 i_309 (.ZN (n_1442), .A1 (n_1661), .A2 (n_1625));
NOR2_X1 i_308 (.ZN (n_1441), .A1 (n_1661), .A2 (n_1628));
NOR2_X1 i_307 (.ZN (n_1440), .A1 (n_1661), .A2 (n_1629));
NOR2_X1 i_306 (.ZN (n_1439), .A1 (n_1661), .A2 (n_1630));
NOR2_X1 i_305 (.ZN (n_1438), .A1 (n_1661), .A2 (n_1631));
NOR2_X1 i_931 (.ZN (n_1437), .A1 (n_1661), .A2 (n_1632));
NOR2_X1 i_930 (.ZN (n_1436), .A1 (n_1661), .A2 (n_1633));
NOR2_X1 i_929 (.ZN (n_1435), .A1 (n_1661), .A2 (n_1634));
NOR2_X1 i_928 (.ZN (n_1434), .A1 (n_1661), .A2 (n_1639));
NOR2_X1 i_304 (.ZN (n_1423), .A1 (n_1661), .A2 (n_1650));
NOR2_X1 i_303 (.ZN (n_1422), .A1 (n_1661), .A2 (n_1651));
NOR2_X1 i_302 (.ZN (n_1421), .A1 (n_1661), .A2 (n_1652));
NOR2_X1 i_301 (.ZN (n_1420), .A1 (n_1661), .A2 (n_1653));
NOR2_X1 i_300 (.ZN (n_1419), .A1 (n_1661), .A2 (n_1654));
NOR2_X1 i_299 (.ZN (n_1418), .A1 (n_1662), .A2 (n_1625));
NOR2_X1 i_298 (.ZN (n_1417), .A1 (n_1662), .A2 (n_1628));
NOR2_X1 i_297 (.ZN (n_1416), .A1 (n_1662), .A2 (n_1629));
NOR2_X1 i_296 (.ZN (n_1415), .A1 (n_1662), .A2 (n_1630));
NOR2_X1 i_908 (.ZN (n_1414), .A1 (n_1662), .A2 (n_1631));
NOR2_X1 i_907 (.ZN (n_1413), .A1 (n_1662), .A2 (n_1632));
NOR2_X1 i_906 (.ZN (n_1412), .A1 (n_1662), .A2 (n_1633));
NOR2_X1 i_905 (.ZN (n_1411), .A1 (n_1662), .A2 (n_1634));
NOR2_X1 i_295 (.ZN (n_1400), .A1 (n_1662), .A2 (n_1649));
NOR2_X1 i_294 (.ZN (n_1399), .A1 (n_1662), .A2 (n_1650));
NOR2_X1 i_293 (.ZN (n_1398), .A1 (n_1662), .A2 (n_1651));
NOR2_X1 i_292 (.ZN (n_1397), .A1 (n_1662), .A2 (n_1652));
NOR2_X1 i_291 (.ZN (n_1396), .A1 (n_1662), .A2 (n_1653));
NOR2_X1 i_290 (.ZN (n_1395), .A1 (n_1662), .A2 (n_1654));
NOR2_X1 i_289 (.ZN (n_1394), .A1 (n_1663), .A2 (n_1625));
NOR2_X1 i_288 (.ZN (n_1393), .A1 (n_1663), .A2 (n_1628));
NOR2_X1 i_287 (.ZN (n_1392), .A1 (n_1663), .A2 (n_1629));
NOR2_X1 i_885 (.ZN (n_1391), .A1 (n_1663), .A2 (n_1630));
NOR2_X1 i_884 (.ZN (n_1390), .A1 (n_1663), .A2 (n_1631));
NOR2_X1 i_883 (.ZN (n_1389), .A1 (n_1663), .A2 (n_1632));
NOR2_X1 i_882 (.ZN (n_1388), .A1 (n_1663), .A2 (n_1633));
NOR2_X1 i_286 (.ZN (n_1377), .A1 (n_1663), .A2 (n_1648));
NOR2_X1 i_285 (.ZN (n_1376), .A1 (n_1663), .A2 (n_1649));
NOR2_X1 i_284 (.ZN (n_1375), .A1 (n_1663), .A2 (n_1650));
NOR2_X1 i_283 (.ZN (n_1374), .A1 (n_1663), .A2 (n_1651));
NOR2_X1 i_282 (.ZN (n_1373), .A1 (n_1663), .A2 (n_1652));
NOR2_X1 i_281 (.ZN (n_1372), .A1 (n_1663), .A2 (n_1653));
NOR2_X1 i_280 (.ZN (n_1371), .A1 (n_1663), .A2 (n_1654));
NOR2_X1 i_279 (.ZN (n_1370), .A1 (n_1664), .A2 (n_1625));
NOR2_X1 i_278 (.ZN (n_1369), .A1 (n_1664), .A2 (n_1628));
NOR2_X1 i_862 (.ZN (n_1368), .A1 (n_1664), .A2 (n_1629));
NOR2_X1 i_861 (.ZN (n_1367), .A1 (n_1664), .A2 (n_1630));
NOR2_X1 i_860 (.ZN (n_1366), .A1 (n_1664), .A2 (n_1631));
NOR2_X1 i_859 (.ZN (n_1365), .A1 (n_1664), .A2 (n_1632));
NOR2_X1 i_277 (.ZN (n_1354), .A1 (n_1664), .A2 (n_1647));
NOR2_X1 i_276 (.ZN (n_1353), .A1 (n_1664), .A2 (n_1648));
NOR2_X1 i_275 (.ZN (n_1352), .A1 (n_1664), .A2 (n_1649));
NOR2_X1 i_274 (.ZN (n_1351), .A1 (n_1664), .A2 (n_1650));
NOR2_X1 i_273 (.ZN (n_1350), .A1 (n_1664), .A2 (n_1651));
NOR2_X1 i_272 (.ZN (n_1349), .A1 (n_1664), .A2 (n_1652));
NOR2_X1 i_271 (.ZN (n_736), .A1 (n_1664), .A2 (n_1653));
NOR2_X1 i_270 (.ZN (n_1346), .A1 (n_1665), .A2 (n_1625));
NOR2_X1 i_839 (.ZN (n_1345), .A1 (n_1665), .A2 (n_1628));
NOR2_X1 i_838 (.ZN (n_1344), .A1 (n_1665), .A2 (n_1629));
NOR2_X1 i_837 (.ZN (n_1343), .A1 (n_1665), .A2 (n_1630));
NOR2_X1 i_836 (.ZN (n_1342), .A1 (n_1665), .A2 (n_1631));
NOR2_X1 i_269 (.ZN (n_1331), .A1 (n_1665), .A2 (n_1646));
NOR2_X1 i_268 (.ZN (n_1330), .A1 (n_1665), .A2 (n_1647));
NOR2_X1 i_267 (.ZN (n_1329), .A1 (n_1665), .A2 (n_1648));
NOR2_X1 i_266 (.ZN (n_1328), .A1 (n_1665), .A2 (n_1649));
NOR2_X1 i_265 (.ZN (n_1327), .A1 (n_1665), .A2 (n_1650));
NOR2_X1 i_264 (.ZN (n_1326), .A1 (n_1665), .A2 (n_1651));
NOR2_X1 i_263 (.ZN (n_734), .A1 (n_1665), .A2 (n_1652));
NOR2_X1 i_816 (.ZN (n_1322), .A1 (n_1666), .A2 (n_1625));
NOR2_X1 i_815 (.ZN (n_1321), .A1 (n_1666), .A2 (n_1628));
NOR2_X1 i_262 (.ZN (n_1320), .A1 (n_1666), .A2 (n_1629));
NOR2_X1 i_813 (.ZN (n_1319), .A1 (n_1666), .A2 (n_1630));
NOR2_X1 i_261 (.ZN (n_1308), .A1 (n_1666), .A2 (n_1645));
NOR2_X1 i_260 (.ZN (n_1307), .A1 (n_1666), .A2 (n_1646));
NOR2_X1 i_259 (.ZN (n_1306), .A1 (n_1666), .A2 (n_1647));
NOR2_X1 i_258 (.ZN (n_1305), .A1 (n_1666), .A2 (n_1648));
NOR2_X1 i_257 (.ZN (n_1304), .A1 (n_1666), .A2 (n_1649));
NOR2_X1 i_256 (.ZN (n_1303), .A1 (n_1666), .A2 (n_1650));
NOR2_X1 i_255 (.ZN (n_731), .A1 (n_1666), .A2 (n_1651));
NOR2_X1 i_792 (.ZN (n_1298), .A1 (n_1667), .A2 (n_1625));
NOR2_X1 i_254 (.ZN (n_1297), .A1 (n_1667), .A2 (n_1628));
NOR2_X1 i_790 (.ZN (n_1296), .A1 (n_1667), .A2 (n_1629));
NOR2_X1 i_253 (.ZN (n_1285), .A1 (n_1667), .A2 (n_1644));
NOR2_X1 i_252 (.ZN (n_1284), .A1 (n_1667), .A2 (n_1645));
NOR2_X1 i_251 (.ZN (n_1283), .A1 (n_1667), .A2 (n_1646));
NOR2_X1 i_250 (.ZN (n_1282), .A1 (n_1667), .A2 (n_1647));
NOR2_X1 i_249 (.ZN (n_1281), .A1 (n_1667), .A2 (n_1648));
NOR2_X1 i_248 (.ZN (n_1280), .A1 (n_1667), .A2 (n_1649));
NOR2_X1 i_247 (.ZN (n_729), .A1 (n_1667), .A2 (n_1650));
NOR2_X1 i_246 (.ZN (n_1274), .A1 (n_1668), .A2 (n_1625));
NOR2_X1 i_767 (.ZN (n_1273), .A1 (n_1668), .A2 (n_1628));
NOR2_X1 i_245 (.ZN (n_705), .A1 (n_1668), .A2 (n_1629));
NOR2_X1 i_244 (.ZN (n_1262), .A1 (n_1668), .A2 (n_1643));
NOR2_X1 i_243 (.ZN (n_1261), .A1 (n_1668), .A2 (n_1644));
NOR2_X1 i_242 (.ZN (n_1260), .A1 (n_1668), .A2 (n_1645));
NOR2_X1 i_241 (.ZN (n_1259), .A1 (n_1668), .A2 (n_1646));
NOR2_X1 i_240 (.ZN (n_1258), .A1 (n_1668), .A2 (n_1647));
NOR2_X1 i_239 (.ZN (n_1257), .A1 (n_1668), .A2 (n_1648));
NOR2_X1 i_238 (.ZN (n_704), .A1 (n_1668), .A2 (n_1649));
NOR2_X1 i_744 (.ZN (n_1250), .A1 (n_1669), .A2 (n_1625));
NOR2_X1 i_237 (.ZN (n_703), .A1 (n_1669), .A2 (n_1628));
NOR2_X1 i_236 (.ZN (n_1239), .A1 (n_1669), .A2 (n_1642));
NOR2_X1 i_235 (.ZN (n_1238), .A1 (n_1669), .A2 (n_1643));
NOR2_X1 i_234 (.ZN (n_1237), .A1 (n_1669), .A2 (n_1644));
NOR2_X1 i_233 (.ZN (n_1236), .A1 (n_1669), .A2 (n_1645));
NOR2_X1 i_232 (.ZN (n_1235), .A1 (n_1669), .A2 (n_1646));
NOR2_X1 i_231 (.ZN (n_1234), .A1 (n_1669), .A2 (n_1647));
NOR2_X1 i_230 (.ZN (n_702), .A1 (n_1669), .A2 (n_1648));
NOR2_X1 i_229 (.ZN (n_700), .A1 (n_1670), .A2 (n_1625));
NOR2_X1 i_228 (.ZN (n_1216), .A1 (n_1670), .A2 (n_1641));
NOR2_X1 i_227 (.ZN (n_1215), .A1 (n_1670), .A2 (n_1642));
NOR2_X1 i_226 (.ZN (n_1214), .A1 (n_1670), .A2 (n_1643));
NOR2_X1 i_225 (.ZN (n_1213), .A1 (n_1670), .A2 (n_1644));
NOR2_X1 i_224 (.ZN (n_1212), .A1 (n_1670), .A2 (n_1645));
NOR2_X1 i_223 (.ZN (n_1211), .A1 (n_1670), .A2 (n_1646));
NOR2_X1 i_222 (.ZN (n_669), .A1 (n_1670), .A2 (n_1647));
NOR2_X1 i_221 (.ZN (n_1193), .A1 (n_1672), .A2 (n_1640));
NOR2_X1 i_220 (.ZN (n_1192), .A1 (n_1672), .A2 (n_1641));
NOR2_X1 i_219 (.ZN (n_1191), .A1 (n_1672), .A2 (n_1642));
NOR2_X1 i_218 (.ZN (n_1190), .A1 (n_1672), .A2 (n_1643));
NOR2_X1 i_217 (.ZN (n_1189), .A1 (n_1672), .A2 (n_1644));
NOR2_X1 i_216 (.ZN (n_1188), .A1 (n_1672), .A2 (n_1645));
NOR2_X1 i_215 (.ZN (n_668), .A1 (n_1672), .A2 (n_1646));
NOR2_X1 i_214 (.ZN (n_1170), .A1 (n_1673), .A2 (n_1639));
NOR2_X1 i_213 (.ZN (n_1169), .A1 (n_1673), .A2 (n_1640));
NOR2_X1 i_212 (.ZN (n_1168), .A1 (n_1673), .A2 (n_1641));
NOR2_X1 i_211 (.ZN (n_1167), .A1 (n_1673), .A2 (n_1642));
NOR2_X1 i_210 (.ZN (n_1166), .A1 (n_1673), .A2 (n_1643));
NOR2_X1 i_209 (.ZN (n_1165), .A1 (n_1673), .A2 (n_1644));
NOR2_X1 i_208 (.ZN (n_667), .A1 (n_1673), .A2 (n_1645));
NOR2_X1 i_207 (.ZN (n_1147), .A1 (n_1674), .A2 (n_1634));
NOR2_X1 i_206 (.ZN (n_1146), .A1 (n_1674), .A2 (n_1639));
NOR2_X1 i_205 (.ZN (n_1145), .A1 (n_1674), .A2 (n_1640));
NOR2_X1 i_204 (.ZN (n_1144), .A1 (n_1674), .A2 (n_1641));
NOR2_X1 i_203 (.ZN (n_1143), .A1 (n_1674), .A2 (n_1642));
NOR2_X1 i_202 (.ZN (n_1142), .A1 (n_1674), .A2 (n_1643));
NOR2_X1 i_201 (.ZN (n_1141), .A1 (n_1674), .A2 (n_1644));
NOR2_X1 i_200 (.ZN (n_1124), .A1 (n_1675), .A2 (n_1633));
NOR2_X1 i_199 (.ZN (n_1123), .A1 (n_1675), .A2 (n_1634));
NOR2_X1 i_198 (.ZN (n_1122), .A1 (n_1675), .A2 (n_1639));
NOR2_X1 i_197 (.ZN (n_1121), .A1 (n_1675), .A2 (n_1640));
NOR2_X1 i_196 (.ZN (n_1120), .A1 (n_1675), .A2 (n_1641));
NOR2_X1 i_195 (.ZN (n_1119), .A1 (n_1675), .A2 (n_1642));
NOR2_X1 i_194 (.ZN (n_1118), .A1 (n_1675), .A2 (n_1643));
NOR2_X1 i_193 (.ZN (n_1101), .A1 (n_1676), .A2 (n_1632));
NOR2_X1 i_192 (.ZN (n_1100), .A1 (n_1676), .A2 (n_1633));
NOR2_X1 i_191 (.ZN (n_1099), .A1 (n_1676), .A2 (n_1634));
NOR2_X1 i_190 (.ZN (n_1098), .A1 (n_1676), .A2 (n_1639));
NOR2_X1 i_189 (.ZN (n_1097), .A1 (n_1676), .A2 (n_1640));
NOR2_X1 i_188 (.ZN (n_1096), .A1 (n_1676), .A2 (n_1641));
NOR2_X1 i_187 (.ZN (n_1095), .A1 (n_1676), .A2 (n_1642));
NOR2_X1 i_186 (.ZN (n_1078), .A1 (n_1677), .A2 (n_1631));
NOR2_X1 i_185 (.ZN (n_1077), .A1 (n_1677), .A2 (n_1632));
NOR2_X1 i_184 (.ZN (n_1076), .A1 (n_1677), .A2 (n_1633));
NOR2_X1 i_183 (.ZN (n_1075), .A1 (n_1677), .A2 (n_1634));
NOR2_X1 i_182 (.ZN (n_1074), .A1 (n_1677), .A2 (n_1639));
NOR2_X1 i_181 (.ZN (n_1073), .A1 (n_1677), .A2 (n_1640));
NOR2_X1 i_180 (.ZN (n_1072), .A1 (n_1677), .A2 (n_1641));
NOR2_X1 i_179 (.ZN (n_1055), .A1 (n_1678), .A2 (n_1630));
NOR2_X1 i_178 (.ZN (n_1054), .A1 (n_1678), .A2 (n_1631));
NOR2_X1 i_177 (.ZN (n_1053), .A1 (n_1678), .A2 (n_1632));
NOR2_X1 i_176 (.ZN (n_1052), .A1 (n_1678), .A2 (n_1633));
NOR2_X1 i_175 (.ZN (n_1051), .A1 (n_1678), .A2 (n_1634));
NOR2_X1 i_174 (.ZN (n_1050), .A1 (n_1678), .A2 (n_1639));
NOR2_X1 i_173 (.ZN (n_1049), .A1 (n_1678), .A2 (n_1640));
NOR2_X1 i_172 (.ZN (n_1032), .A1 (n_1654), .A2 (n_1629));
NOR2_X1 i_171 (.ZN (n_1031), .A1 (n_1654), .A2 (n_1630));
NOR2_X1 i_170 (.ZN (n_1030), .A1 (n_1654), .A2 (n_1631));
NOR2_X1 i_169 (.ZN (n_1029), .A1 (n_1654), .A2 (n_1632));
NOR2_X1 i_168 (.ZN (n_1028), .A1 (n_1654), .A2 (n_1633));
NOR2_X1 i_167 (.ZN (n_1027), .A1 (n_1654), .A2 (n_1634));
NOR2_X1 i_166 (.ZN (n_1026), .A1 (n_1654), .A2 (n_1639));
FA_X1 i_165 (.CO (n_666), .S (n_664), .A (n_782), .B (n_759), .CI (n_757));
FA_X1 i_164 (.CO (n_631), .S (n_629), .A (n_772), .B (n_755), .CI (n_784));
FA_X1 i_163 (.CO (n_549), .S (n_548), .A (n_1690), .B (n_1691), .CI (n_774));
FA_X1 i_162 (.CO (n_547), .S (n_545), .A (n_753), .B (n_751), .CI (n_1688));
FA_X1 i_161 (.CO (n_543), .S (n_784), .A (n_745), .B (n_743), .CI (n_741));
FA_X1 i_160 (.CO (n_541), .S (n_782), .A (n_1371), .B (n_749), .CI (n_747));
FA_X1 i_159 (.CO (n_539), .S (n_774), .A (n_1095), .B (n_1118), .CI (n_1141));
FA_X1 i_158 (.CO (n_537), .S (n_772), .A (n_1026), .B (n_1049), .CI (n_1072));
FA_X1 i_157 (.CO (n_535), .S (n_533), .A (n_733), .B (n_1700), .CI (n_735));
FA_X1 i_156 (.CO (n_531), .S (n_529), .A (n_725), .B (n_723), .CI (n_727));
FA_X1 i_155 (.CO (n_527), .S (n_525), .A (n_740), .B (n_754), .CI (n_752));
FA_X1 i_154 (.CO (n_759), .S (n_523), .A (n_746), .B (n_744), .CI (n_742));
FA_X1 i_153 (.CO (n_757), .S (n_521), .A (n_719), .B (n_750), .CI (n_748));
FA_X1 i_152 (.CO (n_755), .S (n_754), .A (n_709), .B (n_707), .CI (n_721));
FA_X1 i_151 (.CO (n_753), .S (n_752), .A (n_715), .B (n_713), .CI (n_711));
FA_X1 i_150 (.CO (n_751), .S (n_750), .A (n_1372), .B (n_1395), .CI (n_717));
FA_X1 i_149 (.CO (n_749), .S (n_748), .A (n_1303), .B (n_1326), .CI (n_1349));
FA_X1 i_148 (.CO (n_747), .S (n_746), .A (n_1234), .B (n_1257), .CI (n_1280));
FA_X1 i_147 (.CO (n_745), .S (n_744), .A (n_1165), .B (n_1188), .CI (n_1211));
FA_X1 i_146 (.CO (n_743), .S (n_742), .A (n_1096), .B (n_1119), .CI (n_1142));
FA_X1 i_145 (.CO (n_741), .S (n_740), .A (n_1027), .B (n_1050), .CI (n_1073));
FA_X1 i_144 (.CO (n_519), .S (n_517), .A (n_699), .B (n_732), .CI (n_701));
FA_X1 i_143 (.CO (n_735), .S (n_515), .A (n_728), .B (n_697), .CI (n_730));
FA_X1 i_142 (.CO (n_733), .S (n_732), .A (n_693), .B (n_726), .CI (n_724));
FA_X1 i_141 (.CO (n_513), .S (n_730), .A (n_689), .B (n_722), .CI (n_695));
FA_X1 i_140 (.CO (n_511), .S (n_728), .A (n_720), .B (n_718), .CI (n_691));
FA_X1 i_139 (.CO (n_727), .S (n_726), .A (n_708), .B (n_706), .CI (n_687));
FA_X1 i_138 (.CO (n_725), .S (n_724), .A (n_714), .B (n_712), .CI (n_710));
FA_X1 i_137 (.CO (n_723), .S (n_722), .A (n_685), .B (n_683), .CI (n_716));
FA_X1 i_136 (.CO (n_721), .S (n_720), .A (n_675), .B (n_673), .CI (n_671));
FA_X1 i_135 (.CO (n_719), .S (n_718), .A (n_681), .B (n_679), .CI (n_677));
FA_X1 i_134 (.CO (n_717), .S (n_716), .A (n_1373), .B (n_1396), .CI (n_1419));
FA_X1 i_133 (.CO (n_715), .S (n_714), .A (n_1304), .B (n_1327), .CI (n_1350));
FA_X1 i_132 (.CO (n_713), .S (n_712), .A (n_1235), .B (n_1258), .CI (n_1281));
FA_X1 i_131 (.CO (n_711), .S (n_710), .A (n_1166), .B (n_1189), .CI (n_1212));
FA_X1 i_130 (.CO (n_709), .S (n_708), .A (n_1097), .B (n_1120), .CI (n_1143));
FA_X1 i_129 (.CO (n_707), .S (n_706), .A (n_1028), .B (n_1051), .CI (n_1074));
FA_X1 i_128 (.CO (n_509), .S (n_507), .A (n_663), .B (n_698), .CI (n_665));
FA_X1 i_127 (.CO (n_701), .S (n_505), .A (n_692), .B (n_661), .CI (n_696));
FA_X1 i_126 (.CO (n_699), .S (n_698), .A (n_688), .B (n_659), .CI (n_694));
FA_X1 i_125 (.CO (n_697), .S (n_696), .A (n_686), .B (n_657), .CI (n_690));
FA_X1 i_124 (.CO (n_695), .S (n_694), .A (n_655), .B (n_653), .CI (n_651));
FA_X1 i_123 (.CO (n_693), .S (n_692), .A (n_670), .B (n_684), .CI (n_682));
FA_X1 i_122 (.CO (n_691), .S (n_690), .A (n_676), .B (n_674), .CI (n_672));
FA_X1 i_121 (.CO (n_689), .S (n_688), .A (n_645), .B (n_680), .CI (n_678));
FA_X1 i_120 (.CO (n_687), .S (n_686), .A (n_633), .B (n_649), .CI (n_647));
FA_X1 i_119 (.CO (n_685), .S (n_684), .A (n_639), .B (n_637), .CI (n_635));
FA_X1 i_118 (.CO (n_683), .S (n_682), .A (n_1443), .B (n_643), .CI (n_641));
FA_X1 i_117 (.CO (n_681), .S (n_680), .A (n_1374), .B (n_1397), .CI (n_1420));
FA_X1 i_116 (.CO (n_679), .S (n_678), .A (n_1305), .B (n_1328), .CI (n_1351));
FA_X1 i_115 (.CO (n_677), .S (n_676), .A (n_1236), .B (n_1259), .CI (n_1282));
FA_X1 i_114 (.CO (n_675), .S (n_674), .A (n_1167), .B (n_1190), .CI (n_1213));
FA_X1 i_113 (.CO (n_673), .S (n_672), .A (n_1098), .B (n_1121), .CI (n_1144));
FA_X1 i_112 (.CO (n_671), .S (n_670), .A (n_1029), .B (n_1052), .CI (n_1075));
FA_X1 i_111 (.CO (n_504), .S (n_461), .A (n_625), .B (n_662), .CI (n_627));
FA_X1 i_110 (.CO (n_665), .S (n_169), .A (n_656), .B (n_623), .CI (n_660));
FA_X1 i_109 (.CO (n_663), .S (n_662), .A (n_652), .B (n_621), .CI (n_658));
FA_X1 i_108 (.CO (n_661), .S (n_660), .A (n_619), .B (n_617), .CI (n_654));
FA_X1 i_107 (.CO (n_659), .S (n_658), .A (n_615), .B (n_613), .CI (n_650));
FA_X1 i_106 (.CO (n_657), .S (n_656), .A (n_611), .B (n_648), .CI (n_646));
FA_X1 i_105 (.CO (n_655), .S (n_654), .A (n_636), .B (n_634), .CI (n_632));
FA_X1 i_104 (.CO (n_653), .S (n_652), .A (n_642), .B (n_640), .CI (n_638));
FA_X1 i_103 (.CO (n_651), .S (n_650), .A (n_609), .B (n_607), .CI (n_644));
FA_X1 i_102 (.CO (n_649), .S (n_648), .A (n_597), .B (n_595), .CI (n_593));
FA_X1 i_101 (.CO (n_647), .S (n_646), .A (n_603), .B (n_601), .CI (n_599));
FA_X1 i_100 (.CO (n_645), .S (n_644), .A (n_1444), .B (n_1467), .CI (n_605));
FA_X1 i_99 (.CO (n_643), .S (n_642), .A (n_1375), .B (n_1398), .CI (n_1421));
FA_X1 i_98 (.CO (n_641), .S (n_640), .A (n_1306), .B (n_1329), .CI (n_1352));
FA_X1 i_97 (.CO (n_639), .S (n_638), .A (n_1237), .B (n_1260), .CI (n_1283));
FA_X1 i_96 (.CO (n_637), .S (n_636), .A (n_1168), .B (n_1191), .CI (n_1214));
FA_X1 i_95 (.CO (n_635), .S (n_634), .A (n_1099), .B (n_1122), .CI (n_1145));
FA_X1 i_94 (.CO (n_633), .S (n_632), .A (n_1030), .B (n_1053), .CI (n_1076));
FA_X1 i_93 (.CO (n_168), .S (n_630), .A (n_626), .B (n_589), .CI (n_628));
FA_X1 i_92 (.CO (n_167), .S (n_628), .A (n_622), .B (n_624), .CI (n_587));
FA_X1 i_91 (.CO (n_627), .S (n_626), .A (n_583), .B (n_620), .CI (n_585));
FA_X1 i_90 (.CO (n_625), .S (n_624), .A (n_616), .B (n_581), .CI (n_618));
FA_X1 i_89 (.CO (n_623), .S (n_622), .A (n_577), .B (n_614), .CI (n_612));
FA_X1 i_88 (.CO (n_621), .S (n_620), .A (n_571), .B (n_610), .CI (n_579));
FA_X1 i_87 (.CO (n_619), .S (n_618), .A (n_606), .B (n_575), .CI (n_573));
FA_X1 i_86 (.CO (n_617), .S (n_616), .A (n_592), .B (n_569), .CI (n_608));
FA_X1 i_85 (.CO (n_615), .S (n_614), .A (n_598), .B (n_596), .CI (n_594));
FA_X1 i_84 (.CO (n_613), .S (n_612), .A (n_604), .B (n_602), .CI (n_600));
FA_X1 i_83 (.CO (n_611), .S (n_610), .A (n_551), .B (n_567), .CI (n_565));
FA_X1 i_82 (.CO (n_609), .S (n_608), .A (n_557), .B (n_555), .CI (n_553));
FA_X1 i_81 (.CO (n_607), .S (n_606), .A (n_563), .B (n_561), .CI (n_559));
FA_X1 i_80 (.CO (n_605), .S (n_604), .A (n_1445), .B (n_1468), .CI (n_1491));
FA_X1 i_79 (.CO (n_603), .S (n_602), .A (n_1376), .B (n_1399), .CI (n_1422));
FA_X1 i_78 (.CO (n_601), .S (n_600), .A (n_1307), .B (n_1330), .CI (n_1353));
FA_X1 i_77 (.CO (n_599), .S (n_598), .A (n_1238), .B (n_1261), .CI (n_1284));
FA_X1 i_76 (.CO (n_597), .S (n_596), .A (n_1169), .B (n_1192), .CI (n_1215));
FA_X1 i_75 (.CO (n_595), .S (n_594), .A (n_1100), .B (n_1123), .CI (n_1146));
FA_X1 i_74 (.CO (n_593), .S (n_592), .A (n_1031), .B (n_1054), .CI (n_1077));
FA_X1 i_73 (.CO (n_591), .S (n_590), .A (n_586), .B (n_588), .CI (n_879));
FA_X1 i_72 (.CO (n_589), .S (n_588), .A (n_582), .B (n_584), .CI (n_878));
FA_X1 i_71 (.CO (n_587), .S (n_586), .A (n_580), .B (n_855), .CI (n_783));
FA_X1 i_70 (.CO (n_585), .S (n_584), .A (n_578), .B (n_576), .CI (n_792));
FA_X1 i_69 (.CO (n_583), .S (n_582), .A (n_574), .B (n_572), .CI (n_854));
FA_X1 i_68 (.CO (n_581), .S (n_580), .A (n_787), .B (n_570), .CI (n_780));
FA_X1 i_67 (.CO (n_579), .S (n_578), .A (n_564), .B (n_791), .CI (n_828));
FA_X1 i_66 (.CO (n_577), .S (n_576), .A (n_829), .B (n_568), .CI (n_566));
FA_X1 i_65 (.CO (n_575), .S (n_574), .A (n_554), .B (n_552), .CI (n_550));
FA_X1 i_64 (.CO (n_573), .S (n_572), .A (n_560), .B (n_558), .CI (n_556));
FA_X1 i_63 (.CO (n_571), .S (n_570), .A (n_778), .B (n_793), .CI (n_562));
FA_X1 i_62 (.CO (n_569), .S (n_568), .A (n_785), .B (n_786), .CI (n_776));
FA_X1 i_61 (.CO (n_567), .S (n_566), .A (n_788), .B (n_789), .CI (n_790));
FA_X1 i_60 (.CO (n_565), .S (n_564), .A (n_1515), .B (n_800), .CI (n_801));
FA_X1 i_59 (.CO (n_563), .S (n_562), .A (n_1446), .B (n_1469), .CI (n_1492));
FA_X1 i_58 (.CO (n_561), .S (n_560), .A (n_1377), .B (n_1400), .CI (n_1423));
FA_X1 i_55 (.CO (n_559), .S (n_558), .A (n_1308), .B (n_1331), .CI (n_1354));
FA_X1 i_54 (.CO (n_557), .S (n_556), .A (n_1239), .B (n_1262), .CI (n_1285));
FA_X1 i_53 (.CO (n_555), .S (n_554), .A (n_1170), .B (n_1193), .CI (n_1216));
FA_X1 i_52 (.CO (n_553), .S (n_552), .A (n_1101), .B (n_1124), .CI (n_1147));
FA_X1 i_51 (.CO (n_551), .S (n_550), .A (n_1032), .B (n_1055), .CI (n_1078));
FA_X1 i_50 (.CO (n_166), .S (n_165), .A (n_133), .B (n_939), .CI (n_141));
FA_X1 i_49 (.CO (n_164), .S (n_163), .A (n_139), .B (n_137), .CI (n_135));
FA_X1 i_44 (.CO (n_162), .S (n_161), .A (n_1526), .B (n_1549), .CI (n_1570));
FA_X1 i_43 (.CO (n_160), .S (n_159), .A (n_1457), .B (n_1480), .CI (n_1503));
FA_X1 i_42 (.CO (n_158), .S (n_157), .A (n_1388), .B (n_1411), .CI (n_1434));
FA_X1 i_41 (.CO (n_156), .S (n_143), .A (n_1319), .B (n_1342), .CI (n_1365));
FA_X1 i_40 (.CO (n_140), .S (n_138), .A (n_1250), .B (n_1273), .CI (n_1296));
FA_X1 i_39 (.CO (n_141), .S (n_136), .A (n_1550), .B (n_1571), .CI (n_117));
FA_X1 i_38 (.CO (n_139), .S (n_134), .A (n_1481), .B (n_1504), .CI (n_1527));
FA_X1 i_37 (.CO (n_137), .S (n_132), .A (n_1412), .B (n_1435), .CI (n_1458));
FA_X1 i_36 (.CO (n_135), .S (n_119), .A (n_1343), .B (n_1366), .CI (n_1389));
FA_X1 i_35 (.CO (n_133), .S (n_118), .A (n_1274), .B (n_1297), .CI (n_1320));
FA_X1 i_34 (.CO (n_116), .S (n_115), .A (n_1572), .B (n_97), .CI (n_95));
FA_X1 i_33 (.CO (n_117), .S (n_114), .A (n_1505), .B (n_1528), .CI (n_1551));
FA_X1 i_57 (.CO (n_113), .S (n_112), .A (n_1436), .B (n_1459), .CI (n_1482));
FA_X1 i_56 (.CO (n_111), .S (n_110), .A (n_1367), .B (n_1390), .CI (n_1413));
FA_X1 i_32 (.CO (n_99), .S (n_98), .A (n_1298), .B (n_1321), .CI (n_1344));
FA_X1 i_31 (.CO (n_96), .S (n_94), .A (n_77), .B (n_75), .CI (n_73));
FA_X1 i_48 (.CO (n_97), .S (n_93), .A (n_1529), .B (n_1552), .CI (n_1573));
FA_X1 i_47 (.CO (n_95), .S (n_92), .A (n_1460), .B (n_1483), .CI (n_1506));
FA_X1 i_46 (.CO (n_91), .S (n_90), .A (n_1391), .B (n_1414), .CI (n_1437));
FA_X1 i_45 (.CO (n_85), .S (n_84), .A (n_1322), .B (n_1345), .CI (n_1368));
FA_X1 i_30 (.CO (n_83), .S (n_82), .A (n_72), .B (n_80), .CI (n_65));
FA_X1 i_29 (.CO (n_81), .S (n_79), .A (n_78), .B (n_76), .CI (n_74));
FA_X1 i_28 (.CO (n_67), .S (n_80), .A (n_59), .B (n_57), .CI (n_63));
FA_X1 i_27 (.CO (n_66), .S (n_78), .A (n_1553), .B (n_1574), .CI (n_61));
FA_X1 i_26 (.CO (n_77), .S (n_76), .A (n_1484), .B (n_1507), .CI (n_1530));
FA_X1 i_25 (.CO (n_75), .S (n_74), .A (n_1415), .B (n_1438), .CI (n_1461));
FA_X1 i_24 (.CO (n_73), .S (n_72), .A (n_1346), .B (n_1369), .CI (n_1392));
FA_X1 i_23 (.CO (n_64), .S (n_51), .A (n_56), .B (n_49), .CI (n_62));
FA_X1 i_22 (.CO (n_65), .S (n_50), .A (n_43), .B (n_60), .CI (n_58));
FA_X1 i_21 (.CO (n_63), .S (n_62), .A (n_1575), .B (n_47), .CI (n_45));
FA_X1 i_20 (.CO (n_61), .S (n_60), .A (n_1508), .B (n_1531), .CI (n_1554));
FA_X1 i_19 (.CO (n_59), .S (n_58), .A (n_1439), .B (n_1462), .CI (n_1485));
FA_X1 i_18 (.CO (n_57), .S (n_56), .A (n_1370), .B (n_1393), .CI (n_1416));
FA_X1 i_17 (.CO (n_48), .S (n_37), .A (n_46), .B (n_44), .CI (n_42));
FA_X1 i_16 (.CO (n_49), .S (n_36), .A (n_33), .B (n_31), .CI (n_35));
FA_X1 i_15 (.CO (n_47), .S (n_46), .A (n_1532), .B (n_1555), .CI (n_1576));
FA_X1 i_14 (.CO (n_45), .S (n_44), .A (n_1463), .B (n_1486), .CI (n_1509));
FA_X1 i_13 (.CO (n_43), .S (n_42), .A (n_1394), .B (n_1417), .CI (n_1440));
FA_X1 i_12 (.CO (n_32), .S (n_30), .A (n_21), .B (n_25), .CI (n_34));
FA_X1 i_11 (.CO (n_35), .S (n_34), .A (n_1556), .B (n_1577), .CI (n_23));
FA_X1 i_10 (.CO (n_33), .S (n_24), .A (n_1487), .B (n_1510), .CI (n_1533));
FA_X1 i_9 (.CO (n_31), .S (n_22), .A (n_1418), .B (n_1441), .CI (n_1464));
FA_X1 i_8 (.CO (n_25), .S (n_20), .A (n_1578), .B (n_15), .CI (n_13));
FA_X1 i_7 (.CO (n_23), .S (n_14), .A (n_1511), .B (n_1534), .CI (n_1557));
FA_X1 i_6 (.CO (n_21), .S (n_12), .A (n_1442), .B (n_1465), .CI (n_1488));
FA_X1 i_5 (.CO (n_15), .S (n_10), .A (n_1535), .B (n_1558), .CI (n_1579));
FA_X1 i_4 (.CO (n_13), .S (n_9), .A (n_1466), .B (n_1489), .CI (n_1512));
FA_X1 i_3 (.CO (n_8), .S (n_6), .A (n_1559), .B (n_1580), .CI (n_5));
HA_X1 i_2 (.CO (n_5), .S (n_4), .A (n_1581), .B (n_1));
FA_X1 i_1 (.CO (n_3), .S (n_2), .A (n_1514), .B (n_1537), .CI (n_1560));
HA_X1 i_0 (.CO (n_1), .S (n_0), .A (n_1538), .B (n_1723));
BUF_X2 hfn_ipo_c6 (.Z (hfn_ipo_n6), .A (n_1654));

endmodule //datapath__0_2

module VM (clk_CTS_0_PP_4, clk_CTS_0_PP_5, clk_CTS_0_PP_6, Res, OVF, A, B, clk, reset, 
    enable);

output OVF;
output [63:0] Res;
output clk_CTS_0_PP_4;
output clk_CTS_0_PP_5;
input [31:0] A;
input [31:0] B;
input clk;
input enable;
input reset;
input clk_CTS_0_PP_6;
wire \Res_imm[47] ;
wire \Res_imm[46] ;
wire \Res_imm[45] ;
wire \Res_imm[44] ;
wire \Res_imm[43] ;
wire \Res_imm[42] ;
wire \Res_imm[41] ;
wire \Res_imm[40] ;
wire \Res_imm[39] ;
wire \Res_imm[38] ;
wire \Res_imm[37] ;
wire \Res_imm[36] ;
wire \Res_imm[35] ;
wire \Res_imm[34] ;
wire \Res_imm[33] ;
wire \Res_imm[32] ;
wire \Res_imm[31] ;
wire \Res_imm[30] ;
wire \Res_imm[29] ;
wire \Res_imm[28] ;
wire \Res_imm[27] ;
wire \Res_imm[26] ;
wire \Res_imm[25] ;
wire \Res_imm[24] ;
wire \Res_imm[23] ;
wire hfn_ipo_n6;
wire CTS_n12;
wire n_0_0__1;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire uc_8;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_0;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire n_46;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_1;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire uc_28;
wire uc_29;
wire uc_30;
wire uc_31;
wire uc_32;
wire uc_33;
wire uc_34;
wire uc_35;
wire uc_36;
wire uc_37;
wire uc_38;
wire uc_39;
wire uc_40;
wire uc_41;
wire uc_42;
wire uc_43;
wire uc_44;
wire uc_45;
wire uc_46;
wire uc_47;
wire uc_48;
wire uc_49;
wire uc_50;
wire uc_51;
wire uc_52;
wire uc_53;
wire uc_54;
wire uc_55;
wire n_71;
wire n_119;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_118;
wire CTS_n11;
wire n_117;
wire n_116;
wire n_115;
wire n_114;
wire n_113;
wire n_112;
wire n_111;
wire n_110;
wire n_109;
wire n_108;
wire n_107;
wire n_106;
wire n_105;
wire n_104;
wire n_103;
wire n_102;
wire n_101;
wire n_100;
wire n_99;
wire n_98;
wire n_97;
wire n_96;
wire n_94;
wire n_93;
wire n_92;
wire n_91;
wire n_90;
wire n_89;
wire n_88;
wire n_87;
wire n_86;
wire n_85;
wire n_84;
wire n_83;
wire n_82;
wire n_81;
wire n_80;
wire n_79;
wire n_78;
wire n_77;
wire n_76;
wire n_75;
wire n_74;
wire n_73;
wire n_72;


INV_X1 i_0_74 (.ZN (n_0_0__1), .A (reset));
NAND2_X2 i_0_73 (.ZN (n_119), .A1 (n_0_0__1), .A2 (clk_CTS_0_PP_4));
AND2_X1 i_0_72 (.ZN (n_118), .A1 (hfn_ipo_n6), .A2 (B[22]));
AND2_X1 i_0_71 (.ZN (n_117), .A1 (hfn_ipo_n6), .A2 (B[21]));
AND2_X1 i_0_70 (.ZN (n_116), .A1 (hfn_ipo_n6), .A2 (B[20]));
AND2_X1 i_0_69 (.ZN (n_115), .A1 (hfn_ipo_n6), .A2 (B[19]));
AND2_X1 i_0_68 (.ZN (n_114), .A1 (hfn_ipo_n6), .A2 (B[18]));
AND2_X1 i_0_67 (.ZN (n_113), .A1 (hfn_ipo_n6), .A2 (B[17]));
AND2_X1 i_0_66 (.ZN (n_112), .A1 (hfn_ipo_n6), .A2 (B[16]));
AND2_X1 i_0_65 (.ZN (n_111), .A1 (hfn_ipo_n6), .A2 (B[15]));
AND2_X1 i_0_64 (.ZN (n_110), .A1 (hfn_ipo_n6), .A2 (B[14]));
AND2_X1 i_0_63 (.ZN (n_109), .A1 (hfn_ipo_n6), .A2 (B[13]));
AND2_X1 i_0_62 (.ZN (n_108), .A1 (hfn_ipo_n6), .A2 (B[12]));
AND2_X1 i_0_61 (.ZN (n_107), .A1 (hfn_ipo_n6), .A2 (B[11]));
AND2_X1 i_0_60 (.ZN (n_106), .A1 (hfn_ipo_n6), .A2 (B[10]));
AND2_X1 i_0_59 (.ZN (n_105), .A1 (hfn_ipo_n6), .A2 (B[9]));
AND2_X1 i_0_58 (.ZN (n_104), .A1 (hfn_ipo_n6), .A2 (B[8]));
AND2_X1 i_0_57 (.ZN (n_103), .A1 (hfn_ipo_n6), .A2 (B[7]));
AND2_X1 i_0_56 (.ZN (n_102), .A1 (hfn_ipo_n6), .A2 (B[6]));
AND2_X1 i_0_55 (.ZN (n_101), .A1 (hfn_ipo_n6), .A2 (B[5]));
AND2_X1 i_0_54 (.ZN (n_100), .A1 (hfn_ipo_n6), .A2 (B[4]));
AND2_X1 i_0_53 (.ZN (n_99), .A1 (hfn_ipo_n6), .A2 (B[3]));
AND2_X1 i_0_52 (.ZN (n_98), .A1 (hfn_ipo_n6), .A2 (B[2]));
AND2_X1 i_0_51 (.ZN (n_97), .A1 (hfn_ipo_n6), .A2 (B[1]));
AND2_X1 i_0_50 (.ZN (n_96), .A1 (hfn_ipo_n6), .A2 (B[0]));
AOI21_X1 i_0_49 (.ZN (CTS_n12), .A (reset), .B1 (clk_CTS_0_PP_4), .B2 (enable));
INV_X4 CTS_L4_remove_c14 (.ZN (CTS_n11), .A (CTS_n12));
AND2_X1 i_0_47 (.ZN (n_94), .A1 (hfn_ipo_n6), .A2 (A[22]));
AND2_X1 i_0_46 (.ZN (n_93), .A1 (hfn_ipo_n6), .A2 (A[21]));
AND2_X1 i_0_45 (.ZN (n_92), .A1 (hfn_ipo_n6), .A2 (A[20]));
AND2_X1 i_0_44 (.ZN (n_91), .A1 (hfn_ipo_n6), .A2 (A[19]));
AND2_X1 i_0_43 (.ZN (n_90), .A1 (hfn_ipo_n6), .A2 (A[18]));
AND2_X1 i_0_42 (.ZN (n_89), .A1 (hfn_ipo_n6), .A2 (A[17]));
AND2_X1 i_0_41 (.ZN (n_88), .A1 (hfn_ipo_n6), .A2 (A[16]));
AND2_X1 i_0_40 (.ZN (n_87), .A1 (hfn_ipo_n6), .A2 (A[15]));
AND2_X1 i_0_39 (.ZN (n_86), .A1 (hfn_ipo_n6), .A2 (A[14]));
AND2_X1 i_0_38 (.ZN (n_85), .A1 (hfn_ipo_n6), .A2 (A[13]));
AND2_X1 i_0_37 (.ZN (n_84), .A1 (hfn_ipo_n6), .A2 (A[12]));
AND2_X1 i_0_36 (.ZN (n_83), .A1 (hfn_ipo_n6), .A2 (A[11]));
AND2_X1 i_0_35 (.ZN (n_82), .A1 (hfn_ipo_n6), .A2 (A[10]));
AND2_X1 i_0_34 (.ZN (n_81), .A1 (hfn_ipo_n6), .A2 (A[9]));
AND2_X1 i_0_33 (.ZN (n_80), .A1 (hfn_ipo_n6), .A2 (A[8]));
AND2_X1 i_0_32 (.ZN (n_79), .A1 (hfn_ipo_n6), .A2 (A[7]));
AND2_X1 i_0_31 (.ZN (n_78), .A1 (hfn_ipo_n6), .A2 (A[6]));
AND2_X1 i_0_30 (.ZN (n_77), .A1 (hfn_ipo_n6), .A2 (A[5]));
AND2_X1 i_0_29 (.ZN (n_76), .A1 (hfn_ipo_n6), .A2 (A[4]));
AND2_X1 i_0_28 (.ZN (n_75), .A1 (hfn_ipo_n6), .A2 (A[3]));
AND2_X1 i_0_27 (.ZN (n_74), .A1 (hfn_ipo_n6), .A2 (A[2]));
AND2_X1 i_0_26 (.ZN (n_73), .A1 (hfn_ipo_n6), .A2 (A[1]));
AND2_X1 i_0_25 (.ZN (n_72), .A1 (hfn_ipo_n6), .A2 (A[0]));
AND2_X1 i_0_24 (.ZN (n_71), .A1 (n_0_0__1), .A2 (\Res_imm[47] ));
AND2_X1 i_0_23 (.ZN (n_70), .A1 (n_0_0__1), .A2 (\Res_imm[46] ));
AND2_X1 i_0_22 (.ZN (n_69), .A1 (n_0_0__1), .A2 (\Res_imm[45] ));
AND2_X1 i_0_21 (.ZN (n_68), .A1 (n_0_0__1), .A2 (\Res_imm[44] ));
AND2_X1 i_0_20 (.ZN (n_67), .A1 (n_0_0__1), .A2 (\Res_imm[43] ));
AND2_X1 i_0_19 (.ZN (n_66), .A1 (n_0_0__1), .A2 (\Res_imm[42] ));
AND2_X1 i_0_18 (.ZN (n_65), .A1 (n_0_0__1), .A2 (\Res_imm[41] ));
AND2_X1 i_0_17 (.ZN (n_64), .A1 (n_0_0__1), .A2 (\Res_imm[40] ));
AND2_X1 i_0_16 (.ZN (n_63), .A1 (n_0_0__1), .A2 (\Res_imm[39] ));
AND2_X1 i_0_15 (.ZN (n_62), .A1 (n_0_0__1), .A2 (\Res_imm[38] ));
AND2_X1 i_0_14 (.ZN (n_61), .A1 (n_0_0__1), .A2 (\Res_imm[37] ));
AND2_X1 i_0_13 (.ZN (n_60), .A1 (n_0_0__1), .A2 (\Res_imm[36] ));
AND2_X1 i_0_12 (.ZN (n_59), .A1 (n_0_0__1), .A2 (\Res_imm[35] ));
AND2_X1 i_0_11 (.ZN (n_58), .A1 (n_0_0__1), .A2 (\Res_imm[34] ));
AND2_X1 i_0_10 (.ZN (n_57), .A1 (n_0_0__1), .A2 (\Res_imm[33] ));
AND2_X1 i_0_9 (.ZN (n_56), .A1 (n_0_0__1), .A2 (\Res_imm[32] ));
AND2_X1 i_0_8 (.ZN (n_55), .A1 (n_0_0__1), .A2 (\Res_imm[31] ));
AND2_X1 i_0_7 (.ZN (n_54), .A1 (n_0_0__1), .A2 (\Res_imm[30] ));
AND2_X1 i_0_6 (.ZN (n_53), .A1 (n_0_0__1), .A2 (\Res_imm[29] ));
AND2_X1 i_0_5 (.ZN (n_52), .A1 (n_0_0__1), .A2 (\Res_imm[28] ));
AND2_X1 i_0_4 (.ZN (n_51), .A1 (n_0_0__1), .A2 (\Res_imm[27] ));
AND2_X1 i_0_3 (.ZN (n_50), .A1 (n_0_0__1), .A2 (\Res_imm[26] ));
AND2_X1 i_0_2 (.ZN (n_49), .A1 (n_0_0__1), .A2 (\Res_imm[25] ));
AND2_X1 i_0_1 (.ZN (n_48), .A1 (n_0_0__1), .A2 (\Res_imm[24] ));
AND2_X1 i_0_0 (.ZN (n_47), .A1 (n_0_0__1), .A2 (\Res_imm[23] ));
DLH_X1 \A_in_reg[23]  (.Q (n_46), .D (hfn_ipo_n6), .G (CTS_n11));
DLH_X1 \A_in_reg[0]  (.Q (n_1), .D (n_72), .G (CTS_n11));
DLH_X1 \A_in_reg[1]  (.Q (n_45), .D (n_73), .G (CTS_n11));
DLH_X1 \A_in_reg[2]  (.Q (n_44), .D (n_74), .G (CTS_n11));
DLH_X1 \A_in_reg[3]  (.Q (n_43), .D (n_75), .G (CTS_n11));
DLH_X1 \A_in_reg[4]  (.Q (n_42), .D (n_76), .G (CTS_n11));
DLH_X1 \A_in_reg[5]  (.Q (n_41), .D (n_77), .G (CTS_n11));
DLH_X1 \A_in_reg[6]  (.Q (n_40), .D (n_78), .G (CTS_n11));
DLH_X1 \A_in_reg[7]  (.Q (n_39), .D (n_79), .G (CTS_n11));
DLH_X1 \A_in_reg[8]  (.Q (n_38), .D (n_80), .G (CTS_n11));
DLH_X1 \A_in_reg[9]  (.Q (n_37), .D (n_81), .G (CTS_n11));
DLH_X1 \A_in_reg[10]  (.Q (n_36), .D (n_82), .G (CTS_n11));
DLH_X1 \A_in_reg[11]  (.Q (n_35), .D (n_83), .G (CTS_n11));
DLH_X1 \A_in_reg[12]  (.Q (n_34), .D (n_84), .G (CTS_n11));
DLH_X1 \A_in_reg[13]  (.Q (n_33), .D (n_85), .G (CTS_n11));
DLH_X1 \A_in_reg[14]  (.Q (n_32), .D (n_86), .G (CTS_n11));
DLH_X1 \A_in_reg[15]  (.Q (n_31), .D (n_87), .G (CTS_n11));
DLH_X1 \A_in_reg[16]  (.Q (n_30), .D (n_88), .G (CTS_n11));
DLH_X1 \A_in_reg[17]  (.Q (n_29), .D (n_89), .G (CTS_n11));
DLH_X1 \A_in_reg[18]  (.Q (n_28), .D (n_90), .G (CTS_n11));
DLH_X1 \A_in_reg[19]  (.Q (n_27), .D (n_91), .G (CTS_n11));
DLH_X1 \A_in_reg[20]  (.Q (n_26), .D (n_92), .G (CTS_n11));
DLH_X1 \A_in_reg[21]  (.Q (n_25), .D (n_93), .G (CTS_n11));
DLH_X1 \A_in_reg[22]  (.Q (n_24), .D (n_94), .G (CTS_n11));
DLH_X1 \B_in_reg[0]  (.Q (n_0), .D (n_96), .G (CTS_n11));
DLH_X1 \B_in_reg[1]  (.Q (n_23), .D (n_97), .G (CTS_n11));
DLH_X1 \B_in_reg[2]  (.Q (n_22), .D (n_98), .G (CTS_n11));
DLH_X1 \B_in_reg[3]  (.Q (n_21), .D (n_99), .G (CTS_n11));
DLH_X1 \B_in_reg[4]  (.Q (n_20), .D (n_100), .G (CTS_n11));
DLH_X1 \B_in_reg[5]  (.Q (n_19), .D (n_101), .G (CTS_n11));
DLH_X1 \B_in_reg[6]  (.Q (n_18), .D (n_102), .G (CTS_n11));
DLH_X1 \B_in_reg[7]  (.Q (n_17), .D (n_103), .G (CTS_n11));
DLH_X1 \B_in_reg[8]  (.Q (n_16), .D (n_104), .G (CTS_n11));
DLH_X1 \B_in_reg[9]  (.Q (n_15), .D (n_105), .G (CTS_n11));
DLH_X1 \B_in_reg[10]  (.Q (n_14), .D (n_106), .G (CTS_n11));
DLH_X1 \B_in_reg[11]  (.Q (n_13), .D (n_107), .G (CTS_n11));
DLH_X1 \B_in_reg[12]  (.Q (n_12), .D (n_108), .G (CTS_n11));
DLH_X1 \B_in_reg[13]  (.Q (n_11), .D (n_109), .G (CTS_n11));
DLH_X1 \B_in_reg[14]  (.Q (n_10), .D (n_110), .G (CTS_n11));
DLH_X1 \B_in_reg[15]  (.Q (n_9), .D (n_111), .G (CTS_n11));
DLH_X1 \B_in_reg[16]  (.Q (n_8), .D (n_112), .G (CTS_n11));
DLH_X1 \B_in_reg[17]  (.Q (n_7), .D (n_113), .G (CTS_n11));
DLH_X1 \B_in_reg[18]  (.Q (n_6), .D (n_114), .G (CTS_n11));
DLH_X1 \B_in_reg[19]  (.Q (n_5), .D (n_115), .G (CTS_n11));
DLH_X1 \B_in_reg[20]  (.Q (n_4), .D (n_116), .G (CTS_n11));
DLH_X1 \B_in_reg[21]  (.Q (n_3), .D (n_117), .G (CTS_n11));
DLH_X1 \B_in_reg[22]  (.Q (n_2), .D (n_118), .G (CTS_n11));
DLH_X1 \Res_reg[23]  (.Q (Res[23]), .D (n_47), .G (n_119));
DLH_X1 \Res_reg[24]  (.Q (Res[24]), .D (n_48), .G (n_119));
DLH_X1 \Res_reg[25]  (.Q (Res[25]), .D (n_49), .G (n_119));
DLH_X1 \Res_reg[26]  (.Q (Res[26]), .D (n_50), .G (n_119));
DLH_X1 \Res_reg[27]  (.Q (Res[27]), .D (n_51), .G (n_119));
DLH_X1 \Res_reg[28]  (.Q (Res[28]), .D (n_52), .G (n_119));
DLH_X1 \Res_reg[29]  (.Q (Res[29]), .D (n_53), .G (n_119));
DLH_X1 \Res_reg[30]  (.Q (Res[30]), .D (n_54), .G (n_119));
DLH_X1 \Res_reg[31]  (.Q (Res[31]), .D (n_55), .G (n_119));
DLH_X1 \Res_reg[32]  (.Q (Res[32]), .D (n_56), .G (n_119));
DLH_X1 \Res_reg[33]  (.Q (Res[33]), .D (n_57), .G (n_119));
DLH_X1 \Res_reg[34]  (.Q (Res[34]), .D (n_58), .G (n_119));
DLH_X1 \Res_reg[35]  (.Q (Res[35]), .D (n_59), .G (n_119));
DLH_X1 \Res_reg[36]  (.Q (Res[36]), .D (n_60), .G (n_119));
DLH_X1 \Res_reg[37]  (.Q (Res[37]), .D (n_61), .G (n_119));
DLH_X1 \Res_reg[38]  (.Q (Res[38]), .D (n_62), .G (n_119));
DLH_X1 \Res_reg[39]  (.Q (Res[39]), .D (n_63), .G (n_119));
DLH_X1 \Res_reg[40]  (.Q (Res[40]), .D (n_64), .G (n_119));
DLH_X1 \Res_reg[41]  (.Q (Res[41]), .D (n_65), .G (n_119));
DLH_X1 \Res_reg[42]  (.Q (Res[42]), .D (n_66), .G (n_119));
DLH_X1 \Res_reg[43]  (.Q (Res[43]), .D (n_67), .G (n_119));
DLH_X1 \Res_reg[44]  (.Q (Res[44]), .D (n_68), .G (n_119));
DLH_X1 \Res_reg[45]  (.Q (Res[45]), .D (n_69), .G (n_119));
DLH_X1 \Res_reg[46]  (.Q (Res[46]), .D (n_70), .G (n_119));
DLH_X1 \Res_reg[47]  (.Q (Res[47]), .D (n_71), .G (n_119));
datapath__0_2 i_4 (.Res_imm ({uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, 
    uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, uc_32, \Res_imm[47] , \Res_imm[46] , 
    \Res_imm[45] , \Res_imm[44] , \Res_imm[43] , \Res_imm[42] , \Res_imm[41] , \Res_imm[40] , 
    \Res_imm[39] , \Res_imm[38] , \Res_imm[37] , \Res_imm[36] , \Res_imm[35] , \Res_imm[34] , 
    \Res_imm[33] , \Res_imm[32] , \Res_imm[31] , \Res_imm[30] , \Res_imm[29] , \Res_imm[28] , 
    \Res_imm[27] , \Res_imm[26] , \Res_imm[25] , \Res_imm[24] , \Res_imm[23] , uc_33, 
    uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, 
    uc_45, uc_46, uc_47, uc_48, uc_49, uc_50, uc_51, uc_52, uc_53, uc_54, uc_55})
    , .A_imm ({uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, n_46, n_24, 
    n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, 
    n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_1}), .B_imm ({uc_0, uc_1, uc_2, 
    uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, 
    n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, 
    n_0}));
CLKBUF_X3 CTS_L2_c_tid0_41 (.Z (clk_CTS_0_PP_4), .A (clk_CTS_0_PP_5));
CLKBUF_X3 hfn_ipo_c6 (.Z (hfn_ipo_n6), .A (n_0_0__1));
CLKBUF_X1 CTS_L1_c_tid0_42 (.Z (clk_CTS_0_PP_5), .A (clk_CTS_0_PP_6));

endmodule //VM

module FPU_VM (Res, A, B, clk, reset, enable);

output [31:0] Res;
input [31:0] A;
input [31:0] B;
input clk;
input enable;
input reset;
wire CTS_n_tid0_90;
wire CLOCK_slh__n413;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire \M_resultTruncated[22] ;
wire \M_resultTruncated[21] ;
wire \M_resultTruncated[20] ;
wire \M_resultTruncated[19] ;
wire \M_resultTruncated[18] ;
wire \M_resultTruncated[17] ;
wire \M_resultTruncated[16] ;
wire \M_resultTruncated[15] ;
wire \M_resultTruncated[14] ;
wire \M_resultTruncated[13] ;
wire \M_resultTruncated[12] ;
wire \M_resultTruncated[11] ;
wire \M_resultTruncated[10] ;
wire \M_resultTruncated[9] ;
wire \M_resultTruncated[8] ;
wire \M_resultTruncated[7] ;
wire \M_resultTruncated[6] ;
wire \M_resultTruncated[5] ;
wire \M_resultTruncated[4] ;
wire \M_resultTruncated[3] ;
wire \M_resultTruncated[2] ;
wire \M_resultTruncated[1] ;
wire \M_resultTruncated[0] ;
wire \EA[7] ;
wire \EA[6] ;
wire \EA[5] ;
wire \EA[4] ;
wire \EA[3] ;
wire \EA[2] ;
wire \EA[1] ;
wire \EA[0] ;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire \EB[7] ;
wire \EB[6] ;
wire \EB[5] ;
wire \EB[4] ;
wire \EB[3] ;
wire \EB[2] ;
wire \EB[1] ;
wire \EB[0] ;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire A_reg;
wire B_reg;
wire n_0_1_2;
wire n_0_1_3;
wire n_0_1_4;
wire n_0_1_5;
wire n_0_1_6;
wire n_0_1_7;
wire n_0_1_8;
wire n_0_1_9;
wire n_0_1_10;
wire n_0_1_11;
wire n_0_1_12;
wire n_0_1_13;
wire n_0_1_14;
wire n_0_1_15;
wire n_0_1_22;
wire n_0_1_16;
wire n_0_1_23;
wire n_0_1_17;
wire n_0_1_24;
wire n_0_1_18;
wire n_0_1_25;
wire n_0_1_19;
wire n_0_1_26;
wire n_0_1_20;
wire n_0_1_27;
wire n_0_1_21;
wire n_0_1_0;
wire n_0_1_1;
wire n_0_72;
wire n_0_1_32;
wire n_0_73;
wire n_0_1_33;
wire n_0_74;
wire n_0_1_34;
wire n_0_75;
wire n_0_1_35;
wire n_0_76;
wire n_0_1_36;
wire n_0_77;
wire n_0_1_37;
wire n_0_78;
wire n_0_1_38;
wire n_0_79;
wire n_0_1_39;
wire n_0_80;
wire n_0_1_40;
wire n_0_81;
wire n_0_1_41;
wire n_0_82;
wire n_0_1_42;
wire n_0_83;
wire n_0_1_43;
wire n_0_84;
wire n_0_1_44;
wire n_0_85;
wire n_0_1_45;
wire n_0_86;
wire n_0_1_46;
wire n_0_87;
wire n_0_1_47;
wire n_0_88;
wire n_0_1_48;
wire n_0_89;
wire n_0_1_49;
wire n_0_90;
wire n_0_1_50;
wire n_0_91;
wire n_0_1_51;
wire n_0_92;
wire n_0_1_52;
wire n_0_93;
wire n_0_1_53;
wire n_0_1_54;
wire n_0_1_55;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_1_56;
wire n_0_1_57;
wire n_0_1_58;
wire n_0_1_59;
wire n_0_1_60;
wire n_0_1_62;
wire n_0_1_64;
wire n_0_103;
wire CTS_n_tid0_13;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_1_105;
wire n_0_1_106;
wire n_0_1_107;
wire n_0_1_108;
wire n_0_1_109;
wire n_0_1_110;
wire n_0_1_111;
wire n_0_1_112;
wire n_0_1_28;
wire n_0_1_29;
wire n_0_71;
wire n_0_1_30;
wire n_0_1_31;
wire n_0_1_61;
wire n_0_1_63;
wire n_0_1_65;
wire n_0_1_66;
wire n_0_1_67;
wire n_0_1_68;
wire n_0_1_69;
wire n_0_1_70;
wire n_0_1_71;
wire n_0_1_72;
wire n_0_1_73;
wire n_0_1_74;
wire n_0_1_75;
wire n_0_1_76;
wire n_0_1_77;
wire n_0_1_78;
wire n_0_1_79;
wire n_0_1_80;
wire n_0_1_81;
wire n_0_1_82;
wire n_0_1_83;
wire n_0_1_84;
wire n_0_1_85;
wire n_0_1_86;
wire n_0_1_87;
wire n_0_1_88;
wire n_0_1_89;
wire n_0_1_90;
wire n_0_1_91;
wire n_0_1_92;
wire n_0_1_93;
wire n_0_1_94;
wire n_0_1_95;
wire n_0_1_96;
wire n_0_1_97;
wire n_0_1_98;
wire n_0_1_99;
wire n_0_1_100;
wire n_0_1_101;
wire n_0_1_102;
wire CTS_n_tid0_14;
wire n_0_102;
wire n_0_1_104;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire uc_28;
wire uc_29;
wire uc_30;
wire uc_31;
wire uc_32;
wire uc_33;
wire uc_34;
wire uc_35;
wire uc_36;
wire uc_37;
wire uc_38;
wire uc_39;
wire uc_40;
wire uc_41;
wire uc_42;
wire uc_43;
wire uc_44;
wire uc_45;
wire uc_46;
wire uc_47;
wire uc_48;
wire uc_49;
wire uc_50;
wire uc_51;
wire uc_52;
wire uc_53;
wire uc_54;
wire uc_55;
wire uc_56;
wire hfn_ipo_n10;
wire hfn_ipo_n11;
wire CLOCK_slh__n179;
wire CTS_n_tid0_91;
wire CLOCK_slh__n178;
wire CLOCK_slh__n182;
wire CLOCK_slh__n183;
wire CLOCK_slh__n186;
wire CLOCK_slh__n187;
wire CLOCK_slh__n190;
wire CLOCK_slh__n191;
wire CLOCK_slh__n194;
wire CLOCK_slh__n195;
wire CLOCK_slh__n198;
wire CLOCK_slh__n199;
wire CLOCK_slh__n202;
wire CLOCK_slh__n203;
wire CLOCK_slh__n206;
wire CLOCK_slh__n207;
wire CLOCK_slh__n210;
wire CLOCK_slh__n211;
wire CLOCK_slh__n214;
wire CLOCK_slh__n215;
wire CLOCK_slh__n218;
wire CLOCK_slh__n219;
wire CLOCK_slh__n222;
wire CLOCK_slh__n223;
wire CLOCK_slh__n226;
wire CLOCK_slh__n227;
wire CLOCK_slh__n230;
wire CLOCK_slh__n231;
wire CLOCK_slh__n234;
wire CLOCK_slh__n235;
wire CLOCK_slh__n238;
wire CLOCK_slh__n239;
wire CLOCK_slh__n242;
wire CLOCK_slh__n243;
wire CLOCK_slh__n246;
wire CLOCK_slh__n247;
wire CLOCK_slh__n250;
wire CLOCK_slh__n251;
wire CLOCK_slh__n254;
wire CLOCK_slh__n255;
wire CLOCK_slh__n258;
wire CLOCK_slh__n259;
wire CLOCK_slh__n262;
wire CLOCK_slh__n263;
wire CLOCK_slh__n266;
wire CLOCK_slh__n267;
wire CLOCK_slh__n270;
wire CLOCK_slh__n271;
wire CLOCK_slh__n274;
wire CLOCK_slh__n275;
wire CLOCK_slh__n278;
wire CLOCK_slh__n279;
wire CLOCK_slh__n282;
wire CLOCK_slh__n283;
wire CLOCK_slh__n286;
wire CLOCK_slh__n287;
wire CLOCK_slh__n290;
wire CLOCK_slh__n291;
wire CLOCK_slh__n294;
wire CLOCK_slh__n295;
wire CLOCK_slh__n298;
wire CLOCK_slh__n299;
wire CLOCK_slh__n302;
wire CLOCK_slh__n303;
wire CLOCK_slh__n306;
wire CLOCK_slh__n307;
wire CLOCK_slh__n310;
wire CLOCK_slh__n311;
wire CLOCK_slh__n314;
wire CLOCK_slh__n315;
wire CLOCK_slh__n318;
wire CLOCK_slh__n319;
wire CLOCK_slh__n322;
wire CLOCK_slh__n323;
wire CLOCK_slh__n326;
wire CLOCK_slh__n327;
wire CLOCK_slh__n330;
wire CLOCK_slh__n331;
wire CLOCK_slh__n334;
wire CLOCK_slh__n335;
wire CLOCK_slh__n338;
wire CLOCK_slh__n339;
wire CLOCK_slh__n342;
wire CLOCK_slh__n343;
wire CLOCK_slh__n346;
wire CLOCK_slh__n347;
wire CLOCK_slh__n350;
wire CLOCK_slh__n351;
wire CLOCK_slh__n354;
wire CLOCK_slh__n355;
wire CLOCK_slh__n358;
wire CLOCK_slh__n359;
wire CLOCK_slh__n362;
wire CLOCK_slh__n363;
wire CLOCK_slh__n366;
wire CLOCK_slh__n367;
wire CLOCK_slh__n370;
wire CLOCK_slh__n371;
wire CLOCK_slh__n374;
wire CLOCK_slh__n375;
wire CLOCK_slh__n378;
wire CLOCK_slh__n379;
wire CLOCK_slh__n382;
wire CLOCK_slh__n383;
wire CLOCK_slh__n386;
wire CLOCK_slh__n387;
wire CLOCK_slh__n390;
wire CLOCK_slh__n391;
wire CLOCK_slh__n392;
wire CLOCK_slh__n393;
wire CLOCK_slh__n394;
wire CLOCK_slh__n395;
wire CLOCK_slh__n396;
wire CLOCK_slh__n397;
wire CLOCK_slh__n398;
wire CLOCK_slh__n399;
wire CLOCK_slh__n400;
wire CLOCK_slh__n401;
wire CLOCK_slh__n402;
wire CLOCK_slh__n403;
wire CLOCK_slh__n404;
wire CLOCK_slh__n405;
wire CLOCK_slh__n406;
wire CLOCK_slh__n407;
wire CLOCK_slh__n408;
wire CLOCK_slh__n409;
wire CLOCK_slh__n410;
wire CLOCK_slh__n411;
wire CLOCK_slh__n414;
wire CLOCK_slh__n415;
wire CLOCK_slh__n416;
wire CLOCK_slh__n422;
wire CLOCK_slh__n423;
wire CLOCK_slh__n424;
wire CLOCK_slh__n430;
wire CLOCK_slh__n431;
wire CLOCK_slh__n432;
wire CLOCK_slh__n438;
wire CLOCK_slh__n439;
wire CLOCK_slh__n440;
wire CLOCK_slh__n446;
wire CLOCK_slh__n447;
wire CLOCK_slh__n448;
wire CLOCK_slh__n452;
wire CLOCK_slh__n453;
wire CLOCK_slh__n454;
wire CLOCK_slh__n458;
wire CLOCK_slh__n459;
wire CLOCK_slh__n460;
wire CLOCK_slh__n464;
wire CLOCK_slh__n465;
wire CLOCK_slh__n466;
wire CLOCK_slh__n470;
wire CLOCK_slh__n471;
wire CLOCK_slh__n472;


NOR2_X1 i_0_1_196 (.ZN (n_0_1_104), .A1 (B_reg), .A2 (A_reg));
AOI211_X1 i_0_1_124 (.ZN (n_0_102), .A (reset), .B (n_0_1_104), .C1 (B_reg), .C2 (A_reg));
CLKBUF_X3 CTS_L3_c_tid0_15 (.Z (CTS_n_tid0_13), .A (CTS_n_tid0_14));
AND4_X1 i_0_1_122 (.ZN (n_0_1_102), .A1 (\EB[5] ), .A2 (\EB[4] ), .A3 (\EB[3] ), .A4 (\EB[0] ));
AND3_X1 i_0_1_121 (.ZN (n_0_1_101), .A1 (\EB[2] ), .A2 (\EB[1] ), .A3 (n_0_1_102));
NAND3_X1 i_0_1_120 (.ZN (n_0_1_100), .A1 (\EB[7] ), .A2 (n_0_1_101), .A3 (\EB[6] ));
AND4_X1 i_0_1_119 (.ZN (n_0_1_99), .A1 (\EA[5] ), .A2 (\EA[4] ), .A3 (\EA[3] ), .A4 (\EA[0] ));
AND3_X1 i_0_1_118 (.ZN (n_0_1_98), .A1 (\EA[2] ), .A2 (\EA[1] ), .A3 (n_0_1_99));
NAND3_X1 i_0_1_117 (.ZN (n_0_1_97), .A1 (\EA[7] ), .A2 (n_0_1_98), .A3 (\EA[6] ));
OR4_X1 i_0_1_116 (.ZN (n_0_1_96), .A1 (\EA[3] ), .A2 (\EA[2] ), .A3 (\EA[1] ), .A4 (\EA[0] ));
OR2_X1 i_0_1_115 (.ZN (n_0_1_95), .A1 (\EA[7] ), .A2 (\EA[6] ));
OR4_X1 i_0_1_114 (.ZN (n_0_1_94), .A1 (n_0_1_96), .A2 (n_0_1_95), .A3 (\EA[5] ), .A4 (\EA[4] ));
OR4_X1 i_0_1_113 (.ZN (n_0_1_93), .A1 (\EB[3] ), .A2 (\EB[2] ), .A3 (\EB[1] ), .A4 (\EB[0] ));
OR2_X1 i_0_1_112 (.ZN (n_0_1_92), .A1 (\EB[7] ), .A2 (\EB[6] ));
OR4_X1 i_0_1_111 (.ZN (n_0_1_91), .A1 (n_0_1_93), .A2 (n_0_1_92), .A3 (\EB[5] ), .A4 (\EB[4] ));
OAI22_X1 i_0_1_110 (.ZN (n_0_1_90), .A1 (n_0_1_100), .A2 (n_0_1_94), .B1 (n_0_1_97), .B2 (n_0_1_91));
INV_X1 i_0_1_109 (.ZN (n_0_1_89), .A (n_0_1_90));
NOR4_X1 i_0_1_108 (.ZN (n_0_1_88), .A1 (n_0_52), .A2 (n_0_53), .A3 (n_0_54), .A4 (n_0_55));
NOR4_X1 i_0_1_107 (.ZN (n_0_1_87), .A1 (n_0_48), .A2 (n_0_49), .A3 (n_0_50), .A4 (n_0_51));
NOR4_X1 i_0_1_106 (.ZN (n_0_1_86), .A1 (n_0_61), .A2 (n_0_62), .A3 (n_0_56), .A4 (n_0_59));
NOR3_X1 i_0_1_105 (.ZN (n_0_1_85), .A1 (n_0_65), .A2 (n_0_66), .A3 (n_0_69));
NOR4_X1 i_0_1_104 (.ZN (n_0_1_84), .A1 (n_0_60), .A2 (n_0_63), .A3 (n_0_57), .A4 (n_0_58));
NOR4_X1 i_0_1_103 (.ZN (n_0_1_83), .A1 (n_0_68), .A2 (n_0_70), .A3 (n_0_64), .A4 (n_0_67));
AND4_X1 i_0_1_102 (.ZN (n_0_1_82), .A1 (n_0_1_88), .A2 (n_0_1_87), .A3 (n_0_1_84), .A4 (n_0_1_83));
NAND3_X1 i_0_1_101 (.ZN (n_0_1_81), .A1 (n_0_1_86), .A2 (n_0_1_85), .A3 (n_0_1_82));
NOR4_X1 i_0_1_100 (.ZN (n_0_1_80), .A1 (n_0_29), .A2 (n_0_30), .A3 (n_0_31), .A4 (n_0_32));
NOR4_X1 i_0_1_99 (.ZN (n_0_1_79), .A1 (n_0_25), .A2 (n_0_26), .A3 (n_0_27), .A4 (n_0_28));
NOR4_X1 i_0_1_98 (.ZN (n_0_1_78), .A1 (n_0_38), .A2 (n_0_39), .A3 (n_0_33), .A4 (n_0_36));
NOR3_X1 i_0_1_97 (.ZN (n_0_1_77), .A1 (n_0_42), .A2 (n_0_43), .A3 (n_0_46));
NOR4_X1 i_0_1_96 (.ZN (n_0_1_76), .A1 (n_0_37), .A2 (n_0_40), .A3 (n_0_34), .A4 (n_0_35));
NOR4_X1 i_0_1_95 (.ZN (n_0_1_75), .A1 (n_0_45), .A2 (n_0_47), .A3 (n_0_41), .A4 (n_0_44));
AND4_X1 i_0_1_94 (.ZN (n_0_1_74), .A1 (n_0_1_80), .A2 (n_0_1_79), .A3 (n_0_1_76), .A4 (n_0_1_75));
NAND3_X1 i_0_1_93 (.ZN (n_0_1_73), .A1 (n_0_1_78), .A2 (n_0_1_77), .A3 (n_0_1_74));
NOR4_X1 i_0_1_92 (.ZN (n_0_1_72), .A1 (reset), .A2 (n_0_1_73), .A3 (n_0_1_81), .A4 (n_0_1_89));
INV_X1 i_0_1_91 (.ZN (n_0_1_71), .A (n_0_1_72));
OAI22_X1 i_0_1_90 (.ZN (n_0_1_70), .A1 (n_0_1_91), .A2 (n_0_1_81), .B1 (n_0_1_94), .B2 (n_0_1_73));
NOR2_X1 i_0_1_89 (.ZN (n_0_1_69), .A1 (reset), .A2 (n_0_1_70));
AND2_X1 i_0_1_88 (.ZN (n_0_1_68), .A1 (\EA[7] ), .A2 (\EB[7] ));
OAI221_X1 i_0_1_87 (.ZN (n_0_1_67), .A (n_0_1_68), .B1 (\EA[6] ), .B2 (n_0_1_98), .C1 (\EB[6] ), .C2 (n_0_1_101));
OR4_X1 i_0_1_86 (.ZN (n_0_1_66), .A1 (n_0_1_101), .A2 (n_0_1_98), .A3 (n_0_1_92), .A4 (n_0_1_95));
AOI22_X1 i_0_1_85 (.ZN (n_0_1_65), .A1 (n_0_1_29), .A2 (n_0_0), .B1 (n_0_24), .B2 (\M_resultTruncated[0] ));
NAND2_X1 i_0_1_84 (.ZN (n_0_1_63), .A1 (n_0_1_67), .A2 (n_0_1_66));
OAI211_X1 i_0_1_83 (.ZN (n_0_1_61), .A (n_0_1_100), .B (n_0_1_97), .C1 (n_0_1_65), .C2 (n_0_1_63));
INV_X1 i_0_1_82 (.ZN (n_0_1_31), .A (n_0_1_61));
OAI221_X1 i_0_1_81 (.ZN (n_0_1_30), .A (n_0_1_69), .B1 (n_0_1_100), .B2 (n_0_1_81)
    , .C1 (n_0_1_97), .C2 (n_0_1_73));
OAI21_X1 i_0_1_80 (.ZN (n_0_71), .A (n_0_1_71), .B1 (n_0_1_31), .B2 (n_0_1_30));
INV_X1 i_0_1_79 (.ZN (n_0_1_29), .A (n_0_24));
INV_X1 i_0_1_198 (.ZN (n_0_1_28), .A (enable));
INV_X1 i_0_1_78 (.ZN (n_0_1_112), .A (reset));
INV_X1 i_0_1_66 (.ZN (n_0_1_111), .A (n_0_1_14));
INV_X1 i_0_1_195 (.ZN (n_0_1_110), .A (n_0_1_22));
INV_X1 i_0_1_194 (.ZN (n_0_1_109), .A (n_0_1_23));
INV_X1 i_0_1_193 (.ZN (n_0_1_108), .A (n_0_1_24));
INV_X1 i_0_1_192 (.ZN (n_0_1_107), .A (n_0_1_25));
INV_X1 i_0_1_191 (.ZN (n_0_1_106), .A (n_0_1_26));
INV_X1 i_0_1_190 (.ZN (n_0_1_105), .A (n_0_1_27));
OR2_X2 i_0_1_189 (.ZN (n_0_168), .A1 (CTS_n_tid0_90), .A2 (reset));
AND2_X1 i_0_1_188 (.ZN (CLOCK_slh__n226), .A1 (hfn_ipo_n11), .A2 (B[30]));
AND2_X1 i_0_1_187 (.ZN (CLOCK_slh__n222), .A1 (hfn_ipo_n11), .A2 (B[29]));
AND2_X1 i_0_1_186 (.ZN (CLOCK_slh__n214), .A1 (hfn_ipo_n11), .A2 (B[28]));
AND2_X1 i_0_1_185 (.ZN (CLOCK_slh__n210), .A1 (hfn_ipo_n11), .A2 (B[27]));
AND2_X1 i_0_1_184 (.ZN (CLOCK_slh__n206), .A1 (hfn_ipo_n11), .A2 (B[26]));
AND2_X1 i_0_1_183 (.ZN (CLOCK_slh__n202), .A1 (hfn_ipo_n11), .A2 (B[25]));
AND2_X1 i_0_1_182 (.ZN (CLOCK_slh__n178), .A1 (hfn_ipo_n11), .A2 (B[24]));
AND2_X1 i_0_1_181 (.ZN (CLOCK_slh__n310), .A1 (hfn_ipo_n11), .A2 (B[23]));
AND2_X1 i_0_1_180 (.ZN (CLOCK_slh__n258), .A1 (hfn_ipo_n11), .A2 (B[22]));
AND2_X1 i_0_1_179 (.ZN (CLOCK_slh__n266), .A1 (hfn_ipo_n11), .A2 (B[21]));
AND2_X1 i_0_1_178 (.ZN (CLOCK_slh__n246), .A1 (hfn_ipo_n11), .A2 (B[20]));
AND2_X1 i_0_1_177 (.ZN (CLOCK_slh__n254), .A1 (hfn_ipo_n11), .A2 (B[19]));
AND2_X1 i_0_1_176 (.ZN (CLOCK_slh__n294), .A1 (hfn_ipo_n10), .A2 (B[18]));
AND2_X1 i_0_1_175 (.ZN (CLOCK_slh__n374), .A1 (hfn_ipo_n10), .A2 (B[17]));
AND2_X1 i_0_1_174 (.ZN (CLOCK_slh__n318), .A1 (hfn_ipo_n10), .A2 (B[16]));
AND2_X1 i_0_1_173 (.ZN (CLOCK_slh__n398), .A1 (hfn_ipo_n10), .A2 (B[15]));
AND2_X1 i_0_1_172 (.ZN (CLOCK_slh__n362), .A1 (hfn_ipo_n10), .A2 (B[14]));
AND2_X1 i_0_1_171 (.ZN (CLOCK_slh__n370), .A1 (hfn_ipo_n10), .A2 (B[13]));
AND2_X1 i_0_1_170 (.ZN (CLOCK_slh__n354), .A1 (hfn_ipo_n10), .A2 (B[12]));
AND2_X1 i_0_1_169 (.ZN (CLOCK_slh__n392), .A1 (hfn_ipo_n10), .A2 (B[11]));
AND2_X1 i_0_1_168 (.ZN (CLOCK_slh__n298), .A1 (hfn_ipo_n10), .A2 (B[10]));
AND2_X1 i_0_1_167 (.ZN (CLOCK_slh__n334), .A1 (hfn_ipo_n10), .A2 (B[9]));
AND2_X1 i_0_1_166 (.ZN (CLOCK_slh__n270), .A1 (hfn_ipo_n10), .A2 (B[8]));
AND2_X1 i_0_1_165 (.ZN (CLOCK_slh__n330), .A1 (hfn_ipo_n10), .A2 (B[7]));
AND2_X1 i_0_1_164 (.ZN (CLOCK_slh__n314), .A1 (hfn_ipo_n10), .A2 (B[6]));
AND2_X1 i_0_1_163 (.ZN (CLOCK_slh__n306), .A1 (hfn_ipo_n10), .A2 (B[5]));
AND2_X1 i_0_1_162 (.ZN (CLOCK_slh__n302), .A1 (hfn_ipo_n10), .A2 (B[4]));
AND2_X1 i_0_1_161 (.ZN (CLOCK_slh__n282), .A1 (hfn_ipo_n10), .A2 (B[3]));
AND2_X1 i_0_1_160 (.ZN (CLOCK_slh__n390), .A1 (hfn_ipo_n10), .A2 (B[2]));
AND2_X1 i_0_1_159 (.ZN (CLOCK_slh__n338), .A1 (hfn_ipo_n10), .A2 (B[1]));
AND2_X1 i_0_1_158 (.ZN (CLOCK_slh__n386), .A1 (hfn_ipo_n10), .A2 (B[0]));
AND2_X1 i_0_1_157 (.ZN (CLOCK_slh__n234), .A1 (hfn_ipo_n11), .A2 (A[30]));
AND2_X1 i_0_1_156 (.ZN (CLOCK_slh__n238), .A1 (hfn_ipo_n11), .A2 (A[29]));
AND2_X1 i_0_1_155 (.ZN (CLOCK_slh__n218), .A1 (hfn_ipo_n11), .A2 (A[28]));
AND2_X1 i_0_1_154 (.ZN (CLOCK_slh__n186), .A1 (hfn_ipo_n11), .A2 (A[27]));
AND2_X1 i_0_1_153 (.ZN (CLOCK_slh__n198), .A1 (hfn_ipo_n11), .A2 (A[26]));
AND2_X1 i_0_1_152 (.ZN (CLOCK_slh__n194), .A1 (hfn_ipo_n11), .A2 (A[25]));
AND2_X1 i_0_1_151 (.ZN (CLOCK_slh__n190), .A1 (hfn_ipo_n11), .A2 (A[24]));
AND2_X1 i_0_1_150 (.ZN (CLOCK_slh__n182), .A1 (hfn_ipo_n11), .A2 (A[23]));
AND2_X1 i_0_1_149 (.ZN (CLOCK_slh__n358), .A1 (hfn_ipo_n11), .A2 (A[22]));
AND2_X1 i_0_1_148 (.ZN (CLOCK_slh__n250), .A1 (hfn_ipo_n11), .A2 (A[21]));
AND2_X1 i_0_1_147 (.ZN (CLOCK_slh__n242), .A1 (hfn_ipo_n11), .A2 (A[20]));
AND2_X1 i_0_1_146 (.ZN (CLOCK_slh__n262), .A1 (hfn_ipo_n11), .A2 (A[19]));
AND2_X1 i_0_1_145 (.ZN (CLOCK_slh__n410), .A1 (hfn_ipo_n10), .A2 (A[18]));
AND2_X1 i_0_1_144 (.ZN (CLOCK_slh__n274), .A1 (hfn_ipo_n11), .A2 (A[17]));
AND2_X1 i_0_1_143 (.ZN (CLOCK_slh__n408), .A1 (hfn_ipo_n10), .A2 (A[16]));
AND2_X1 i_0_1_142 (.ZN (CLOCK_slh__n326), .A1 (hfn_ipo_n10), .A2 (A[15]));
AND2_X1 i_0_1_141 (.ZN (CLOCK_slh__n346), .A1 (hfn_ipo_n11), .A2 (A[14]));
AND2_X1 i_0_1_140 (.ZN (CLOCK_slh__n342), .A1 (hfn_ipo_n11), .A2 (A[13]));
AND2_X1 i_0_1_139 (.ZN (CLOCK_slh__n406), .A1 (hfn_ipo_n10), .A2 (A[12]));
AND2_X1 i_0_1_138 (.ZN (CLOCK_slh__n402), .A1 (hfn_ipo_n10), .A2 (A[11]));
AND2_X1 i_0_1_137 (.ZN (CLOCK_slh__n404), .A1 (hfn_ipo_n11), .A2 (A[10]));
AND2_X1 i_0_1_136 (.ZN (CLOCK_slh__n396), .A1 (hfn_ipo_n10), .A2 (A[9]));
AND2_X1 i_0_1_135 (.ZN (CLOCK_slh__n394), .A1 (hfn_ipo_n11), .A2 (A[8]));
AND2_X1 i_0_1_134 (.ZN (CLOCK_slh__n322), .A1 (hfn_ipo_n10), .A2 (A[7]));
AND2_X1 i_0_1_133 (.ZN (CLOCK_slh__n366), .A1 (hfn_ipo_n10), .A2 (A[6]));
AND2_X1 i_0_1_132 (.ZN (CLOCK_slh__n278), .A1 (hfn_ipo_n10), .A2 (A[5]));
AND2_X1 i_0_1_131 (.ZN (CLOCK_slh__n290), .A1 (hfn_ipo_n10), .A2 (A[4]));
AND2_X1 i_0_1_130 (.ZN (CLOCK_slh__n382), .A1 (hfn_ipo_n10), .A2 (A[3]));
AND2_X1 i_0_1_129 (.ZN (CLOCK_slh__n378), .A1 (hfn_ipo_n10), .A2 (A[2]));
AND2_X1 i_0_1_128 (.ZN (CLOCK_slh__n350), .A1 (hfn_ipo_n10), .A2 (A[1]));
AND2_X1 i_0_1_127 (.ZN (CLOCK_slh__n400), .A1 (hfn_ipo_n10), .A2 (A[0]));
AND2_X1 i_0_1_126 (.ZN (CLOCK_slh__n286), .A1 (hfn_ipo_n11), .A2 (B[31]));
OAI21_X4 i_0_1_125 (.ZN (CTS_n_tid0_14), .A (hfn_ipo_n11), .B1 (n_0_1_28), .B2 (CTS_n_tid0_91));
AND2_X1 i_0_1_65 (.ZN (CLOCK_slh__n230), .A1 (hfn_ipo_n11), .A2 (A[31]));
NAND3_X1 i_0_1_64 (.ZN (n_0_1_64), .A1 (n_0_1_100), .A2 (n_0_1_97), .A3 (n_0_1_67));
AOI21_X1 i_0_1_21 (.ZN (n_0_1_62), .A (n_0_1_72), .B1 (n_0_1_69), .B2 (n_0_1_64));
NAND2_X1 i_0_1_20 (.ZN (n_0_1_60), .A1 (n_0_1_69), .A2 (n_0_1_66));
NOR2_X1 i_0_1_77 (.ZN (n_0_1_59), .A1 (\EB[7] ), .A2 (\EA[7] ));
NOR2_X1 i_0_1_76 (.ZN (n_0_1_58), .A1 (n_0_1_68), .A2 (n_0_1_59));
XNOR2_X1 i_0_1_75 (.ZN (n_0_1_57), .A (n_0_1_13), .B (n_0_1_21));
XNOR2_X1 i_0_1_74 (.ZN (n_0_1_56), .A (n_0_1_58), .B (n_0_1_57));
OAI21_X1 i_0_1_73 (.ZN (n_0_101), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_56));
OAI21_X1 i_0_1_72 (.ZN (n_0_100), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_105));
OAI21_X1 i_0_1_71 (.ZN (n_0_99), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_106));
OAI21_X1 i_0_1_70 (.ZN (n_0_98), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_107));
OAI21_X1 i_0_1_69 (.ZN (n_0_97), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_108));
OAI21_X1 i_0_1_68 (.ZN (n_0_96), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_109));
OAI21_X1 i_0_1_67 (.ZN (n_0_95), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_110));
OAI21_X1 i_0_1_19 (.ZN (n_0_94), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_111));
NOR3_X4 i_0_1_18 (.ZN (n_0_1_55), .A1 (n_0_1_29), .A2 (n_0_1_64), .A3 (n_0_1_60));
NOR3_X4 i_0_1_17 (.ZN (n_0_1_54), .A1 (n_0_1_60), .A2 (n_0_24), .A3 (n_0_1_64));
AOI22_X1 i_0_1_63 (.ZN (n_0_1_53), .A1 (\M_resultTruncated[22] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_22));
INV_X1 i_0_1_62 (.ZN (n_0_93), .A (n_0_1_53));
AOI22_X1 i_0_1_61 (.ZN (n_0_1_52), .A1 (\M_resultTruncated[21] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_21));
INV_X1 i_0_1_60 (.ZN (n_0_92), .A (n_0_1_52));
AOI22_X1 i_0_1_59 (.ZN (n_0_1_51), .A1 (\M_resultTruncated[20] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_20));
INV_X1 i_0_1_58 (.ZN (n_0_91), .A (n_0_1_51));
AOI22_X1 i_0_1_57 (.ZN (n_0_1_50), .A1 (\M_resultTruncated[19] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_19));
INV_X1 i_0_1_56 (.ZN (n_0_90), .A (n_0_1_50));
AOI22_X1 i_0_1_55 (.ZN (n_0_1_49), .A1 (\M_resultTruncated[18] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_18));
INV_X1 i_0_1_54 (.ZN (n_0_89), .A (n_0_1_49));
AOI22_X1 i_0_1_53 (.ZN (n_0_1_48), .A1 (\M_resultTruncated[17] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_17));
INV_X1 i_0_1_52 (.ZN (n_0_88), .A (n_0_1_48));
AOI22_X1 i_0_1_51 (.ZN (n_0_1_47), .A1 (\M_resultTruncated[16] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_16));
INV_X1 i_0_1_50 (.ZN (n_0_87), .A (n_0_1_47));
AOI22_X1 i_0_1_49 (.ZN (n_0_1_46), .A1 (\M_resultTruncated[15] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_15));
INV_X1 i_0_1_48 (.ZN (n_0_86), .A (n_0_1_46));
AOI22_X1 i_0_1_47 (.ZN (n_0_1_45), .A1 (\M_resultTruncated[14] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_14));
INV_X1 i_0_1_46 (.ZN (n_0_85), .A (n_0_1_45));
AOI22_X1 i_0_1_45 (.ZN (n_0_1_44), .A1 (\M_resultTruncated[13] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_13));
INV_X1 i_0_1_44 (.ZN (n_0_84), .A (n_0_1_44));
AOI22_X1 i_0_1_43 (.ZN (n_0_1_43), .A1 (\M_resultTruncated[12] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_12));
INV_X1 i_0_1_42 (.ZN (n_0_83), .A (n_0_1_43));
AOI22_X1 i_0_1_41 (.ZN (n_0_1_42), .A1 (\M_resultTruncated[11] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_11));
INV_X1 i_0_1_40 (.ZN (n_0_82), .A (n_0_1_42));
AOI22_X1 i_0_1_39 (.ZN (n_0_1_41), .A1 (\M_resultTruncated[10] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_10));
INV_X1 i_0_1_38 (.ZN (n_0_81), .A (n_0_1_41));
AOI22_X1 i_0_1_37 (.ZN (n_0_1_40), .A1 (\M_resultTruncated[9] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_9));
INV_X1 i_0_1_36 (.ZN (n_0_80), .A (n_0_1_40));
AOI22_X1 i_0_1_35 (.ZN (n_0_1_39), .A1 (\M_resultTruncated[8] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_8));
INV_X1 i_0_1_34 (.ZN (n_0_79), .A (n_0_1_39));
AOI22_X1 i_0_1_33 (.ZN (n_0_1_38), .A1 (\M_resultTruncated[7] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_7));
INV_X1 i_0_1_32 (.ZN (n_0_78), .A (n_0_1_38));
AOI22_X1 i_0_1_31 (.ZN (n_0_1_37), .A1 (\M_resultTruncated[6] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_6));
INV_X1 i_0_1_30 (.ZN (n_0_77), .A (n_0_1_37));
AOI22_X1 i_0_1_29 (.ZN (n_0_1_36), .A1 (\M_resultTruncated[5] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_5));
INV_X1 i_0_1_28 (.ZN (n_0_76), .A (n_0_1_36));
AOI22_X1 i_0_1_27 (.ZN (n_0_1_35), .A1 (\M_resultTruncated[4] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_4));
INV_X1 i_0_1_26 (.ZN (n_0_75), .A (n_0_1_35));
AOI22_X1 i_0_1_25 (.ZN (n_0_1_34), .A1 (\M_resultTruncated[3] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_3));
INV_X1 i_0_1_24 (.ZN (n_0_74), .A (n_0_1_34));
AOI22_X1 i_0_1_23 (.ZN (n_0_1_33), .A1 (\M_resultTruncated[2] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_2));
INV_X1 i_0_1_22 (.ZN (n_0_73), .A (n_0_1_33));
AOI22_X1 i_0_1_16 (.ZN (n_0_1_32), .A1 (\M_resultTruncated[1] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_1));
INV_X1 i_0_1_15 (.ZN (n_0_72), .A (n_0_1_32));
OR2_X1 i_0_1_14 (.ZN (n_0_1_1), .A1 (\EB[0] ), .A2 (n_0_24));
XNOR2_X1 i_0_1_13 (.ZN (n_0_1_0), .A (\EB[0] ), .B (n_0_24));
FA_X1 i_0_1_12 (.CO (n_0_1_21), .S (n_0_1_27), .A (n_0_1_11), .B (n_0_1_12), .CI (n_0_1_20));
FA_X1 i_0_1_11 (.CO (n_0_1_20), .S (n_0_1_26), .A (n_0_1_9), .B (n_0_1_10), .CI (n_0_1_19));
FA_X1 i_0_1_10 (.CO (n_0_1_19), .S (n_0_1_25), .A (n_0_1_7), .B (n_0_1_8), .CI (n_0_1_18));
FA_X1 i_0_1_9 (.CO (n_0_1_18), .S (n_0_1_24), .A (n_0_1_5), .B (n_0_1_6), .CI (n_0_1_17));
FA_X1 i_0_1_8 (.CO (n_0_1_17), .S (n_0_1_23), .A (n_0_1_3), .B (n_0_1_4), .CI (n_0_1_16));
FA_X1 i_0_1_7 (.CO (n_0_1_16), .S (n_0_1_22), .A (n_0_1_1), .B (n_0_1_2), .CI (n_0_1_15));
HA_X1 i_0_1_6 (.CO (n_0_1_15), .S (n_0_1_14), .A (\EA[0] ), .B (n_0_1_0));
HA_X1 i_0_1_5 (.CO (n_0_1_13), .S (n_0_1_12), .A (\EB[6] ), .B (\EA[6] ));
HA_X1 i_0_1_4 (.CO (n_0_1_11), .S (n_0_1_10), .A (\EB[5] ), .B (\EA[5] ));
HA_X1 i_0_1_3 (.CO (n_0_1_9), .S (n_0_1_8), .A (\EB[4] ), .B (\EA[4] ));
HA_X1 i_0_1_2 (.CO (n_0_1_7), .S (n_0_1_6), .A (\EB[3] ), .B (\EA[3] ));
HA_X1 i_0_1_1 (.CO (n_0_1_5), .S (n_0_1_4), .A (\EB[2] ), .B (\EA[2] ));
HA_X1 i_0_1_0 (.CO (n_0_1_3), .S (n_0_1_2), .A (\EB[1] ), .B (\EA[1] ));
DLH_X1 \B_reg_reg[31]  (.Q (B_reg), .D (n_0_105), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[31]  (.Q (A_reg), .D (n_0_103), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[0]  (.Q (n_0_70), .D (n_0_137), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[1]  (.Q (n_0_69), .D (n_0_138), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[2]  (.Q (n_0_68), .D (n_0_139), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[3]  (.Q (n_0_67), .D (n_0_140), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[4]  (.Q (n_0_66), .D (n_0_141), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[5]  (.Q (n_0_65), .D (n_0_142), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[6]  (.Q (n_0_64), .D (n_0_143), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[7]  (.Q (n_0_63), .D (n_0_144), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[8]  (.Q (n_0_62), .D (n_0_145), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[9]  (.Q (n_0_61), .D (n_0_146), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[10]  (.Q (n_0_60), .D (n_0_147), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[11]  (.Q (n_0_59), .D (n_0_148), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[12]  (.Q (n_0_58), .D (n_0_149), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[13]  (.Q (n_0_57), .D (n_0_150), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[14]  (.Q (n_0_56), .D (n_0_151), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[15]  (.Q (n_0_55), .D (n_0_152), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[16]  (.Q (n_0_54), .D (n_0_153), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[17]  (.Q (n_0_53), .D (n_0_154), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[18]  (.Q (n_0_52), .D (n_0_155), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[19]  (.Q (n_0_51), .D (n_0_156), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[20]  (.Q (n_0_50), .D (n_0_157), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[21]  (.Q (n_0_49), .D (n_0_158), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[22]  (.Q (n_0_48), .D (n_0_159), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[23]  (.Q (\EB[0] ), .D (n_0_160), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[24]  (.Q (\EB[1] ), .D (n_0_161), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[25]  (.Q (\EB[2] ), .D (n_0_162), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[26]  (.Q (\EB[3] ), .D (n_0_163), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[27]  (.Q (\EB[4] ), .D (n_0_164), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[28]  (.Q (\EB[5] ), .D (n_0_165), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[29]  (.Q (\EB[6] ), .D (n_0_166), .G (CTS_n_tid0_13));
DLH_X1 \B_reg_reg[30]  (.Q (\EB[7] ), .D (n_0_167), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[0]  (.Q (n_0_47), .D (n_0_106), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[1]  (.Q (n_0_46), .D (n_0_107), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[2]  (.Q (n_0_45), .D (n_0_108), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[3]  (.Q (n_0_44), .D (n_0_109), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[4]  (.Q (n_0_43), .D (n_0_110), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[5]  (.Q (n_0_42), .D (n_0_111), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[6]  (.Q (n_0_41), .D (n_0_112), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[7]  (.Q (n_0_40), .D (n_0_113), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[8]  (.Q (n_0_39), .D (n_0_114), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[9]  (.Q (n_0_38), .D (n_0_115), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[10]  (.Q (n_0_37), .D (n_0_116), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[11]  (.Q (n_0_36), .D (n_0_117), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[12]  (.Q (n_0_35), .D (n_0_118), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[13]  (.Q (n_0_34), .D (n_0_119), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[14]  (.Q (n_0_33), .D (n_0_120), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[15]  (.Q (n_0_32), .D (n_0_121), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[16]  (.Q (n_0_31), .D (n_0_122), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[17]  (.Q (n_0_30), .D (n_0_123), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[18]  (.Q (n_0_29), .D (n_0_124), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[19]  (.Q (n_0_28), .D (n_0_125), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[20]  (.Q (n_0_27), .D (n_0_126), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[21]  (.Q (n_0_26), .D (n_0_127), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[22]  (.Q (n_0_25), .D (n_0_128), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[23]  (.Q (\EA[0] ), .D (n_0_129), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[24]  (.Q (\EA[1] ), .D (n_0_130), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[25]  (.Q (\EA[2] ), .D (n_0_131), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[26]  (.Q (\EA[3] ), .D (n_0_132), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[27]  (.Q (\EA[4] ), .D (n_0_133), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[28]  (.Q (\EA[5] ), .D (n_0_134), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[29]  (.Q (\EA[6] ), .D (n_0_135), .G (CTS_n_tid0_13));
DLH_X1 \A_reg_reg[30]  (.Q (\EA[7] ), .D (n_0_136), .G (CTS_n_tid0_13));
DLH_X1 \Res_reg[0]  (.Q (Res[0]), .D (n_0_71), .G (n_0_168));
DLH_X1 \Res_reg[1]  (.Q (Res[1]), .D (n_0_72), .G (n_0_168));
DLH_X1 \Res_reg[2]  (.Q (Res[2]), .D (n_0_73), .G (n_0_168));
DLH_X1 \Res_reg[3]  (.Q (Res[3]), .D (n_0_74), .G (n_0_168));
DLH_X1 \Res_reg[4]  (.Q (Res[4]), .D (n_0_75), .G (n_0_168));
DLH_X1 \Res_reg[5]  (.Q (Res[5]), .D (n_0_76), .G (n_0_168));
DLH_X1 \Res_reg[6]  (.Q (Res[6]), .D (n_0_77), .G (n_0_168));
DLH_X1 \Res_reg[7]  (.Q (Res[7]), .D (n_0_78), .G (n_0_168));
DLH_X1 \Res_reg[8]  (.Q (Res[8]), .D (n_0_79), .G (n_0_168));
DLH_X1 \Res_reg[9]  (.Q (Res[9]), .D (n_0_80), .G (n_0_168));
DLH_X1 \Res_reg[10]  (.Q (Res[10]), .D (n_0_81), .G (n_0_168));
DLH_X1 \Res_reg[11]  (.Q (Res[11]), .D (n_0_82), .G (n_0_168));
DLH_X1 \Res_reg[12]  (.Q (Res[12]), .D (n_0_83), .G (n_0_168));
DLH_X1 \Res_reg[13]  (.Q (Res[13]), .D (n_0_84), .G (n_0_168));
DLH_X1 \Res_reg[14]  (.Q (Res[14]), .D (n_0_85), .G (n_0_168));
DLH_X1 \Res_reg[15]  (.Q (Res[15]), .D (n_0_86), .G (n_0_168));
DLH_X1 \Res_reg[16]  (.Q (Res[16]), .D (n_0_87), .G (n_0_168));
DLH_X1 \Res_reg[17]  (.Q (Res[17]), .D (n_0_88), .G (n_0_168));
DLH_X1 \Res_reg[18]  (.Q (Res[18]), .D (n_0_89), .G (n_0_168));
DLH_X1 \Res_reg[19]  (.Q (Res[19]), .D (n_0_90), .G (n_0_168));
DLH_X1 \Res_reg[20]  (.Q (Res[20]), .D (n_0_91), .G (n_0_168));
DLH_X1 \Res_reg[21]  (.Q (Res[21]), .D (n_0_92), .G (n_0_168));
DLH_X1 \Res_reg[22]  (.Q (Res[22]), .D (n_0_93), .G (n_0_168));
DLH_X1 \Res_reg[23]  (.Q (Res[23]), .D (n_0_94), .G (n_0_168));
DLH_X1 \Res_reg[24]  (.Q (Res[24]), .D (n_0_95), .G (n_0_168));
DLH_X1 \Res_reg[25]  (.Q (Res[25]), .D (n_0_96), .G (n_0_168));
DLH_X1 \Res_reg[26]  (.Q (Res[26]), .D (n_0_97), .G (n_0_168));
DLH_X1 \Res_reg[27]  (.Q (Res[27]), .D (n_0_98), .G (n_0_168));
DLH_X1 \Res_reg[28]  (.Q (Res[28]), .D (n_0_99), .G (n_0_168));
DLH_X1 \Res_reg[29]  (.Q (Res[29]), .D (n_0_100), .G (n_0_168));
DLH_X1 \Res_reg[30]  (.Q (Res[30]), .D (n_0_101), .G (n_0_168));
DLH_X1 \Res_reg[31]  (.Q (Res[31]), .D (n_0_102), .G (n_0_168));
datapath__0_13 i_0_0 (.M_resultTruncated ({\M_resultTruncated[22] , \M_resultTruncated[21] , 
    \M_resultTruncated[20] , \M_resultTruncated[19] , \M_resultTruncated[18] , \M_resultTruncated[17] , 
    \M_resultTruncated[16] , \M_resultTruncated[15] , \M_resultTruncated[14] , \M_resultTruncated[13] , 
    \M_resultTruncated[12] , \M_resultTruncated[11] , \M_resultTruncated[10] , \M_resultTruncated[9] , 
    \M_resultTruncated[8] , \M_resultTruncated[7] , \M_resultTruncated[6] , \M_resultTruncated[5] , 
    \M_resultTruncated[4] , \M_resultTruncated[3] , \M_resultTruncated[2] , \M_resultTruncated[1] , 
    \M_resultTruncated[0] }), .M_multiplied (n_0_0), .p_0 ({n_0_23, n_0_22, n_0_21, 
    n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, 
    n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1}));
VM multiplier (.Res ({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, uc_9, 
    uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, 
    n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, 
    n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, uc_16, 
    uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, 
    uc_28, uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, uc_38})
    , .clk_CTS_0_PP_4 (CTS_n_tid0_90), .clk_CTS_0_PP_5 (CTS_n_tid0_91), .A ({uc_39, 
    uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, n_0_25, n_0_26, n_0_27, 
    n_0_28, n_0_29, n_0_30, n_0_31, n_0_32, n_0_33, n_0_34, n_0_35, n_0_36, n_0_37, 
    n_0_38, n_0_39, n_0_40, n_0_41, n_0_42, n_0_43, n_0_44, n_0_45, n_0_46, n_0_47})
    , .B ({uc_48, uc_49, uc_50, uc_51, uc_52, uc_53, uc_54, uc_55, uc_56, n_0_48, 
    n_0_49, n_0_50, n_0_51, n_0_52, n_0_53, n_0_54, n_0_55, n_0_56, n_0_57, n_0_58, 
    n_0_59, n_0_60, n_0_61, n_0_62, n_0_63, n_0_64, n_0_65, n_0_66, n_0_67, n_0_68, 
    n_0_69, n_0_70}), .enable (CLOCK_slh__n413), .reset (reset), .clk_CTS_0_PP_6 (clk));
CLKBUF_X3 hfn_ipo_c10 (.Z (hfn_ipo_n10), .A (n_0_1_112));
CLKBUF_X1 hfn_ipo_c11 (.Z (hfn_ipo_n11), .A (n_0_1_112));
CLKBUF_X1 CLOCK_slh__c78 (.Z (n_0_161), .A (CLOCK_slh__n179));
CLKBUF_X1 CLOCK_slh__c77 (.Z (CLOCK_slh__n179), .A (CLOCK_slh__n178));
CLKBUF_X1 CLOCK_slh__c81 (.Z (CLOCK_slh__n183), .A (CLOCK_slh__n182));
CLKBUF_X1 CLOCK_slh__c82 (.Z (n_0_129), .A (CLOCK_slh__n183));
CLKBUF_X1 CLOCK_slh__c85 (.Z (CLOCK_slh__n187), .A (CLOCK_slh__n186));
CLKBUF_X1 CLOCK_slh__c86 (.Z (n_0_133), .A (CLOCK_slh__n187));
CLKBUF_X1 CLOCK_slh__c89 (.Z (CLOCK_slh__n191), .A (CLOCK_slh__n190));
CLKBUF_X1 CLOCK_slh__c90 (.Z (n_0_130), .A (CLOCK_slh__n191));
CLKBUF_X1 CLOCK_slh__c93 (.Z (CLOCK_slh__n195), .A (CLOCK_slh__n194));
CLKBUF_X1 CLOCK_slh__c94 (.Z (n_0_131), .A (CLOCK_slh__n195));
CLKBUF_X1 CLOCK_slh__c97 (.Z (CLOCK_slh__n199), .A (CLOCK_slh__n198));
CLKBUF_X1 CLOCK_slh__c98 (.Z (n_0_132), .A (CLOCK_slh__n199));
CLKBUF_X1 CLOCK_slh__c101 (.Z (CLOCK_slh__n203), .A (CLOCK_slh__n202));
CLKBUF_X1 CLOCK_slh__c102 (.Z (n_0_162), .A (CLOCK_slh__n203));
CLKBUF_X1 CLOCK_slh__c105 (.Z (CLOCK_slh__n207), .A (CLOCK_slh__n206));
CLKBUF_X1 CLOCK_slh__c106 (.Z (n_0_163), .A (CLOCK_slh__n207));
CLKBUF_X1 CLOCK_slh__c109 (.Z (CLOCK_slh__n211), .A (CLOCK_slh__n210));
CLKBUF_X1 CLOCK_slh__c110 (.Z (n_0_164), .A (CLOCK_slh__n211));
CLKBUF_X1 CLOCK_slh__c113 (.Z (CLOCK_slh__n215), .A (CLOCK_slh__n214));
CLKBUF_X1 CLOCK_slh__c114 (.Z (n_0_165), .A (CLOCK_slh__n215));
CLKBUF_X1 CLOCK_slh__c117 (.Z (CLOCK_slh__n219), .A (CLOCK_slh__n218));
CLKBUF_X1 CLOCK_slh__c118 (.Z (n_0_134), .A (CLOCK_slh__n219));
CLKBUF_X1 CLOCK_slh__c121 (.Z (CLOCK_slh__n223), .A (CLOCK_slh__n222));
CLKBUF_X1 CLOCK_slh__c122 (.Z (n_0_166), .A (CLOCK_slh__n223));
CLKBUF_X1 CLOCK_slh__c125 (.Z (CLOCK_slh__n227), .A (CLOCK_slh__n226));
CLKBUF_X1 CLOCK_slh__c126 (.Z (n_0_167), .A (CLOCK_slh__n227));
CLKBUF_X1 CLOCK_slh__c129 (.Z (CLOCK_slh__n231), .A (CLOCK_slh__n230));
CLKBUF_X1 CLOCK_slh__c130 (.Z (n_0_103), .A (CLOCK_slh__n231));
CLKBUF_X1 CLOCK_slh__c133 (.Z (CLOCK_slh__n235), .A (CLOCK_slh__n234));
CLKBUF_X1 CLOCK_slh__c134 (.Z (n_0_136), .A (CLOCK_slh__n235));
CLKBUF_X1 CLOCK_slh__c137 (.Z (CLOCK_slh__n239), .A (CLOCK_slh__n238));
CLKBUF_X1 CLOCK_slh__c138 (.Z (n_0_135), .A (CLOCK_slh__n239));
CLKBUF_X1 CLOCK_slh__c141 (.Z (CLOCK_slh__n243), .A (CLOCK_slh__n242));
CLKBUF_X1 CLOCK_slh__c142 (.Z (n_0_126), .A (CLOCK_slh__n243));
CLKBUF_X1 CLOCK_slh__c145 (.Z (CLOCK_slh__n247), .A (CLOCK_slh__n246));
CLKBUF_X1 CLOCK_slh__c146 (.Z (n_0_157), .A (CLOCK_slh__n247));
CLKBUF_X1 CLOCK_slh__c149 (.Z (CLOCK_slh__n251), .A (CLOCK_slh__n250));
CLKBUF_X1 CLOCK_slh__c150 (.Z (n_0_127), .A (CLOCK_slh__n251));
CLKBUF_X1 CLOCK_slh__c153 (.Z (CLOCK_slh__n255), .A (CLOCK_slh__n254));
CLKBUF_X1 CLOCK_slh__c154 (.Z (n_0_156), .A (CLOCK_slh__n255));
CLKBUF_X1 CLOCK_slh__c157 (.Z (CLOCK_slh__n259), .A (CLOCK_slh__n258));
CLKBUF_X1 CLOCK_slh__c158 (.Z (n_0_159), .A (CLOCK_slh__n259));
CLKBUF_X1 CLOCK_slh__c161 (.Z (CLOCK_slh__n263), .A (CLOCK_slh__n262));
CLKBUF_X1 CLOCK_slh__c162 (.Z (n_0_125), .A (CLOCK_slh__n263));
CLKBUF_X1 CLOCK_slh__c165 (.Z (CLOCK_slh__n267), .A (CLOCK_slh__n266));
CLKBUF_X1 CLOCK_slh__c166 (.Z (n_0_158), .A (CLOCK_slh__n267));
CLKBUF_X1 CLOCK_slh__c169 (.Z (CLOCK_slh__n271), .A (CLOCK_slh__n270));
CLKBUF_X1 CLOCK_slh__c170 (.Z (n_0_145), .A (CLOCK_slh__n271));
CLKBUF_X1 CLOCK_slh__c173 (.Z (CLOCK_slh__n275), .A (CLOCK_slh__n274));
CLKBUF_X1 CLOCK_slh__c174 (.Z (n_0_123), .A (CLOCK_slh__n275));
CLKBUF_X1 CLOCK_slh__c177 (.Z (CLOCK_slh__n279), .A (CLOCK_slh__n278));
CLKBUF_X1 CLOCK_slh__c178 (.Z (n_0_111), .A (CLOCK_slh__n279));
CLKBUF_X1 CLOCK_slh__c181 (.Z (CLOCK_slh__n283), .A (CLOCK_slh__n282));
CLKBUF_X1 CLOCK_slh__c182 (.Z (n_0_140), .A (CLOCK_slh__n283));
CLKBUF_X1 CLOCK_slh__c185 (.Z (CLOCK_slh__n287), .A (CLOCK_slh__n286));
CLKBUF_X1 CLOCK_slh__c186 (.Z (n_0_105), .A (CLOCK_slh__n287));
CLKBUF_X1 CLOCK_slh__c189 (.Z (CLOCK_slh__n291), .A (CLOCK_slh__n290));
CLKBUF_X1 CLOCK_slh__c190 (.Z (n_0_110), .A (CLOCK_slh__n291));
CLKBUF_X1 CLOCK_slh__c193 (.Z (CLOCK_slh__n295), .A (CLOCK_slh__n294));
CLKBUF_X1 CLOCK_slh__c194 (.Z (n_0_155), .A (CLOCK_slh__n295));
CLKBUF_X1 CLOCK_slh__c197 (.Z (CLOCK_slh__n299), .A (CLOCK_slh__n298));
CLKBUF_X1 CLOCK_slh__c198 (.Z (n_0_147), .A (CLOCK_slh__n299));
CLKBUF_X1 CLOCK_slh__c201 (.Z (CLOCK_slh__n303), .A (CLOCK_slh__n302));
CLKBUF_X1 CLOCK_slh__c202 (.Z (n_0_141), .A (CLOCK_slh__n303));
CLKBUF_X1 CLOCK_slh__c205 (.Z (CLOCK_slh__n307), .A (CLOCK_slh__n306));
CLKBUF_X1 CLOCK_slh__c206 (.Z (n_0_142), .A (CLOCK_slh__n307));
CLKBUF_X1 CLOCK_slh__c209 (.Z (CLOCK_slh__n311), .A (CLOCK_slh__n310));
CLKBUF_X1 CLOCK_slh__c210 (.Z (n_0_160), .A (CLOCK_slh__n311));
CLKBUF_X1 CLOCK_slh__c213 (.Z (CLOCK_slh__n315), .A (CLOCK_slh__n314));
CLKBUF_X1 CLOCK_slh__c214 (.Z (n_0_143), .A (CLOCK_slh__n315));
CLKBUF_X1 CLOCK_slh__c217 (.Z (CLOCK_slh__n319), .A (CLOCK_slh__n318));
CLKBUF_X1 CLOCK_slh__c218 (.Z (n_0_153), .A (CLOCK_slh__n319));
CLKBUF_X1 CLOCK_slh__c221 (.Z (CLOCK_slh__n323), .A (CLOCK_slh__n322));
CLKBUF_X1 CLOCK_slh__c222 (.Z (n_0_113), .A (CLOCK_slh__n323));
CLKBUF_X1 CLOCK_slh__c225 (.Z (CLOCK_slh__n327), .A (CLOCK_slh__n326));
CLKBUF_X1 CLOCK_slh__c226 (.Z (n_0_121), .A (CLOCK_slh__n327));
CLKBUF_X1 CLOCK_slh__c229 (.Z (CLOCK_slh__n331), .A (CLOCK_slh__n330));
CLKBUF_X1 CLOCK_slh__c230 (.Z (n_0_144), .A (CLOCK_slh__n331));
CLKBUF_X1 CLOCK_slh__c233 (.Z (CLOCK_slh__n335), .A (CLOCK_slh__n334));
CLKBUF_X1 CLOCK_slh__c234 (.Z (n_0_146), .A (CLOCK_slh__n335));
CLKBUF_X1 CLOCK_slh__c237 (.Z (CLOCK_slh__n339), .A (CLOCK_slh__n338));
CLKBUF_X1 CLOCK_slh__c238 (.Z (n_0_138), .A (CLOCK_slh__n339));
CLKBUF_X1 CLOCK_slh__c241 (.Z (CLOCK_slh__n343), .A (CLOCK_slh__n342));
CLKBUF_X1 CLOCK_slh__c242 (.Z (n_0_119), .A (CLOCK_slh__n343));
CLKBUF_X1 CLOCK_slh__c245 (.Z (CLOCK_slh__n347), .A (CLOCK_slh__n346));
CLKBUF_X1 CLOCK_slh__c246 (.Z (n_0_120), .A (CLOCK_slh__n347));
CLKBUF_X1 CLOCK_slh__c249 (.Z (CLOCK_slh__n351), .A (CLOCK_slh__n350));
CLKBUF_X1 CLOCK_slh__c250 (.Z (n_0_107), .A (CLOCK_slh__n351));
CLKBUF_X1 CLOCK_slh__c253 (.Z (CLOCK_slh__n355), .A (CLOCK_slh__n354));
CLKBUF_X1 CLOCK_slh__c254 (.Z (n_0_149), .A (CLOCK_slh__n355));
CLKBUF_X1 CLOCK_slh__c257 (.Z (CLOCK_slh__n359), .A (CLOCK_slh__n358));
CLKBUF_X1 CLOCK_slh__c258 (.Z (n_0_128), .A (CLOCK_slh__n359));
CLKBUF_X1 CLOCK_slh__c261 (.Z (CLOCK_slh__n363), .A (CLOCK_slh__n362));
CLKBUF_X1 CLOCK_slh__c262 (.Z (n_0_151), .A (CLOCK_slh__n363));
CLKBUF_X1 CLOCK_slh__c265 (.Z (CLOCK_slh__n367), .A (CLOCK_slh__n366));
CLKBUF_X1 CLOCK_slh__c266 (.Z (n_0_112), .A (CLOCK_slh__n367));
CLKBUF_X1 CLOCK_slh__c269 (.Z (CLOCK_slh__n371), .A (CLOCK_slh__n370));
CLKBUF_X1 CLOCK_slh__c270 (.Z (n_0_150), .A (CLOCK_slh__n371));
CLKBUF_X1 CLOCK_slh__c273 (.Z (CLOCK_slh__n375), .A (CLOCK_slh__n374));
CLKBUF_X1 CLOCK_slh__c274 (.Z (n_0_154), .A (CLOCK_slh__n375));
CLKBUF_X1 CLOCK_slh__c277 (.Z (CLOCK_slh__n379), .A (CLOCK_slh__n378));
CLKBUF_X1 CLOCK_slh__c278 (.Z (n_0_108), .A (CLOCK_slh__n379));
CLKBUF_X1 CLOCK_slh__c281 (.Z (CLOCK_slh__n383), .A (CLOCK_slh__n382));
CLKBUF_X1 CLOCK_slh__c282 (.Z (n_0_109), .A (CLOCK_slh__n383));
CLKBUF_X1 CLOCK_slh__c285 (.Z (CLOCK_slh__n387), .A (CLOCK_slh__n386));
CLKBUF_X1 CLOCK_slh__c286 (.Z (n_0_137), .A (CLOCK_slh__n387));
CLKBUF_X1 CLOCK_slh__c289 (.Z (CLOCK_slh__n391), .A (CLOCK_slh__n390));
CLKBUF_X1 CLOCK_slh__c290 (.Z (n_0_139), .A (CLOCK_slh__n391));
CLKBUF_X1 CLOCK_slh__c291 (.Z (CLOCK_slh__n393), .A (CLOCK_slh__n392));
CLKBUF_X1 CLOCK_slh__c292 (.Z (n_0_148), .A (CLOCK_slh__n393));
CLKBUF_X1 CLOCK_slh__c293 (.Z (CLOCK_slh__n395), .A (CLOCK_slh__n394));
CLKBUF_X1 CLOCK_slh__c294 (.Z (n_0_114), .A (CLOCK_slh__n395));
CLKBUF_X1 CLOCK_slh__c295 (.Z (CLOCK_slh__n397), .A (CLOCK_slh__n396));
CLKBUF_X1 CLOCK_slh__c296 (.Z (n_0_115), .A (CLOCK_slh__n397));
CLKBUF_X1 CLOCK_slh__c297 (.Z (CLOCK_slh__n399), .A (CLOCK_slh__n398));
CLKBUF_X1 CLOCK_slh__c298 (.Z (n_0_152), .A (CLOCK_slh__n399));
CLKBUF_X1 CLOCK_slh__c299 (.Z (CLOCK_slh__n401), .A (CLOCK_slh__n400));
CLKBUF_X1 CLOCK_slh__c300 (.Z (n_0_106), .A (CLOCK_slh__n401));
CLKBUF_X1 CLOCK_slh__c301 (.Z (CLOCK_slh__n403), .A (CLOCK_slh__n402));
CLKBUF_X1 CLOCK_slh__c302 (.Z (n_0_117), .A (CLOCK_slh__n403));
CLKBUF_X1 CLOCK_slh__c303 (.Z (CLOCK_slh__n405), .A (CLOCK_slh__n404));
CLKBUF_X1 CLOCK_slh__c304 (.Z (n_0_116), .A (CLOCK_slh__n405));
CLKBUF_X1 CLOCK_slh__c305 (.Z (CLOCK_slh__n407), .A (CLOCK_slh__n406));
CLKBUF_X1 CLOCK_slh__c306 (.Z (n_0_118), .A (CLOCK_slh__n407));
CLKBUF_X1 CLOCK_slh__c307 (.Z (CLOCK_slh__n409), .A (CLOCK_slh__n408));
CLKBUF_X1 CLOCK_slh__c308 (.Z (n_0_122), .A (CLOCK_slh__n409));
CLKBUF_X1 CLOCK_slh__c309 (.Z (CLOCK_slh__n411), .A (CLOCK_slh__n410));
CLKBUF_X1 CLOCK_slh__c310 (.Z (n_0_124), .A (CLOCK_slh__n411));
CLKBUF_X1 CLOCK_slh__c311 (.Z (CLOCK_slh__n414), .A (enable));
CLKBUF_X1 CLOCK_slh__c312 (.Z (CLOCK_slh__n415), .A (CLOCK_slh__n414));
CLKBUF_X1 CLOCK_slh__c313 (.Z (CLOCK_slh__n416), .A (CLOCK_slh__n415));
CLKBUF_X1 CLOCK_slh__c314 (.Z (CLOCK_slh__n422), .A (CLOCK_slh__n416));
CLKBUF_X1 CLOCK_slh__c320 (.Z (CLOCK_slh__n423), .A (CLOCK_slh__n422));
CLKBUF_X1 CLOCK_slh__c321 (.Z (CLOCK_slh__n424), .A (CLOCK_slh__n423));
CLKBUF_X1 CLOCK_slh__c322 (.Z (CLOCK_slh__n430), .A (CLOCK_slh__n424));
CLKBUF_X1 CLOCK_slh__c328 (.Z (CLOCK_slh__n431), .A (CLOCK_slh__n430));
CLKBUF_X1 CLOCK_slh__c329 (.Z (CLOCK_slh__n432), .A (CLOCK_slh__n431));
CLKBUF_X1 CLOCK_slh__c330 (.Z (CLOCK_slh__n438), .A (CLOCK_slh__n432));
CLKBUF_X1 CLOCK_slh__c336 (.Z (CLOCK_slh__n439), .A (CLOCK_slh__n438));
CLKBUF_X1 CLOCK_slh__c337 (.Z (CLOCK_slh__n440), .A (CLOCK_slh__n439));
CLKBUF_X1 CLOCK_slh__c338 (.Z (CLOCK_slh__n446), .A (CLOCK_slh__n440));
CLKBUF_X1 CLOCK_slh__c344 (.Z (CLOCK_slh__n447), .A (CLOCK_slh__n446));
CLKBUF_X1 CLOCK_slh__c345 (.Z (CLOCK_slh__n448), .A (CLOCK_slh__n447));
CLKBUF_X1 CLOCK_slh__c346 (.Z (CLOCK_slh__n452), .A (CLOCK_slh__n448));
CLKBUF_X1 CLOCK_slh__c350 (.Z (CLOCK_slh__n453), .A (CLOCK_slh__n452));
CLKBUF_X1 CLOCK_slh__c351 (.Z (CLOCK_slh__n454), .A (CLOCK_slh__n453));
CLKBUF_X1 CLOCK_slh__c352 (.Z (CLOCK_slh__n458), .A (CLOCK_slh__n454));
CLKBUF_X1 CLOCK_slh__c356 (.Z (CLOCK_slh__n459), .A (CLOCK_slh__n458));
CLKBUF_X1 CLOCK_slh__c357 (.Z (CLOCK_slh__n460), .A (CLOCK_slh__n459));
CLKBUF_X1 CLOCK_slh__c358 (.Z (CLOCK_slh__n464), .A (CLOCK_slh__n460));
CLKBUF_X1 CLOCK_slh__c362 (.Z (CLOCK_slh__n465), .A (CLOCK_slh__n464));
CLKBUF_X1 CLOCK_slh__c363 (.Z (CLOCK_slh__n466), .A (CLOCK_slh__n465));
CLKBUF_X1 CLOCK_slh__c364 (.Z (CLOCK_slh__n470), .A (CLOCK_slh__n466));
CLKBUF_X1 CLOCK_slh__c368 (.Z (CLOCK_slh__n471), .A (CLOCK_slh__n470));
CLKBUF_X1 CLOCK_slh__c369 (.Z (CLOCK_slh__n472), .A (CLOCK_slh__n471));
CLKBUF_X1 CLOCK_slh__c370 (.Z (CLOCK_slh__n413), .A (CLOCK_slh__n472));

endmodule //FPU_VM


