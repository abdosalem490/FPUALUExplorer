* SPICE NETLIST
***************************************

.SUBCKT MGC_via1_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via1_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X2
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT WELLTAP
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_3
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUF_X1 A VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
M0 VSS A 5 VSS NMOS_VTL L=5e-08 W=9.5e-08 AD=2.03e-14 AS=9.975e-15 PD=6.7e-07 PS=4e-07 $X=165 $Y=160 $D=1
M1 Z 5 VSS VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.03e-14 PD=6e-07 PS=6.7e-07 $X=355 $Y=160 $D=1
M2 VDD A 5 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=165 $Y=995 $D=0
M3 Z 5 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=355 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=2 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT AND2_X1 A1 A2 VSS VDD ZN
** N=7 EP=5 IP=0 FDC=6
M0 7 A1 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 6 A1 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV_X2 A ZN VSS VDD
** N=4 EP=4 IP=0 FDC=4
M0 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X4
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_12
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7
** N=7 EP=7 IP=9 FDC=10
X0 1 2 3 4 CLKBUF_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 5 6 2 3 7 AND2_X1 $T=-760 0 0 0 $X=-875 $Y=-115
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT via1_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DLH_X1 G Q D VSS VDD
** N=13 EP=5 IP=0 FDC=16
M0 VSS G 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07 $X=170 $Y=90 $D=1
M1 Q 8 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS 6 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=755 $Y=215 $D=1
M3 12 D VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=945 $Y=215 $D=1
M4 8 7 12 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1135 $Y=215 $D=1
M5 13 6 8 VSS NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07 $X=1325 $Y=335 $D=1
M6 VSS 9 13 VSS NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=1515 $Y=335 $D=1
M7 9 8 VSS VSS NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14 PD=3.9e-07 PS=4.6e-07 $X=1705 $Y=335 $D=1
M8 VDD G 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=170 $Y=995 $D=0
M9 Q 8 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M10 VDD 6 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=755 $Y=815 $D=0
M11 10 D VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=945 $Y=815 $D=0
M12 8 6 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1135 $Y=815 $D=0
M13 11 7 8 VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07 $X=1325 $Y=1040 $D=0
M14 VDD 9 11 VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=1515 $Y=1040 $D=0
M15 9 8 VDD VDD PMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14 PD=3.9e-07 PS=4.6e-07 $X=1705 $Y=1040 $D=0
.ENDS
***************************************
.SUBCKT FILLCELL_X8
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_20
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT INV_X4 A ZN VSS VDD
** N=4 EP=4 IP=0 FDC=8
M0 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=2 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT NOR2_X1 A2 VDD A1 ZN VSS 6
** N=7 EP=6 IP=0 FDC=4
M0 ZN A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A1 ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 7 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 ZN A1 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_23 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=4
X1 3 2 4 5 1 1 NOR2_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=4
X1 1 2 3 4 5 ICV_23 $T=380 0 0 0 $X=265 $Y=-115
.ENDS
***************************************
.SUBCKT HA_X1 S B A VSS VDD CO
** N=12 EP=6 IP=0 FDC=16
M0 11 B VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 S A 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS 8 S VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.48e-14 AS=5.81e-14 PD=1.12e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 8 B VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.48e-14 PD=7e-07 PS=1.12e-06 $X=760 $Y=90 $D=1
M4 VSS A 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=950 $Y=90 $D=1
M5 12 A 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1320 $Y=90 $D=1
M6 VSS B 12 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=1510 $Y=90 $D=1
M7 CO 9 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1700 $Y=90 $D=1
M8 S B 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M9 7 A S VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M10 VDD 8 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.7725e-14 AS=8.82e-14 PD=1.55e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M11 10 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.7725e-14 PD=9.1e-07 PS=1.55e-06 $X=760 $Y=870 $D=0
M12 8 A 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=950 $Y=870 $D=0
M13 9 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1320 $Y=870 $D=0
M14 VDD B 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=1510 $Y=870 $D=0
M15 CO 9 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1700 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_25
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=16
X1 3 4 5 1 2 DLH_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=16
X1 3 4 5 1 2 DLH_X1 $T=380 0 0 0 $X=265 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_28
** N=2 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT AOI22_X1 B2 B1 VDD A1 ZN A2 VSS
** N=10 EP=7 IP=0 FDC=8
M0 9 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN B1 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 10 A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 VSS A2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 VDD B2 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 8 B1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 ZN A1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 8 A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_29
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_30
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_31
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_32
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_33
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FA_X1 CO CI B A VDD VSS S 8
** N=20 EP=8 IP=0 FDC=28
M0 VSS 9 CO 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 18 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06 $X=360 $Y=215 $D=1
M2 9 A 18 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=550 $Y=215 $D=1
M3 10 CI 9 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07 $X=740 $Y=215 $D=1
M4 VSS A 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07 $X=935 $Y=215 $D=1
M5 10 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1125 $Y=215 $D=1
M6 12 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1465 $Y=90 $D=1
M7 VSS CI 12 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1655 $Y=90 $D=1
M8 12 A VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1845 $Y=90 $D=1
M9 14 9 12 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07 $X=2035 $Y=90 $D=1
M10 19 CI 14 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.15e-14 PD=7e-07 PS=7.2e-07 $X=2235 $Y=90 $D=1
M11 20 B 19 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2425 $Y=90 $D=1
M12 VSS A 20 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=2615 $Y=90 $D=1
M13 S 14 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=2805 $Y=90 $D=1
M14 VDD 9 CO VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M15 15 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.54e-06 $X=360 $Y=870 $D=0
M16 9 A 15 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=550 $Y=870 $D=0
M17 11 CI 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06 PS=9.1e-07 $X=740 $Y=870 $D=0
M18 VDD A 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.53e-14 PD=9.1e-07 PS=1.07e-06 $X=935 $Y=945 $D=0
M19 11 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1125 $Y=945 $D=0
M20 13 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1465 $Y=995 $D=0
M21 VDD CI 13 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1655 $Y=995 $D=0
M22 13 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1845 $Y=995 $D=0
M23 14 9 13 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07 $X=2035 $Y=995 $D=0
M24 16 CI 14 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.725e-14 PD=9.1e-07 PS=9.3e-07 $X=2235 $Y=995 $D=0
M25 17 B 16 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=2425 $Y=995 $D=0
M26 VDD A 17 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2615 $Y=995 $D=0
M27 S 14 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2805 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_34
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT NOR4_X1 A4 VDD A3 A2 A1 ZN VSS
** N=10 EP=7 IP=0 FDC=8
M0 ZN A4 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A3 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 8 A4 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 9 A3 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 10 A2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 ZN A1 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI21_X1 B2 B1 ZN A VSS VDD
** N=8 EP=6 IP=0 FDC=6
M0 8 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN B1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M4 7 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M5 VDD A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI21_X1 B2 B1 ZN A VSS VDD
** N=8 EP=6 IP=0 FDC=6
M0 ZN B2 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 7 B1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS A 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=550 $Y=90 $D=1
M3 8 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M4 ZN B1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M5 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=550 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_35 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=28
X1 3 4 5 6 2 1 7 1 FA_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_36
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_37
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT INV_X1 A VSS VDD ZN
** N=4 EP=4 IP=0 FDC=2
M0 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI221_X1 B2 B1 VSS A C2 VDD C1 ZN
** N=12 EP=8 IP=0 FDC=10
M0 VSS B2 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 9 B1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 10 A 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN C2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 10 C1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 11 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 ZN B1 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 12 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 ZN C1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI211_X1 C2 C1 B VSS A ZN VDD
** N=10 EP=7 IP=0 FDC=8
M0 10 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN C1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS B ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 ZN C2 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 8 C1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 9 B 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 VDD A 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_38
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_39
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_40
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X16
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_41
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_42
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_43
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_44
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_45
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_46
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_47 1 2 3 4 5 6
** N=6 EP=6 IP=9 FDC=4
X1 3 2 4 5 1 6 NOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_48 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=4
X1 1 2 3 4 5 1 ICV_47 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_49 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=4
X1 1 2 3 4 5 ICV_23 $T=1140 0 0 0 $X=1025 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_50 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=16
X1 3 4 5 1 2 DLH_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_51
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_52 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=4
X1 1 2 3 4 5 1 ICV_47 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_53 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=4
X1 3 2 4 5 1 1 NOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI222_X1 C2 C1 VSS B1 B2 A2 VDD A1 ZN
** N=14 EP=9 IP=0 FDC=12
M0 10 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=155 $Y=90 $D=1
M1 VSS C1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=345 $Y=90 $D=1
M2 10 B1 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=710 $Y=90 $D=1
M3 11 B2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=900 $Y=90 $D=1
M4 ZN A2 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1090 $Y=90 $D=1
M5 11 A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1280 $Y=90 $D=1
M6 12 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=155 $Y=680 $D=0
M7 ZN C1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=1.9845e-13 AS=8.82e-14 PD=1.89e-06 PS=1.54e-06 $X=345 $Y=680 $D=0
M8 13 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.9845e-13 PD=1.54e-06 PS=1.89e-06 $X=710 $Y=680 $D=0
M9 VDD B2 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=900 $Y=680 $D=0
M10 14 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1090 $Y=680 $D=0
M11 ZN A1 14 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1280 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_54
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_55 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=32
X0 1 2 3 4 5 DLH_X1 $T=0 0 1 180 $X=-2015 $Y=-115
X1 1 6 7 4 5 DLH_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_56
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_57 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=14 FDC=32
X0 1 2 3 4 5 5 NOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 6 7 8 9 2 5 10 5 FA_X1 $T=570 0 0 0 $X=455 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_58 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=8
X0 1 2 3 4 5 5 NOR2_X1 $T=0 0 1 180 $X=-685 $Y=-115
X1 6 2 7 8 5 5 NOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT OR4_X1 A1 A2 A3 A4 VSS VDD ZN
** N=11 EP=7 IP=0 FDC=10
M0 8 A1 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 8 A3 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 VSS A4 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=715 $Y=90 $D=1
M4 ZN 8 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 9 A1 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 10 A2 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 11 A3 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M8 VDD A4 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=715 $Y=995 $D=0
M9 ZN 8 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_59
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_60
** N=2 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT ICV_61 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=4
X1 3 2 4 5 1 1 NOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT CLKBUF_X3 A VSS VDD Z
** N=5 EP=4 IP=0 FDC=8
M0 VSS A 5 VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07 $X=145 $Y=90 $D=1
M1 Z 5 VSS VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=335 $Y=90 $D=1
M2 VSS 5 Z VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=525 $Y=90 $D=1
M3 Z 5 VSS VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=715 $Y=90 $D=1
M4 VDD A 5 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 Z 5 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 VDD 5 Z VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 Z 5 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OR2_X1 A1 A2 VSS VDD ZN
** N=7 EP=5 IP=0 FDC=6
M0 6 A1 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 A1 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR3_X1 A3 VDD A2 A1 VSS ZN
** N=8 EP=6 IP=0 FDC=6
M0 ZN A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 8 A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_62
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT AND3_X1 A1 A2 A3 VSS VDD ZN
** N=9 EP=6 IP=0 FDC=8
M0 8 A1 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 9 A2 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 VSS A3 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=525 $Y=90 $D=1
M3 ZN 7 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 VDD A1 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M5 7 A2 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M6 VDD A3 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=525 $Y=995 $D=0
M7 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_63
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_64
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT MGC_AUTO_NDR_MGC_CLK_NDR_1.0w2.0s_via2_single_MA_north
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3_X1 A3 VSS A2 A1 VDD ZN
** N=8 EP=6 IP=0 FDC=6
M0 7 A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 8 A2 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 VDD A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI22_X1 B2 B1 VSS ZN A1 A2 VDD
** N=10 EP=7 IP=0 FDC=8
M0 VSS B2 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 8 B1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 8 A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 9 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 ZN B1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 10 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 VDD A2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_65
** N=2 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT ICV_66 1 2 3 4 5 6 7 8 9 10 11 12 13
** N=13 EP=13 IP=16 FDC=56
X0 1 2 3 4 5 6 7 13 FA_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 8 9 10 11 5 6 12 13 FA_X1 $T=3040 0 0 0 $X=2925 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_67 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=32
X0 1 2 3 4 5 11 NOR2_X1 $T=3610 0 1 180 $X=2925 $Y=-115
X1 6 7 8 9 2 5 10 11 FA_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT AND4_X1 A1 A2 A3 A4 VSS VDD ZN
** N=11 EP=7 IP=0 FDC=10
M0 9 A1 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 10 A2 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 11 A3 10 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 VSS A4 11 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=715 $Y=90 $D=1
M4 ZN 8 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 8 A1 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD A2 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 8 A3 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M8 VDD A4 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=715 $Y=995 $D=0
M9 ZN 8 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_68
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X32
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_69 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=4
X1 3 2 4 5 1 1 NOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_70 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=16
X0 1 2 3 4 5 DLH_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_71 1 2 3 4 5 6 7
** N=7 EP=7 IP=11 FDC=28
X1 3 4 5 6 2 1 7 1 FA_X1 $T=3230 0 1 180 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_72 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=6
X0 1 2 3 4 5 AND2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_73 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=4
X1 3 2 4 5 1 1 NOR2_X1 $T=950 0 0 0 $X=835 $Y=-115
.ENDS
***************************************
.SUBCKT INV_X8 A ZN VSS VDD
** N=4 EP=4 IP=0 FDC=16
M0 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1095 $Y=90 $D=1
M6 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1285 $Y=90 $D=1
M7 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1475 $Y=90 $D=1
M8 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M9 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M10 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M11 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M12 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
M13 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1095 $Y=680 $D=0
M14 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1285 $Y=680 $D=0
M15 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1475 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_74
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_75 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=32
X0 1 2 3 4 5 11 NOR2_X1 $T=3040 0 0 0 $X=2925 $Y=-115
X1 6 7 8 9 2 5 10 11 FA_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_76
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT NAND2_X1 A2 VSS A1 ZN VDD
** N=6 EP=5 IP=0 FDC=4
M0 6 A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN A1 6 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_77
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_78
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_79
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT OAI211_X1 C2 C1 A VDD B ZN VSS
** N=10 EP=7 IP=0 FDC=8
M0 ZN C2 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 8 C1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 10 A 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS B 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 9 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN C1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 ZN B VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_80
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_81 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=4
X1 3 2 4 5 1 1 NOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_82 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=4
X1 3 2 4 5 1 1 NOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_83 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=4
X1 3 2 4 5 1 1 NOR2_X1 $T=760 0 1 180 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_84
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_85
** N=2 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT XNOR2_X1 VSS A ZN B VDD
** N=9 EP=5 IP=0 FDC=10
M0 9 A 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=155 $Y=90 $D=1
M1 VSS B 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=345 $Y=90 $D=1
M2 7 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=540 $Y=90 $D=1
M3 ZN A 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 7 B ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 6 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=155 $Y=995 $D=0
M6 VDD B 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=345 $Y=995 $D=0
M7 ZN 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=540 $Y=680 $D=0
M8 8 A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M9 VDD B 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_86 1 2 3 4 5 6 7
** N=7 EP=7 IP=11 FDC=28
X1 3 4 5 6 2 1 7 1 FA_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_87 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=8
X0 1 2 3 4 5 5 NOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 6 2 7 8 5 5 NOR2_X1 $T=570 0 0 0 $X=455 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_88 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=14 FDC=32
X0 1 2 3 4 5 5 NOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 6 7 8 9 2 5 10 5 FA_X1 $T=0 0 1 180 $X=-3155 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_89
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_90 1 2 3 4 5 6 7
** N=7 EP=7 IP=11 FDC=28
X1 3 4 5 6 2 1 7 1 FA_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_91 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=11 FDC=28
X0 1 2 3 4 5 6 7 8 FA_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_92 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=28
X1 3 4 5 6 2 1 7 1 FA_X1 $T=380 0 0 0 $X=265 $Y=-115
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_93 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=4
X1 1 2 3 5 4 ICV_81 $T=0 0 0 0 $X=-875 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_94 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=28
X0 1 2 3 4 5 6 7 6 FA_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2_X1 VDD A Z B VSS
** N=9 EP=5 IP=0 FDC=10
M0 6 A VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 9 A Z VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 8 A 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 7 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 7 B Z VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI211_X2 A VDD B C1 ZN C2 VSS
** N=12 EP=7 IP=0 FDC=16
M0 ZN B VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=150 $Y=90 $D=1
M1 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=340 $Y=90 $D=1
M2 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=530 $Y=90 $D=1
M3 VSS B ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=7.2625e-14 AS=5.81e-14 PD=1.18e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 11 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=7.2625e-14 PD=1.11e-06 PS=1.18e-06 $X=945 $Y=90 $D=1
M5 ZN C1 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1135 $Y=90 $D=1
M6 12 C1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1325 $Y=90 $D=1
M7 VSS C2 12 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1515 $Y=90 $D=1
M8 9 B 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=150 $Y=680 $D=0
M9 VDD A 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=340 $Y=680 $D=0
M10 10 A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=530 $Y=680 $D=0
M11 8 B 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=1.1025e-13 AS=8.82e-14 PD=1.61e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M12 ZN C2 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.1025e-13 PD=1.54e-06 PS=1.61e-06 $X=945 $Y=680 $D=0
M13 8 C1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1135 $Y=680 $D=0
M14 ZN C1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1325 $Y=680 $D=0
M15 8 C2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1515 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XOR2_X2 Z B A VSS VDD
** N=10 EP=5 IP=0 FDC=16
M0 7 A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=175 $Y=90 $D=1
M1 VSS B 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=365 $Y=90 $D=1
M2 Z 7 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=555 $Y=90 $D=1
M3 9 A Z VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=745 $Y=90 $D=1
M4 VSS B 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=935 $Y=90 $D=1
M5 10 B VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1125 $Y=90 $D=1
M6 Z A 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1315 $Y=90 $D=1
M7 VSS 7 Z VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1505 $Y=90 $D=1
M8 8 A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=175 $Y=680 $D=0
M9 VDD B 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=365 $Y=680 $D=0
M10 6 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=555 $Y=680 $D=0
M11 Z A 6 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=745 $Y=680 $D=0
M12 6 B Z VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=935 $Y=680 $D=0
M13 Z B 6 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1125 $Y=680 $D=0
M14 6 A Z VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1315 $Y=680 $D=0
M15 VDD 7 6 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1505 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI21_X2 A VDD B1 ZN B2 VSS
** N=9 EP=6 IP=0 FDC=12
M0 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 8 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 9 B1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=945 $Y=90 $D=1
M5 VSS B2 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1135 $Y=90 $D=1
M6 VDD A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M7 7 A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M8 ZN B2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M9 7 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
M10 ZN B1 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=945 $Y=680 $D=0
M11 7 B2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1135 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR2_X2 A1 ZN A2 VSS VDD
** N=7 EP=5 IP=0 FDC=8
M0 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 6 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN A1 6 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 7 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 VDD A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI221_X2 B2 B1 VDD A ZN C1 C2 VSS
** N=14 EP=8 IP=0 FDC=20
M0 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 11 B1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 VSS B2 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 12 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN B1 12 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=6.225e-14 AS=5.81e-14 PD=1.13e-06 PS=1.11e-06 $X=1095 $Y=90 $D=1
M6 13 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=6.225e-14 PD=1.11e-06 PS=1.13e-06 $X=1295 $Y=90 $D=1
M7 ZN C1 13 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1485 $Y=90 $D=1
M8 14 C1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1675 $Y=90 $D=1
M9 VSS C2 14 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1865 $Y=90 $D=1
M10 9 A 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M11 VDD B1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M12 9 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M13 VDD B2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M14 9 B1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
M15 10 A 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=9.45e-14 AS=8.82e-14 PD=1.56e-06 PS=1.54e-06 $X=1095 $Y=680 $D=0
M16 ZN C2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=9.45e-14 PD=1.54e-06 PS=1.56e-06 $X=1295 $Y=680 $D=0
M17 10 C1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1485 $Y=680 $D=0
M18 ZN C1 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1675 $Y=680 $D=0
M19 10 C2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1865 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR3_X4 A1 A2 A3 ZN VDD VSS
** N=8 EP=6 IP=0 FDC=24
M0 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1095 $Y=90 $D=1
M6 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1285 $Y=90 $D=1
M7 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1475 $Y=90 $D=1
M8 ZN A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=1850 $Y=90 $D=1
M9 VSS A3 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=2040 $Y=90 $D=1
M10 ZN A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=2230 $Y=90 $D=1
M11 VSS A3 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=2420 $Y=90 $D=1
M12 ZN A1 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M13 7 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M14 ZN A1 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M15 7 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M16 8 A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
M17 7 A2 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1095 $Y=680 $D=0
M18 8 A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1285 $Y=680 $D=0
M19 7 A2 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1475 $Y=680 $D=0
M20 8 A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=1850 $Y=680 $D=0
M21 VDD A3 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=2040 $Y=680 $D=0
M22 8 A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=2230 $Y=680 $D=0
M23 VDD A3 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=2420 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NAND2_X2 A1 ZN A2 VSS VDD
** N=7 EP=5 IP=0 FDC=8
M0 6 A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 ZN A1 6 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 7 A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=550 $Y=90 $D=1
M3 VSS A2 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=740 $Y=90 $D=1
M4 ZN A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M5 VDD A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M6 ZN A1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=550 $Y=680 $D=0
M7 VDD A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=740 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FPU_VM reset A[0] B[21] B[19] B[23] B[22] A[19] A[17] B[20] A[21] A[20] A[22] B[25] B[24] A[14] A[13] B[11] A[10] B[14] B[9]
+ B[26] B[13] B[8] B[12] B[4] A[25] B[29] A[29] A[30] B[1] A[2] B[5] A[23] B[7] B[10] A[15] A[24] A[6] B[31] A[12]
+ A[3] A[1] A[11] B[27] A[4] A[31] B[18] B[6] B[3] B[16] A[9] A[28] A[26] B[0] A[8] A[27] B[28] B[2] B[17] A[7]
+ A[16] Res[10] Res[12] Res[19] Res[14] Res[22] Res[24] Res[26] Res[13] Res[9] Res[31] Res[16] Res[4] Res[11] Res[27] Res[7] Res[8] Res[18] Res[17] Res[20]
+ Res[23] Res[25] Res[28] enable B[15] Res[0] A[18] A[5] B[30] Res[2] Res[3] Res[5] Res[1] Res[6] Res[15] Res[21] Res[29] Res[30] clk
** N=2528 EP=99 IP=30622 FDC=23226
M0 939 941 931 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=4945 $Y=34095 $D=1
M1 931 64 939 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=5135 $Y=34095 $D=1
M2 939 937 931 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=5325 $Y=34095 $D=1
M3 931 937 939 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=5515 $Y=34095 $D=1
M4 939 64 931 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=5705 $Y=34095 $D=1
M5 931 941 939 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=5895 $Y=34095 $D=1
M6 167 956 931 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=13345 $Y=50895 $D=1
M7 931 956 167 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=13535 $Y=50895 $D=1
M8 956 161 931 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=13725 $Y=50895 $D=1
M9 931 166 956 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=13915 $Y=50895 $D=1
M10 956 143 931 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=14105 $Y=50895 $D=1
M11 931 962 958 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=16195 $Y=59295 $D=1
M12 962 198 931 931 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06 $X=16385 $Y=59500 $D=1
M13 931 201 962 931 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=16575 $Y=59500 $D=1
M14 962 205 931 931 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=16765 $Y=59500 $D=1
M15 2526 966 970 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=17520 $Y=14495 $D=1
M16 931 215 2526 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=17710 $Y=14495 $D=1
M17 2527 215 931 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=6.0175e-14 AS=5.81e-14 PD=1.12e-06 PS=1.11e-06 $X=17900 $Y=14495 $D=1
M18 970 966 2527 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=6.0175e-14 PD=1.11e-06 PS=1.12e-06 $X=18095 $Y=14495 $D=1
M19 155 969 970 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=18285 $Y=14495 $D=1
M20 970 967 155 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=18475 $Y=14495 $D=1
M21 155 967 970 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=18665 $Y=14495 $D=1
M22 970 969 155 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=18855 $Y=14495 $D=1
M23 1004 1002 931 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=30025 $Y=82290 $D=1
M24 931 reset 1004 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=30215 $Y=82290 $D=1
M25 1005 1004 931 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=30405 $Y=82290 $D=1
M26 931 1004 1005 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=30595 $Y=82290 $D=1
M27 931 524 1060 931 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07 $X=55485 $Y=59890 $D=1
M28 1009 1060 931 931 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=55675 $Y=59890 $D=1
M29 931 1060 1009 931 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=55865 $Y=59890 $D=1
M30 931 1077 1079 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=66885 $Y=81695 $D=1
M31 1079 1077 931 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=67075 $Y=81695 $D=1
M32 931 1077 1079 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=67265 $Y=81695 $D=1
M33 1079 1077 931 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=67455 $Y=81695 $D=1
M34 1085 674 1079 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=67645 $Y=81695 $D=1
M35 1079 1084 1085 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=67835 $Y=81695 $D=1
M36 1085 1084 1079 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=68025 $Y=81695 $D=1
M37 1079 674 1085 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=68215 $Y=81695 $D=1
M38 1085 674 1079 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=68405 $Y=81695 $D=1
M39 1079 1084 1085 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=68595 $Y=81695 $D=1
M40 1085 1084 1079 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=68785 $Y=81695 $D=1
M41 1079 674 1085 931 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=68975 $Y=81695 $D=1
M42 2511 941 A[0] A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=4945 $Y=33290 $D=0
M43 2512 64 2511 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=5135 $Y=33290 $D=0
M44 939 937 2512 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=5325 $Y=33290 $D=0
M45 2513 937 939 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=5515 $Y=33290 $D=0
M46 2514 64 2513 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=5705 $Y=33290 $D=0
M47 A[0] 941 2514 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=5895 $Y=33290 $D=0
M48 167 956 A[0] A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=13345 $Y=50090 $D=0
M49 A[0] 956 167 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=13535 $Y=50090 $D=0
M50 2515 161 A[0] A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=13725 $Y=50090 $D=0
M51 2516 166 2515 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=13915 $Y=50090 $D=0
M52 956 143 2516 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=14105 $Y=50090 $D=0
M53 A[0] 962 958 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=16195 $Y=58490 $D=0
M54 2517 198 A[0] A[0] PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.54e-06 $X=16385 $Y=58490 $D=0
M55 2518 201 2517 A[0] PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=16575 $Y=58490 $D=0
M56 962 205 2518 A[0] PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=16765 $Y=58490 $D=0
M57 155 966 A[0] A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=17520 $Y=13690 $D=0
M58 A[0] 215 155 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=17710 $Y=13690 $D=0
M59 155 215 A[0] A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=9.135e-14 AS=8.82e-14 PD=1.55e-06 PS=1.54e-06 $X=17900 $Y=13690 $D=0
M60 A[0] 966 155 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=9.135e-14 PD=1.54e-06 PS=1.55e-06 $X=18095 $Y=13690 $D=0
M61 2519 969 A[0] A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=18285 $Y=13690 $D=0
M62 155 967 2519 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=18475 $Y=13690 $D=0
M63 2520 967 155 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=18665 $Y=13690 $D=0
M64 A[0] 969 2520 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=18855 $Y=13690 $D=0
M65 2521 1002 1004 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=30025 $Y=82880 $D=0
M66 A[0] reset 2521 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=30215 $Y=82880 $D=0
M67 1005 1004 A[0] A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=30405 $Y=82880 $D=0
M68 A[0] 1004 1005 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=30595 $Y=82880 $D=0
M69 A[0] 524 1060 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=55485 $Y=60480 $D=0
M70 1009 1060 A[0] A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=55675 $Y=60480 $D=0
M71 A[0] 1060 1009 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=55865 $Y=60480 $D=0
M72 1085 1077 A[0] A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=66885 $Y=80890 $D=0
M73 A[0] 1077 1085 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=67075 $Y=80890 $D=0
M74 1085 1077 A[0] A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=67265 $Y=80890 $D=0
M75 A[0] 1077 1085 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=67455 $Y=80890 $D=0
M76 2522 674 A[0] A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=67645 $Y=80890 $D=0
M77 1085 1084 2522 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=67835 $Y=80890 $D=0
M78 2523 1084 1085 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=68025 $Y=80890 $D=0
M79 A[0] 674 2523 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=68215 $Y=80890 $D=0
M80 2524 674 A[0] A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=68405 $Y=80890 $D=0
M81 1085 1084 2524 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=68595 $Y=80890 $D=0
M82 2525 1084 1085 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=68785 $Y=80890 $D=0
M83 A[0] 674 2525 A[0] PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=68975 $Y=80890 $D=0
X15374 674 931 A[0] 1002 CLKBUF_X1 $T=37100 73800 0 0 $X=36985 $Y=73685
X15375 2152 931 A[0] 585 CLKBUF_X1 $T=59520 79400 1 0 $X=59405 $Y=77885
X15376 2169 931 A[0] 586 CLKBUF_X1 $T=63700 79400 0 180 $X=63015 $Y=77885
X15377 1860 931 A[0] 621 CLKBUF_X1 $T=63130 82200 0 0 $X=63015 $Y=82085
X15378 1485 931 A[0] 599 CLKBUF_X1 $T=64270 76600 0 180 $X=63585 $Y=75085
X15379 1071 931 A[0] 1099 CLKBUF_X1 $T=64080 37400 0 0 $X=63965 $Y=37285
X15380 1865 931 A[0] 623 CLKBUF_X1 $T=64840 71000 0 180 $X=64155 $Y=69485
X15381 1875 931 A[0] 639 CLKBUF_X1 $T=65030 73800 1 0 $X=64915 $Y=72285
X15382 2331 931 A[0] 2176 CLKBUF_X1 $T=65410 37400 1 0 $X=65295 $Y=35885
X15383 871 931 A[0] 2331 CLKBUF_X1 $T=65410 37400 0 0 $X=65295 $Y=37285
X15384 2332 931 A[0] 831 CLKBUF_X1 $T=65980 37400 1 0 $X=65865 $Y=35885
X15385 1100 931 A[0] 1103 CLKBUF_X1 $T=65980 37400 0 0 $X=65865 $Y=37285
X15386 1569 931 A[0] 2353 CLKBUF_X1 $T=66550 37400 0 0 $X=66435 $Y=37285
X15387 1936 931 A[0] 2363 CLKBUF_X1 $T=67120 37400 0 0 $X=67005 $Y=37285
X15388 2197 931 A[0] 707 CLKBUF_X1 $T=76240 65400 0 180 $X=75555 $Y=63885
X15389 1554 931 A[0] 780 CLKBUF_X1 $T=75670 82200 1 0 $X=75555 $Y=80685
X15390 2347 931 A[0] 743 CLKBUF_X1 $T=76810 45800 1 180 $X=76125 $Y=45685
X15391 2349 931 A[0] 796 CLKBUF_X1 $T=77190 65400 1 0 $X=77075 $Y=63885
X15392 783 931 A[0] 1077 CLKBUF_X1 $T=77760 68200 1 180 $X=77075 $Y=68085
X15393 1565 931 A[0] 810 CLKBUF_X1 $T=78140 82200 0 0 $X=78025 $Y=82085
X15394 1096 931 A[0] 857 CLKBUF_X1 $T=78520 65400 1 0 $X=78405 $Y=63885
X15395 2351 931 A[0] 805 CLKBUF_X1 $T=79470 48600 0 180 $X=78785 $Y=47085
X15396 1928 931 A[0] 1569 CLKBUF_X1 $T=79660 65400 0 180 $X=78975 $Y=63885
X15397 1918 931 A[0] 817 CLKBUF_X1 $T=79660 68200 0 180 $X=78975 $Y=66685
X15398 2354 931 A[0] 795 CLKBUF_X1 $T=80040 54200 1 180 $X=79355 $Y=54085
X15399 1570 931 A[0] 723 CLKBUF_X1 $T=80230 43000 1 180 $X=79545 $Y=42885
X15400 831 931 A[0] 843 CLKBUF_X1 $T=79660 65400 1 0 $X=79545 $Y=63885
X15401 2353 931 A[0] 2209 CLKBUF_X1 $T=79660 65400 0 0 $X=79545 $Y=65285
X15402 832 931 A[0] 912 CLKBUF_X1 $T=79660 68200 1 0 $X=79545 $Y=66685
X15403 2208 931 A[0] 860 CLKBUF_X1 $T=79850 82200 0 0 $X=79735 $Y=82085
X15404 2356 931 A[0] 767 CLKBUF_X1 $T=80800 48600 0 180 $X=80115 $Y=47085
X15405 843 931 A[0] 1071 CLKBUF_X1 $T=80800 65400 1 180 $X=80115 $Y=65285
X15406 2355 931 A[0] 1580 CLKBUF_X1 $T=80230 68200 1 0 $X=80115 $Y=66685
X15407 2358 931 A[0] 733 CLKBUF_X1 $T=81180 59800 0 180 $X=80495 $Y=58285
X15408 1921 931 A[0] 865 CLKBUF_X1 $T=80800 45800 1 0 $X=80685 $Y=44285
X15409 1925 931 A[0] 836 CLKBUF_X1 $T=81370 48600 0 180 $X=80685 $Y=47085
X15410 1931 931 A[0] 808 CLKBUF_X1 $T=81370 51400 1 180 $X=80685 $Y=51285
X15411 1937 931 A[0] 867 CLKBUF_X1 $T=80800 62600 0 0 $X=80685 $Y=62485
X15412 1590 931 A[0] 2332 CLKBUF_X1 $T=81370 65400 1 180 $X=80685 $Y=65285
X15413 1927 931 A[0] 2426 CLKBUF_X1 $T=80800 68200 1 0 $X=80685 $Y=66685
X15414 1574 931 A[0] 818 CLKBUF_X1 $T=81370 71000 0 180 $X=80685 $Y=69485
X15415 1922 931 A[0] 839 CLKBUF_X1 $T=81370 79400 0 180 $X=80685 $Y=77885
X15416 2426 931 A[0] 895 CLKBUF_X1 $T=80990 65400 1 0 $X=80875 $Y=63885
X15417 1919 931 A[0] 822 CLKBUF_X1 $T=81560 71000 1 180 $X=80875 $Y=70885
X15418 1583 931 A[0] 754 CLKBUF_X1 $T=81940 43000 1 180 $X=81255 $Y=42885
X15419 1579 931 A[0] 851 CLKBUF_X1 $T=81370 45800 1 0 $X=81255 $Y=44285
X15420 2215 931 A[0] 811 CLKBUF_X1 $T=81940 48600 0 180 $X=81255 $Y=47085
X15421 1098 931 A[0] 814 CLKBUF_X1 $T=81940 51400 1 180 $X=81255 $Y=51285
X15422 1929 931 A[0] 1927 CLKBUF_X1 $T=81940 62600 1 180 $X=81255 $Y=62485
X15423 enable 931 A[0] 871 CLKBUF_X1 $T=81940 65400 1 180 $X=81255 $Y=65285
X15424 1099 931 A[0] 1928 CLKBUF_X1 $T=81940 68200 0 180 $X=81255 $Y=66685
X15425 872 931 A[0] 899 CLKBUF_X1 $T=81370 71000 1 0 $X=81255 $Y=69485
X15426 2359 931 A[0] 913 CLKBUF_X1 $T=81370 79400 0 0 $X=81255 $Y=79285
X15427 1580 931 A[0] 1929 CLKBUF_X1 $T=82130 68200 1 180 $X=81445 $Y=68085
X15428 1935 931 A[0] 854 CLKBUF_X1 $T=81940 54200 0 0 $X=81825 $Y=54085
X15429 1586 931 A[0] 790 CLKBUF_X1 $T=82700 45800 1 180 $X=82015 $Y=45685
X15430 2221 931 A[0] 745 CLKBUF_X1 $T=82890 54200 0 180 $X=82205 $Y=52685
X15431 1932 931 A[0] 855 CLKBUF_X1 $T=82890 57000 1 180 $X=82205 $Y=56885
X15432 2363 931 A[0] 1590 CLKBUF_X1 $T=82890 65400 0 180 $X=82205 $Y=63885
X15433 1596 931 A[0] 1934 CLKBUF_X1 $T=82890 65400 1 180 $X=82205 $Y=65285
X15434 2214 931 A[0] 819 CLKBUF_X1 $T=82890 76600 0 180 $X=82205 $Y=75085
X15435 2362 931 A[0] 901 CLKBUF_X1 $T=82320 82200 0 0 $X=82205 $Y=82085
X15436 1102 931 A[0] 908 CLKBUF_X1 $T=82700 45800 1 0 $X=82585 $Y=44285
X15437 887 931 A[0] 897 CLKBUF_X1 $T=82700 45800 0 0 $X=82585 $Y=45685
X15438 889 931 A[0] 909 CLKBUF_X1 $T=82700 48600 0 0 $X=82585 $Y=48485
X15439 2218 931 A[0] 852 CLKBUF_X1 $T=83270 51400 1 180 $X=82585 $Y=51285
X15440 2364 931 A[0] 856 CLKBUF_X1 $T=83270 59800 0 180 $X=82585 $Y=58285
X15441 2219 931 A[0] 842 CLKBUF_X1 $T=83270 73800 0 180 $X=82585 $Y=72285
X15442 1593 931 A[0] 765 CLKBUF_X1 $T=83460 59800 1 180 $X=82775 $Y=59685
X15443 1595 931 A[0] 1936 CLKBUF_X1 $T=83460 65400 0 180 $X=82775 $Y=63885
X15444 895 931 A[0] 911 CLKBUF_X1 $T=82890 65400 0 0 $X=82775 $Y=65285
X15445 2220 931 A[0] 898 CLKBUF_X1 $T=83650 48600 0 180 $X=82965 $Y=47085
X15446 1588 931 A[0] 789 CLKBUF_X1 $T=83650 51400 0 180 $X=82965 $Y=49885
X15447 1940 931 A[0] 815 CLKBUF_X1 $T=83650 57000 1 180 $X=82965 $Y=56885
X15448 1933 931 A[0] 816 CLKBUF_X1 $T=83650 62600 0 180 $X=82965 $Y=61085
X15449 1597 931 A[0] 858 CLKBUF_X1 $T=83650 71000 1 180 $X=82965 $Y=70885
X15450 2217 931 A[0] 885 CLKBUF_X1 $T=83840 76600 0 180 $X=83155 $Y=75085
X15451 2367 931 A[0] 837 CLKBUF_X1 $T=84030 54200 1 180 $X=83345 $Y=54085
X15452 1104 931 A[0] 741 CLKBUF_X1 $T=84030 59800 1 180 $X=83345 $Y=59685
X15453 2176 931 A[0] 1595 CLKBUF_X1 $T=84030 65400 0 180 $X=83345 $Y=63885
X15454 911 931 A[0] 1596 CLKBUF_X1 $T=83460 65400 0 0 $X=83345 $Y=65285
X15455 1103 931 A[0] 2355 CLKBUF_X1 $T=84030 71000 0 180 $X=83345 $Y=69485
X15456 1585 931 A[0] 803 CLKBUF_X1 $T=84410 76600 0 180 $X=83725 $Y=75085
X15549 93 11 931 A[0] 27 AND2_X1 $T=3090 37400 1 180 $X=2215 $Y=37285
X15550 93 12 931 A[0] 5 AND2_X1 $T=3090 40200 0 180 $X=2215 $Y=38685
X15551 93 14 931 A[0] 6 AND2_X1 $T=3090 48600 1 180 $X=2215 $Y=48485
X15552 93 10 931 A[0] 28 AND2_X1 $T=2330 51400 0 0 $X=2215 $Y=51285
X15553 93 54 931 A[0] 36 AND2_X1 $T=5940 51400 1 180 $X=5065 $Y=51285
X15554 93 65 931 A[0] 46 AND2_X1 $T=5940 51400 0 0 $X=5825 $Y=51285
X15555 948 78 931 A[0] 48 AND2_X1 $T=6700 43000 0 0 $X=6585 $Y=42885
X15556 93 97 931 A[0] 89 AND2_X1 $T=8980 54200 1 180 $X=8105 $Y=54085
X15557 93 103 931 A[0] 96 AND2_X1 $T=9360 48600 1 180 $X=8485 $Y=48485
X15558 93 118 931 A[0] 105 AND2_X1 $T=10880 62600 0 180 $X=10005 $Y=61085
X15559 93 123 931 A[0] 117 AND2_X1 $T=11070 59800 0 180 $X=10195 $Y=58285
X15560 93 125 931 A[0] 113 AND2_X1 $T=11640 57000 1 180 $X=10765 $Y=56885
X15561 93 130 931 A[0] 112 AND2_X1 $T=11830 54200 1 180 $X=10955 $Y=54085
X15562 93 134 931 A[0] 139 AND2_X1 $T=11450 62600 0 0 $X=11335 $Y=62485
X15563 93 178 931 A[0] 162 AND2_X1 $T=15440 76600 1 180 $X=14565 $Y=76485
X15564 93 179 931 A[0] 158 AND2_X1 $T=15630 71000 1 180 $X=14755 $Y=70885
X15565 93 180 931 A[0] 181 AND2_X1 $T=15630 73800 1 180 $X=14755 $Y=73685
X15566 93 186 931 A[0] 190 AND2_X1 $T=15250 65400 1 0 $X=15135 $Y=63885
X15567 931 192 931 A[0] 138 AND2_X1 $T=15820 48600 0 0 $X=15705 $Y=48485
X15568 1219 152 931 A[0] 214 AND2_X1 $T=16010 57000 0 0 $X=15895 $Y=56885
X15569 93 209 931 A[0] 213 AND2_X1 $T=16960 73800 0 0 $X=16845 $Y=73685
X15570 93 225 931 A[0] 226 AND2_X1 $T=18290 82200 1 0 $X=18175 $Y=80685
X15571 93 271 931 A[0] 257 AND2_X1 $T=22470 82200 0 180 $X=21595 $Y=80685
X15572 93 295 931 A[0] 288 AND2_X1 $T=24940 82200 0 180 $X=24065 $Y=80685
X15573 1271 301 931 A[0] 273 AND2_X1 $T=25510 73800 0 180 $X=24635 $Y=72285
X15574 292 302 931 A[0] 1710 AND2_X1 $T=24940 76600 0 0 $X=24825 $Y=76485
X15575 93 320 931 A[0] 328 AND2_X1 $T=27220 82200 1 0 $X=27105 $Y=80685
X15576 538 547 931 A[0] 2403 AND2_X1 $T=57620 73800 1 0 $X=57505 $Y=72285
X15577 538 551 931 A[0] 541 AND2_X1 $T=58570 73800 1 180 $X=57695 $Y=73685
X15578 538 573 931 A[0] 550 AND2_X1 $T=60090 71000 1 180 $X=59215 $Y=70885
X15579 538 579 931 A[0] 583 AND2_X1 $T=60660 68200 1 0 $X=60545 $Y=66685
X15580 538 590 931 A[0] 580 AND2_X1 $T=61040 71000 0 0 $X=60925 $Y=70885
X15581 538 598 931 A[0] 595 AND2_X1 $T=63130 62600 1 180 $X=62255 $Y=62485
X15582 1077 B[22] 931 A[0] 2169 AND2_X1 $T=63130 79400 0 180 $X=62255 $Y=77885
X15583 1077 B[23] 931 A[0] 1860 AND2_X1 $T=62370 82200 0 0 $X=62255 $Y=82085
X15584 1077 A[19] 931 A[0] 1485 AND2_X1 $T=62940 76600 1 0 $X=62825 $Y=75085
X15585 1077 A[17] 931 A[0] 1865 AND2_X1 $T=63700 71000 0 0 $X=63585 $Y=70885
X15586 538 625 931 A[0] 616 AND2_X1 $T=65030 68200 0 180 $X=64155 $Y=66685
X15587 538 629 931 A[0] 582 AND2_X1 $T=64840 65400 1 0 $X=64725 $Y=63885
X15588 538 635 931 A[0] 617 AND2_X1 $T=65600 71000 0 180 $X=64725 $Y=69485
X15589 538 665 931 A[0] 652 AND2_X1 $T=68070 54200 1 180 $X=67195 $Y=54085
X15590 538 672 931 A[0] 613 AND2_X1 $T=67690 57000 1 0 $X=67575 $Y=55485
X15591 538 681 931 A[0] 668 AND2_X1 $T=69590 45800 1 180 $X=68715 $Y=45685
X15592 538 684 931 A[0] 651 AND2_X1 $T=69210 48600 1 0 $X=69095 $Y=47085
X15593 538 687 931 A[0] 678 AND2_X1 $T=70160 65400 0 180 $X=69285 $Y=63885
X15594 538 694 931 A[0] 669 AND2_X1 $T=70540 59800 1 180 $X=69665 $Y=59685
X15595 538 693 931 A[0] 633 AND2_X1 $T=69970 59800 1 0 $X=69855 $Y=58285
X15596 538 695 931 A[0] 657 AND2_X1 $T=69970 62600 0 0 $X=69855 $Y=62485
X15597 538 699 931 A[0] 676 AND2_X1 $T=71110 51400 0 180 $X=70235 $Y=49885
X15598 538 703 931 A[0] 677 AND2_X1 $T=71300 54200 0 180 $X=70425 $Y=52685
X15599 538 700 931 A[0] 615 AND2_X1 $T=70540 59800 0 0 $X=70425 $Y=59685
X15600 538 706 931 A[0] 666 AND2_X1 $T=70920 62600 1 0 $X=70805 $Y=61085
X15601 538 708 931 A[0] 685 AND2_X1 $T=71680 65400 1 180 $X=70805 $Y=65285
X15602 1534 710 931 A[0] 736 AND2_X1 $T=71110 73800 1 0 $X=70995 $Y=72285
X15603 538 715 931 A[0] 712 AND2_X1 $T=72250 37400 0 180 $X=71375 $Y=35885
X15604 538 716 931 A[0] 698 AND2_X1 $T=72250 43000 1 180 $X=71375 $Y=42885
X15605 538 717 931 A[0] 675 AND2_X1 $T=72440 43000 0 180 $X=71565 $Y=41485
X15606 538 719 931 A[0] 697 AND2_X1 $T=72630 37400 1 180 $X=71755 $Y=37285
X15607 538 721 931 A[0] 705 AND2_X1 $T=72630 59800 0 180 $X=71755 $Y=58285
X15608 538 728 931 A[0] 726 AND2_X1 $T=73010 54200 0 0 $X=72895 $Y=54085
X15609 538 738 931 A[0] 689 AND2_X1 $T=74720 34600 0 180 $X=73845 $Y=33085
X15610 538 740 931 A[0] 773 AND2_X1 $T=74910 34600 1 180 $X=74035 $Y=34485
X15611 538 749 931 A[0] 748 AND2_X1 $T=74910 34600 0 0 $X=74795 $Y=34485
X15612 1077 A[22] 931 A[0] 2197 AND2_X1 $T=74910 65400 1 0 $X=74795 $Y=63885
X15613 538 755 931 A[0] 725 AND2_X1 $T=75100 48600 1 0 $X=74985 $Y=47085
X15614 538 758 931 A[0] 764 AND2_X1 $T=75860 51400 1 180 $X=74985 $Y=51285
X15615 538 761 931 A[0] 729 AND2_X1 $T=76050 57000 1 180 $X=75175 $Y=56885
X15616 538 760 931 A[0] 696 AND2_X1 $T=75480 57000 1 0 $X=75365 $Y=55485
X15617 538 774 931 A[0] 794 AND2_X1 $T=76240 34600 0 0 $X=76125 $Y=34485
X15618 538 775 931 A[0] 731 AND2_X1 $T=76240 40200 1 0 $X=76125 $Y=38685
X15619 1077 B[25] 931 A[0] 1554 AND2_X1 $T=77000 82200 0 180 $X=76125 $Y=80685
X15620 538 785 931 A[0] 800 AND2_X1 $T=77000 34600 0 0 $X=76885 $Y=34485
X15621 1077 B[24] 931 A[0] 1565 AND2_X1 $T=77380 82200 1 0 $X=77265 $Y=80685
X15622 1077 A[14] 931 A[0] 1096 AND2_X1 $T=77760 65400 1 0 $X=77645 $Y=63885
X15623 820 799 931 A[0] 2205 AND2_X1 $T=78900 23400 1 180 $X=78025 $Y=23285
X15624 870 B[9] 931 A[0] 2347 AND2_X1 $T=79470 45800 1 180 $X=78595 $Y=45685
X15625 1077 A[10] 931 A[0] 2206 AND2_X1 $T=78710 62600 1 0 $X=78595 $Y=61085
X15626 870 B[14] 931 A[0] 1570 AND2_X1 $T=78900 43000 0 0 $X=78785 $Y=42885
X15627 538 827 931 A[0] 848 AND2_X1 $T=79850 34600 0 180 $X=78975 $Y=33085
X15628 1077 B[26] 931 A[0] 2208 AND2_X1 $T=79090 82200 0 0 $X=78975 $Y=82085
X15629 870 B[8] 931 A[0] 2351 AND2_X1 $T=80230 45800 1 180 $X=79355 $Y=45685
X15630 870 B[13] 931 A[0] 2356 AND2_X1 $T=79470 48600 1 0 $X=79355 $Y=47085
X15631 870 B[4] 931 A[0] 1579 AND2_X1 $T=80040 45800 1 0 $X=79925 $Y=44285
X15632 1077 B[29] 931 A[0] 1574 AND2_X1 $T=80800 71000 0 180 $X=79925 $Y=69485
X15633 1077 A[25] 931 A[0] 1922 AND2_X1 $T=80040 79400 1 0 $X=79925 $Y=77885
X15634 1077 A[29] 931 A[0] 1918 AND2_X1 $T=80990 65400 0 180 $X=80115 $Y=63885
X15635 1077 A[30] 931 A[0] 1919 AND2_X1 $T=80990 71000 1 180 $X=80115 $Y=70885
X15636 538 844 931 A[0] 850 AND2_X1 $T=80420 37400 1 0 $X=80305 $Y=35885
X15637 870 B[1] 931 A[0] 1583 AND2_X1 $T=80610 43000 0 0 $X=80495 $Y=42885
X15638 870 A[2] 931 A[0] 1921 AND2_X1 $T=81370 45800 1 180 $X=80495 $Y=45685
X15639 538 876 931 A[0] 849 AND2_X1 $T=81940 34600 0 180 $X=81065 $Y=33085
X15640 870 B[10] 931 A[0] 1925 AND2_X1 $T=81940 48600 1 180 $X=81065 $Y=48485
X15641 870 B[15] 931 A[0] 2354 AND2_X1 $T=81940 57000 0 180 $X=81065 $Y=55485
X15642 870 A[15] 931 A[0] 2358 AND2_X1 $T=81940 59800 0 180 $X=81065 $Y=58285
X15643 1077 A[23] 931 A[0] 1585 AND2_X1 $T=81180 76600 1 0 $X=81065 $Y=75085
X15644 870 B[7] 931 A[0] 1586 AND2_X1 $T=81370 45800 0 0 $X=81255 $Y=45685
X15645 1077 A[24] 931 A[0] 2214 AND2_X1 $T=81370 79400 1 0 $X=81255 $Y=77885
X15646 870 A[6] 931 A[0] 1588 AND2_X1 $T=81560 51400 1 0 $X=81445 $Y=49885
X15647 1077 B[31] 931 A[0] 832 AND2_X1 $T=82320 65400 0 180 $X=81445 $Y=63885
X15648 870 A[12] 931 A[0] 1593 AND2_X1 $T=82130 59800 0 0 $X=82015 $Y=59685
X15649 538 886 931 A[0] 893 AND2_X1 $T=82320 34600 1 0 $X=82205 $Y=33085
X15650 870 A[3] 931 A[0] 2215 AND2_X1 $T=83080 48600 0 180 $X=82205 $Y=47085
X15651 870 A[1] 931 A[0] 1931 AND2_X1 $T=83080 51400 0 180 $X=82205 $Y=49885
X15652 870 A[5] 931 A[0] 1932 AND2_X1 $T=83080 57000 0 180 $X=82205 $Y=55485
X15653 870 A[11] 931 A[0] 1933 AND2_X1 $T=83080 62600 0 180 $X=82205 $Y=61085
X15654 1077 B[27] 931 A[0] 2362 AND2_X1 $T=83080 79400 1 180 $X=82205 $Y=79285
X15655 870 A[4] 931 A[0] 1935 AND2_X1 $T=83270 54200 1 180 $X=82395 $Y=54085
X15656 1077 A[31] 931 A[0] 872 AND2_X1 $T=83460 71000 0 180 $X=82585 $Y=69485
X15657 870 B[18] 931 A[0] 1098 AND2_X1 $T=83650 54200 0 180 $X=82775 $Y=52685
X15658 538 907 931 A[0] 896 AND2_X1 $T=83080 34600 1 0 $X=82965 $Y=33085
X15659 870 B[6] 931 A[0] 1102 AND2_X1 $T=83270 45800 1 0 $X=83155 $Y=44285
X15660 870 B[3] 931 A[0] 887 AND2_X1 $T=83270 45800 0 0 $X=83155 $Y=45685
X15661 870 B[0] 931 A[0] 889 AND2_X1 $T=84030 48600 1 180 $X=83155 $Y=48485
X15662 870 A[0] 931 A[0] 2218 AND2_X1 $T=83270 51400 0 0 $X=83155 $Y=51285
X15663 870 B[16] 931 A[0] 2367 AND2_X1 $T=83270 57000 1 0 $X=83155 $Y=55485
X15664 870 A[9] 931 A[0] 2364 AND2_X1 $T=83270 59800 1 0 $X=83155 $Y=58285
X15665 1077 A[28] 931 A[0] 2219 AND2_X1 $T=83270 73800 1 0 $X=83155 $Y=72285
X15666 1077 A[27] 931 A[0] 2217 AND2_X1 $T=84030 73800 1 180 $X=83155 $Y=73685
X15667 1077 A[26] 931 A[0] 2359 AND2_X1 $T=83270 79400 0 0 $X=83155 $Y=79285
X15668 870 B[2] 931 A[0] 2220 AND2_X1 $T=83650 48600 1 0 $X=83535 $Y=47085
X15669 870 B[17] 931 A[0] 2221 AND2_X1 $T=83650 54200 1 0 $X=83535 $Y=52685
X15670 870 A[7] 931 A[0] 1940 AND2_X1 $T=83650 57000 0 0 $X=83535 $Y=56885
X15671 870 A[16] 931 A[0] 1104 AND2_X1 $T=83650 62600 1 0 $X=83535 $Y=61085
X15672 1077 B[30] 931 A[0] 1597 AND2_X1 $T=83650 71000 0 0 $X=83535 $Y=70885
X15828 2231 2235 931 A[0] INV_X2 $T=9170 37400 0 0 $X=9055 $Y=37285
X15829 1438 995 931 A[0] INV_X2 $T=56100 76600 1 0 $X=55985 $Y=75085
X15830 1449 980 931 A[0] INV_X2 $T=57430 71000 1 180 $X=56745 $Y=70885
X15831 1469 1014 931 A[0] INV_X2 $T=59710 68200 1 180 $X=59025 $Y=68085
X15832 1465 1022 931 A[0] INV_X2 $T=60090 65400 0 180 $X=59405 $Y=63885
X15833 1467 973 931 A[0] INV_X2 $T=60850 62600 0 180 $X=60165 $Y=61085
X15834 1482 931 931 A[0] INV_X2 $T=62940 71000 1 0 $X=62825 $Y=69485
X15835 2333 660 931 A[0] INV_X2 $T=66550 65400 1 180 $X=65865 $Y=65285
X15836 1083 664 931 A[0] INV_X2 $T=68070 57000 0 0 $X=67955 $Y=56885
X15837 2346 788 931 A[0] INV_X2 $T=74150 31800 0 0 $X=74035 $Y=31685
X15838 1905 1011 931 A[0] INV_X2 $T=74530 29000 0 0 $X=74415 $Y=28885
X15839 2352 1029 931 A[0] INV_X2 $T=79660 29000 0 180 $X=78975 $Y=27485
X15840 2366 997 931 A[0] INV_X2 $T=83460 26200 1 0 $X=83345 $Y=24685
X16558 1857 931 A[0] 584 1077 B[19] 1857 ICV_16 $T=62180 76600 0 180 $X=61495 $Y=75085
X16559 2486 931 A[0] 618 1077 B[20] 2486 ICV_16 $T=64270 73800 1 180 $X=63585 $Y=73685
X16560 2178 931 A[0] 634 1077 A[20] 2178 ICV_16 $T=66550 71000 0 180 $X=65865 $Y=69485
X16561 1915 931 A[0] 777 1077 A[13] 1915 ICV_16 $T=77950 62600 0 180 $X=77265 $Y=61085
X16562 1916 931 A[0] 702 870 B[11] 1916 ICV_16 $T=78140 48600 0 180 $X=77455 $Y=47085
X16563 1571 931 A[0] 768 870 B[12] 1571 ICV_16 $T=79470 51400 0 180 $X=78785 $Y=49885
X16564 2206 931 A[0] 802 1077 A[18] 2349 ICV_16 $T=80040 62600 1 180 $X=79355 $Y=62485
X16565 2211 931 A[0] 828 870 B[5] 2211 ICV_16 $T=80800 51400 0 180 $X=80115 $Y=49885
X16566 2209 931 A[0] 1100 870 A[8] 1937 ICV_16 $T=83270 62600 1 180 $X=82585 $Y=62485
X16567 1938 931 A[0] 859 1077 B[28] 1938 ICV_16 $T=83270 76600 1 180 $X=82585 $Y=76485
X16868 104 1941 5 931 A[0] DLH_X1 $T=1000 40200 0 0 $X=885 $Y=40085
X16869 104 29 6 931 A[0] DLH_X1 $T=1000 51400 1 0 $X=885 $Y=49885
X16870 1005 Res[2] 8 931 A[0] DLH_X1 $T=1000 65400 1 0 $X=885 $Y=63885
X16871 1005 Res[10] 3 931 A[0] DLH_X1 $T=2900 68200 1 180 $X=885 $Y=68085
X16872 1005 Res[8] 4 931 A[0] DLH_X1 $T=2900 73800 1 180 $X=885 $Y=73685
X16873 1005 Res[7] 9 931 A[0] DLH_X1 $T=1000 79400 1 0 $X=885 $Y=77885
X16874 1005 Res[3] 30 931 A[0] DLH_X1 $T=2330 59800 1 0 $X=2215 $Y=58285
X16875 1005 Res[6] 26 931 A[0] DLH_X1 $T=4230 71000 1 180 $X=2215 $Y=70885
X16876 1005 Res[16] 32 931 A[0] DLH_X1 $T=2330 76600 1 0 $X=2215 $Y=75085
X16877 104 55 36 931 A[0] DLH_X1 $T=2900 54200 0 0 $X=2785 $Y=54085
X16878 1005 Res[13] 39 931 A[0] DLH_X1 $T=3470 73800 1 0 $X=3355 $Y=72285
X16879 1005 Res[18] 45 931 A[0] DLH_X1 $T=3850 82200 0 0 $X=3735 $Y=82085
X16880 1005 Res[11] 51 931 A[0] DLH_X1 $T=4230 65400 0 0 $X=4115 $Y=65285
X16881 1005 Res[12] 66 931 A[0] DLH_X1 $T=5180 68200 0 0 $X=5065 $Y=68085
X16882 1005 Res[9] 69 931 A[0] DLH_X1 $T=5370 73800 1 0 $X=5255 $Y=72285
X16883 1005 Res[17] 72 931 A[0] DLH_X1 $T=7650 82200 1 180 $X=5635 $Y=82085
X16884 1005 Res[19] 84 931 A[0] DLH_X1 $T=6130 82200 1 0 $X=6015 $Y=80685
X16885 1005 Res[15] 98 931 A[0] DLH_X1 $T=9740 76600 1 180 $X=7725 $Y=76485
X16886 104 106 113 931 A[0] DLH_X1 $T=8980 57000 0 0 $X=8865 $Y=56885
X16887 1005 Res[14] 140 931 A[0] DLH_X1 $T=10880 76600 0 0 $X=10765 $Y=76485
X16888 104 67 162 931 A[0] DLH_X1 $T=12780 76600 0 0 $X=12665 $Y=76485
X16889 104 124 190 931 A[0] DLH_X1 $T=16960 65400 1 180 $X=14945 $Y=65285
X16890 104 114 200 931 A[0] DLH_X1 $T=15440 79400 0 0 $X=15325 $Y=79285
X16891 1005 Res[22] 202 931 A[0] DLH_X1 $T=17720 82200 1 180 $X=15705 $Y=82085
X16892 104 92 226 931 A[0] DLH_X1 $T=19620 82200 1 180 $X=17605 $Y=82085
X16893 104 2012 288 931 A[0] DLH_X1 $T=22280 82200 0 0 $X=22165 $Y=82085
X16894 104 543 328 931 A[0] DLH_X1 $T=29880 82200 1 180 $X=27865 $Y=82085
X16895 1436 1438 541 931 A[0] DLH_X1 $T=55910 73800 0 0 $X=55795 $Y=73685
X16896 1436 1447 550 931 A[0] DLH_X1 $T=57240 68200 0 0 $X=57125 $Y=68085
X16897 1436 1449 2403 931 A[0] DLH_X1 $T=57430 71000 0 0 $X=57315 $Y=70885
X16898 1436 1067 578 931 A[0] DLH_X1 $T=61990 59800 1 180 $X=59975 $Y=59685
X16899 1436 1469 580 931 A[0] DLH_X1 $T=61990 68200 1 180 $X=59975 $Y=68085
X16900 1436 1467 595 931 A[0] DLH_X1 $T=61230 62600 1 0 $X=61115 $Y=61085
X16901 883 579 599 931 A[0] DLH_X1 $T=61800 71000 0 0 $X=61685 $Y=70885
X16902 1436 1477 616 931 A[0] DLH_X1 $T=62370 68200 1 0 $X=62255 $Y=66685
X16903 1005 Res[29] 619 931 A[0] DLH_X1 $T=62370 76600 0 0 $X=62255 $Y=76485
X16904 883 747 621 931 A[0] DLH_X1 $T=64840 82200 0 180 $X=62825 $Y=80685
X16905 883 598 623 931 A[0] DLH_X1 $T=63130 62600 0 0 $X=63015 $Y=62485
X16906 883 625 634 931 A[0] DLH_X1 $T=64270 68200 0 0 $X=64155 $Y=68085
X16907 883 635 639 931 A[0] DLH_X1 $T=64460 71000 0 0 $X=64345 $Y=70885
X16908 1436 2177 651 931 A[0] DLH_X1 $T=65410 48600 0 0 $X=65295 $Y=48485
X16909 1436 1500 652 931 A[0] DLH_X1 $T=65410 54200 0 0 $X=65295 $Y=54085
X16910 1005 Res[30] 662 931 A[0] DLH_X1 $T=66360 71000 0 0 $X=66245 $Y=70885
X16911 1436 1506 666 931 A[0] DLH_X1 $T=66740 62600 1 0 $X=66625 $Y=61085
X16912 1436 1877 667 931 A[0] DLH_X1 $T=66930 43000 0 0 $X=66815 $Y=42885
X16913 1436 2335 668 931 A[0] DLH_X1 $T=66930 45800 0 0 $X=66815 $Y=45685
X16914 1436 1878 669 931 A[0] DLH_X1 $T=66930 59800 0 0 $X=66815 $Y=59685
X16915 1436 1512 676 931 A[0] DLH_X1 $T=67500 51400 1 0 $X=67385 $Y=49885
X16916 1436 1513 677 931 A[0] DLH_X1 $T=67500 54200 1 0 $X=67385 $Y=52685
X16917 1436 2333 678 931 A[0] DLH_X1 $T=67500 65400 1 0 $X=67385 $Y=63885
X16918 1436 1521 675 931 A[0] DLH_X1 $T=69590 40200 0 180 $X=67575 $Y=38685
X16919 1436 1517 685 931 A[0] DLH_X1 $T=70540 68200 0 180 $X=68525 $Y=66685
X16920 1005 Res[27] 688 931 A[0] DLH_X1 $T=68830 82200 0 0 $X=68715 $Y=82085
X16921 1436 2415 689 931 A[0] DLH_X1 $T=71110 31800 0 180 $X=69095 $Y=30285
X16922 1436 1524 696 931 A[0] DLH_X1 $T=69400 57000 1 0 $X=69285 $Y=55485
X16923 1436 1886 697 931 A[0] DLH_X1 $T=69590 37400 1 0 $X=69475 $Y=35885
X16924 1436 1522 698 931 A[0] DLH_X1 $T=69780 43000 1 0 $X=69665 $Y=41485
X16925 883 681 702 931 A[0] DLH_X1 $T=69970 48600 1 0 $X=69855 $Y=47085
X16926 883 629 707 931 A[0] DLH_X1 $T=70160 65400 1 0 $X=70045 $Y=63885
X16927 1436 1535 720 931 A[0] DLH_X1 $T=71300 48600 0 0 $X=71185 $Y=48485
X16928 883 683 723 931 A[0] DLH_X1 $T=73770 45800 0 180 $X=71755 $Y=44285
X16929 1436 1896 726 931 A[0] DLH_X1 $T=72060 51400 0 0 $X=71945 $Y=51285
X16930 1436 1902 731 931 A[0] DLH_X1 $T=74530 37400 1 180 $X=72515 $Y=37285
X16931 883 706 733 931 A[0] DLH_X1 $T=72630 59800 1 0 $X=72515 $Y=58285
X16932 883 703 745 931 A[0] DLH_X1 $T=73960 54200 1 0 $X=73845 $Y=52685
X16933 883 749 754 931 A[0] DLH_X1 $T=74340 40200 1 0 $X=74225 $Y=38685
X16934 1436 1910 764 931 A[0] DLH_X1 $T=74910 43000 0 0 $X=74795 $Y=42885
X16935 883 699 768 931 A[0] DLH_X1 $T=75290 51400 1 0 $X=75175 $Y=49885
X16936 1005 Res[0] 766 931 A[0] DLH_X1 $T=77190 65400 1 180 $X=75175 $Y=65285
X16937 883 756 780 931 A[0] DLH_X1 $T=75670 82200 0 0 $X=75555 $Y=82085
X16938 883 715 789 931 A[0] DLH_X1 $T=78710 43000 1 180 $X=76695 $Y=42885
X16939 883 719 790 931 A[0] DLH_X1 $T=78710 45800 1 180 $X=76695 $Y=45685
X16940 1005 Res[31] 792 931 A[0] DLH_X1 $T=76810 68200 1 0 $X=76695 $Y=66685
X16941 1436 1562 794 931 A[0] DLH_X1 $T=77190 34600 1 0 $X=77075 $Y=33085
X16942 883 708 796 931 A[0] DLH_X1 $T=77190 65400 0 0 $X=77075 $Y=65285
X16943 883 694 802 931 A[0] DLH_X1 $T=77570 62600 0 0 $X=77455 $Y=62485
X16944 883 557 803 931 A[0] DLH_X1 $T=77570 76600 1 0 $X=77455 $Y=75085
X16945 883 654 814 931 A[0] DLH_X1 $T=78140 54200 1 0 $X=78025 $Y=52685
X16946 883 769 817 931 A[0] DLH_X1 $T=78140 68200 0 0 $X=78025 $Y=68085
X16947 883 787 819 931 A[0] DLH_X1 $T=78140 76600 0 0 $X=78025 $Y=76485
X16948 883 734 810 931 A[0] DLH_X1 $T=80040 82200 0 180 $X=78025 $Y=80685
X16949 883 738 811 931 A[0] DLH_X1 $T=80230 40200 1 180 $X=78215 $Y=40085
X16950 883 740 828 931 A[0] DLH_X1 $T=78520 37400 1 0 $X=78405 $Y=35885
X16951 883 776 842 931 A[0] DLH_X1 $T=79470 73800 0 0 $X=79355 $Y=73685
X16952 883 758 855 931 A[0] DLH_X1 $T=80040 54200 0 0 $X=79925 $Y=54085
X16953 883 722 860 931 A[0] DLH_X1 $T=80040 82200 1 0 $X=79925 $Y=80685
X16954 1436 931 849 931 A[0] DLH_X1 $T=82130 31800 1 180 $X=80115 $Y=31685
X16955 883 774 865 931 A[0] DLH_X1 $T=80230 40200 0 0 $X=80115 $Y=40085
X16956 883 778 885 931 A[0] DLH_X1 $T=81370 73800 0 0 $X=81255 $Y=73685
X16957 1436 2366 893 931 A[0] DLH_X1 $T=84030 26200 1 180 $X=82015 $Y=26085
X16958 883 844 908 931 A[0] DLH_X1 $T=82320 40200 1 0 $X=82205 $Y=38685
X16959 883 840 912 931 A[0] DLH_X1 $T=82320 68200 1 0 $X=82205 $Y=66685
X17096 1447 986 931 A[0] INV_X4 $T=57620 71000 0 180 $X=56555 $Y=69485
X17097 1453 392 931 A[0] INV_X4 $T=58380 68200 1 0 $X=58265 $Y=66685
X17098 1067 503 931 A[0] INV_X4 $T=60660 59800 0 180 $X=59595 $Y=58285
X17099 1477 399 931 A[0] INV_X4 $T=62370 68200 0 180 $X=61305 $Y=66685
X17100 1483 1000 931 A[0] INV_X4 $T=63130 62600 1 0 $X=63015 $Y=61085
X17101 1488 501 931 A[0] INV_X4 $T=64270 59800 1 0 $X=64155 $Y=58285
X17102 1504 985 931 A[0] INV_X4 $T=65980 62600 1 180 $X=64915 $Y=62485
X17103 2177 975 931 A[0] INV_X4 $T=65790 48600 1 0 $X=65675 $Y=47085
X17104 1506 448 931 A[0] INV_X4 $T=66740 62600 0 180 $X=65675 $Y=61085
X17105 1877 976 931 A[0] INV_X4 $T=66930 43000 1 180 $X=65865 $Y=42885
X17106 2335 655 931 A[0] INV_X4 $T=66930 45800 1 180 $X=65865 $Y=45685
X17107 1878 1033 931 A[0] INV_X4 $T=66930 59800 1 180 $X=65865 $Y=59685
X17108 1512 338 931 A[0] INV_X4 $T=67500 51400 0 180 $X=66435 $Y=49885
X17109 1513 981 931 A[0] INV_X4 $T=67500 54200 0 180 $X=66435 $Y=52685
X17110 2337 1436 931 A[0] INV_X4 $T=67500 76600 1 0 $X=67385 $Y=75085
X17111 1517 1007 931 A[0] INV_X4 $T=68640 68200 0 180 $X=67575 $Y=66685
X17112 1522 1025 931 A[0] INV_X4 $T=69780 43000 0 180 $X=68715 $Y=41485
X17113 1535 164 931 A[0] INV_X4 $T=70160 48600 1 180 $X=69095 $Y=48485
X17114 1886 965 931 A[0] INV_X4 $T=70350 37400 1 180 $X=69285 $Y=37285
X17115 1521 1020 931 A[0] INV_X4 $T=69590 40200 1 0 $X=69475 $Y=38685
X17116 1524 506 931 A[0] INV_X4 $T=69590 54200 0 0 $X=69475 $Y=54085
X17117 1538 258 931 A[0] INV_X4 $T=72440 57000 1 0 $X=72325 $Y=55485
X17118 1902 991 931 A[0] INV_X4 $T=73960 37400 1 0 $X=73845 $Y=35885
X17119 1910 931 931 A[0] INV_X4 $T=74910 43000 1 180 $X=73845 $Y=42885
X17120 1563 1036 931 A[0] INV_X4 $T=78140 29000 1 180 $X=77075 $Y=28885
X17121 1562 428 931 A[0] INV_X4 $T=77380 31800 0 0 $X=77265 $Y=31685
X17122 1577 1012 931 A[0] INV_X4 $T=80040 34600 1 180 $X=78975 $Y=34485
X17123 931 1056 931 A[0] INV_X4 $T=80420 31800 0 180 $X=79355 $Y=30285
X17124 2361 983 931 A[0] INV_X4 $T=82320 31800 1 0 $X=82205 $Y=30285
X17141 936 A[0] 13 1600 931 931 NOR2_X1 $T=1380 45800 1 0 $X=1265 $Y=44285
X17142 1108 A[0] 937 1949 931 931 NOR2_X1 $T=2710 31800 0 0 $X=2595 $Y=31685
X17143 35 A[0] 1128 2368 931 931 NOR2_X1 $T=4230 45800 1 0 $X=4115 $Y=44285
X17144 48 A[0] 1151 2443 931 931 NOR2_X1 $T=5560 48600 1 0 $X=5445 $Y=47085
X17145 1600 A[0] 942 1175 931 931 NOR2_X1 $T=6890 45800 1 180 $X=6205 $Y=45685
X17146 1160 A[0] 1149 68 931 931 NOR2_X1 $T=8030 31800 1 0 $X=7915 $Y=30285
X17147 94 A[0] 91 1167 931 931 NOR2_X1 $T=8410 48600 1 0 $X=8295 $Y=47085
X17148 985 A[0] 1012 1974 931 931 NOR2_X1 $T=10120 3800 0 0 $X=10005 $Y=3685
X17149 1000 A[0] 965 2237 931 931 NOR2_X1 $T=10690 3800 0 0 $X=10575 $Y=3685
X17150 1000 A[0] 1020 2371 931 931 NOR2_X1 $T=11640 15000 0 180 $X=10955 $Y=13485
X17151 501 A[0] 1020 85 931 931 NOR2_X1 $T=11830 3800 1 180 $X=11145 $Y=3685
X17152 664 A[0] 1012 1646 931 931 NOR2_X1 $T=12210 15000 0 180 $X=11525 $Y=13485
X17153 664 A[0] 965 119 931 931 NOR2_X1 $T=11640 26200 1 0 $X=11525 $Y=24685
X17154 1667 A[0] 129 1189 931 931 NOR2_X1 $T=12400 51400 1 180 $X=11715 $Y=51285
X17155 985 A[0] 1020 2436 931 931 NOR2_X1 $T=12780 26200 0 180 $X=12095 $Y=24685
X17156 1033 A[0] 164 1195 931 931 NOR2_X1 $T=14680 17800 0 180 $X=13995 $Y=16285
X17157 931 A[0] 192 957 931 931 NOR2_X1 $T=15250 48600 0 0 $X=15135 $Y=48485
X17158 1663 A[0] 198 2372 931 931 NOR2_X1 $T=15250 62600 1 0 $X=15135 $Y=61085
X17159 501 A[0] 1012 191 931 931 NOR2_X1 $T=15820 6600 1 0 $X=15705 $Y=5085
X17160 664 A[0] 1020 2448 931 931 NOR2_X1 $T=15820 34600 1 0 $X=15705 $Y=33085
X17161 1668 A[0] 205 1193 931 931 NOR2_X1 $T=16580 62600 1 180 $X=15895 $Y=62485
X17162 1000 A[0] 1012 1209 931 931 NOR2_X1 $T=16580 3800 1 0 $X=16465 $Y=2285
X17163 958 A[0] 1995 185 931 931 NOR2_X1 $T=16770 57000 0 0 $X=16655 $Y=56885
X17164 1367 A[0] 2095 166 931 931 NOR2_X1 $T=17150 54200 1 0 $X=17035 $Y=52685
X17165 258 A[0] 1025 222 931 931 NOR2_X1 $T=17340 12200 1 0 $X=17225 $Y=10685
X17166 258 A[0] 164 233 931 931 NOR2_X1 $T=17910 6600 1 0 $X=17795 $Y=5085
X17167 501 A[0] 655 968 931 931 NOR2_X1 $T=17910 51400 1 0 $X=17795 $Y=49885
X17168 744 A[0] 338 1993 931 931 NOR2_X1 $T=18290 12200 0 0 $X=18175 $Y=12085
X17169 660 A[0] 788 1218 931 931 NOR2_X1 $T=18290 17800 0 0 $X=18175 $Y=17685
X17170 1033 A[0] 338 1997 931 931 NOR2_X1 $T=18290 51400 0 0 $X=18175 $Y=51285
X17171 1216 A[0] 1213 205 931 931 NOR2_X1 $T=18860 62600 0 180 $X=18175 $Y=61085
X17172 212 A[0] 1688 218 931 931 NOR2_X1 $T=18860 65400 1 180 $X=18175 $Y=65285
X17173 223 A[0] 1215 1995 931 931 NOR2_X1 $T=18670 54200 0 0 $X=18555 $Y=54085
X17174 1994 A[0] 1241 247 931 931 NOR2_X1 $T=18670 71000 0 0 $X=18555 $Y=70885
X17175 224 A[0] 221 201 931 931 NOR2_X1 $T=19620 57000 1 180 $X=18935 $Y=56885
X17176 1000 A[0] 164 1227 931 931 NOR2_X1 $T=19240 34600 1 0 $X=19125 $Y=33085
X17177 230 A[0] 1697 1999 931 931 NOR2_X1 $T=19430 71000 1 0 $X=19315 $Y=69485
X17178 985 A[0] 1025 2451 931 931 NOR2_X1 $T=19810 34600 1 0 $X=19695 $Y=33085
X17179 404 A[0] 655 2003 931 931 NOR2_X1 $T=20190 6600 0 0 $X=20075 $Y=6485
X17180 2251 A[0] 1231 250 931 931 NOR2_X1 $T=20190 82200 1 0 $X=20075 $Y=80685
X17181 931 A[0] 976 235 931 931 NOR2_X1 $T=20570 20600 1 0 $X=20455 $Y=19085
X17182 1220 A[0] 248 2376 931 931 NOR2_X1 $T=21330 73800 0 180 $X=20645 $Y=72285
X17183 1233 A[0] 1239 1242 931 931 NOR2_X1 $T=20760 79400 1 0 $X=20645 $Y=77885
X17184 258 A[0] 976 251 931 931 NOR2_X1 $T=20950 51400 1 0 $X=20835 $Y=49885
X17185 448 A[0] 1029 1243 931 931 NOR2_X1 $T=21900 3800 0 180 $X=21215 $Y=2285
X17186 931 A[0] 338 259 931 931 NOR2_X1 $T=21900 15000 0 180 $X=21215 $Y=13485
X17187 1231 A[0] 1242 1226 931 931 NOR2_X1 $T=21900 79400 0 180 $X=21215 $Y=77885
X17188 1024 A[0] 976 2248 931 931 NOR2_X1 $T=23040 15000 1 180 $X=22355 $Y=14885
X17189 1265 A[0] 1710 276 931 931 NOR2_X1 $T=22660 76600 1 0 $X=22545 $Y=75085
X17190 660 A[0] 983 2008 931 931 NOR2_X1 $T=23040 3800 1 0 $X=22925 $Y=2285
X17191 1080 A[0] 975 2015 931 931 NOR2_X1 $T=23610 15000 1 180 $X=22925 $Y=14885
X17192 428 A[0] 986 266 931 931 NOR2_X1 $T=23040 29000 1 0 $X=22925 $Y=27485
X17193 991 A[0] 980 1693 931 931 NOR2_X1 $T=23040 31800 1 0 $X=22925 $Y=30285
X17194 274 A[0] 2009 254 931 931 NOR2_X1 $T=23040 73800 0 0 $X=22925 $Y=73685
X17195 1080 A[0] 1015 1695 931 931 NOR2_X1 $T=23420 17800 0 0 $X=23305 $Y=17685
X17196 1036 A[0] 980 1255 931 931 NOR2_X1 $T=24180 31800 0 180 $X=23495 $Y=30285
X17197 1024 A[0] 1015 2253 931 931 NOR2_X1 $T=23800 20600 0 0 $X=23685 $Y=20485
X17198 501 A[0] 1009 1258 931 931 NOR2_X1 $T=23800 54200 0 0 $X=23685 $Y=54085
X17199 1000 A[0] 995 1257 931 931 NOR2_X1 $T=24750 51400 1 180 $X=24065 $Y=51285
X17200 1036 A[0] 1014 1263 931 931 NOR2_X1 $T=24370 29000 1 0 $X=24255 $Y=27485
X17201 258 A[0] 989 988 931 931 NOR2_X1 $T=24370 45800 0 0 $X=24255 $Y=45685
X17202 1036 A[0] 986 1267 931 931 NOR2_X1 $T=25130 23400 1 180 $X=24445 $Y=23285
X17203 991 A[0] 986 1254 931 931 NOR2_X1 $T=25130 26200 0 180 $X=24445 $Y=24685
X17204 301 A[0] 1271 248 931 931 NOR2_X1 $T=25320 73800 1 180 $X=24635 $Y=73685
X17205 664 A[0] 1014 1273 931 931 NOR2_X1 $T=25890 65400 0 180 $X=25205 $Y=63885
X17206 985 A[0] 1029 1275 931 2528 NOR2_X1 $T=26270 1000 1 180 $X=25585 $Y=885
X17207 428 A[0] 980 311 931 931 NOR2_X1 $T=25700 37400 1 0 $X=25585 $Y=35885
X17208 338 A[0] 1009 2025 931 931 NOR2_X1 $T=26270 54200 1 0 $X=26155 $Y=52685
X17209 973 A[0] 1015 1281 931 931 NOR2_X1 $T=27410 48600 1 180 $X=26725 $Y=48485
X17210 991 A[0] 981 1286 931 931 NOR2_X1 $T=27790 17800 0 180 $X=27105 $Y=16285
X17211 660 A[0] 1029 992 931 931 NOR2_X1 $T=27980 20600 0 180 $X=27295 $Y=19085
X17212 404 A[0] 976 2027 931 931 NOR2_X1 $T=28170 23400 0 180 $X=27485 $Y=21885
X17213 660 A[0] 981 2263 931 931 NOR2_X1 $T=28170 48600 0 180 $X=27485 $Y=47085
X17214 448 A[0] 788 2261 931 931 NOR2_X1 $T=28360 17800 0 180 $X=27675 $Y=16285
X17215 975 A[0] 1022 2433 931 931 NOR2_X1 $T=28360 54200 1 180 $X=27675 $Y=54085
X17216 1007 A[0] 1029 2031 931 931 NOR2_X1 $T=29120 29000 1 180 $X=28435 $Y=28885
X17217 1007 A[0] 997 305 931 931 NOR2_X1 $T=29500 9400 0 180 $X=28815 $Y=7885
X17218 744 A[0] 989 2264 931 931 NOR2_X1 $T=29690 23400 0 180 $X=29005 $Y=21885
X17219 744 A[0] 503 996 931 931 NOR2_X1 $T=29690 43000 1 180 $X=29005 $Y=42885
X17220 931 A[0] 975 1296 931 931 NOR2_X1 $T=29880 17800 0 180 $X=29195 $Y=16285
X17221 392 A[0] 983 1282 931 931 NOR2_X1 $T=30070 31800 0 180 $X=29385 $Y=30285
X17222 995 A[0] 1022 1288 931 931 NOR2_X1 $T=29500 71000 0 0 $X=29385 $Y=70885
X17223 392 A[0] 989 325 931 931 NOR2_X1 $T=30450 65400 1 180 $X=29765 $Y=65285
X17224 973 A[0] 1056 252 931 931 NOR2_X1 $T=30070 3800 0 0 $X=29955 $Y=3685
X17225 338 A[0] 1022 345 931 931 NOR2_X1 $T=30070 59800 0 0 $X=29955 $Y=59685
X17226 399 A[0] 997 327 931 931 NOR2_X1 $T=30260 23400 1 0 $X=30145 $Y=21885
X17227 448 A[0] 503 344 931 931 NOR2_X1 $T=30260 54200 0 0 $X=30145 $Y=54085
X17228 448 A[0] 980 331 931 931 NOR2_X1 $T=30450 68200 0 0 $X=30335 $Y=68085
X17229 1007 A[0] 1011 1302 931 931 NOR2_X1 $T=30640 9400 1 0 $X=30525 $Y=7885
X17230 428 A[0] 995 2037 931 931 NOR2_X1 $T=31210 37400 0 180 $X=30525 $Y=35885
X17231 319 A[0] 931 1304 931 931 NOR2_X1 $T=30640 73800 1 0 $X=30525 $Y=72285
X17232 931 A[0] 986 1292 931 931 NOR2_X1 $T=31400 43000 1 180 $X=30715 $Y=42885
X17233 506 A[0] 976 2267 931 931 NOR2_X1 $T=31210 45800 0 0 $X=31095 $Y=45685
X17234 399 A[0] 319 2384 931 931 NOR2_X1 $T=32350 76600 1 180 $X=31665 $Y=76485
X17235 991 A[0] 1009 2043 931 931 NOR2_X1 $T=32540 37400 0 180 $X=31855 $Y=35885
X17236 973 A[0] 1011 368 931 931 NOR2_X1 $T=32730 9400 0 180 $X=32045 $Y=7885
X17237 973 A[0] 997 334 931 931 NOR2_X1 $T=32350 3800 0 0 $X=32235 $Y=3685
X17238 392 A[0] 1011 1300 931 931 NOR2_X1 $T=32920 20600 0 180 $X=32235 $Y=19085
X17239 985 A[0] 164 2036 931 931 NOR2_X1 $T=32920 34600 0 180 $X=32235 $Y=33085
X17240 1080 A[0] 1014 1013 931 931 NOR2_X1 $T=32350 43000 1 0 $X=32235 $Y=41485
X17241 1007 A[0] 1015 2494 931 931 NOR2_X1 $T=32920 65400 0 180 $X=32235 $Y=63885
X17242 976 A[0] 392 2044 931 931 NOR2_X1 $T=32730 48600 0 0 $X=32615 $Y=48485
X17243 392 A[0] 1029 2053 931 931 NOR2_X1 $T=33110 26200 1 0 $X=32995 $Y=24685
X17244 660 A[0] 1056 2046 931 931 NOR2_X1 $T=34060 6600 0 180 $X=33375 $Y=5085
X17245 985 A[0] 1014 2049 931 931 NOR2_X1 $T=34440 51400 1 180 $X=33755 $Y=51285
X17246 976 A[0] 319 2050 931 931 NOR2_X1 $T=33870 68200 1 0 $X=33755 $Y=66685
X17247 448 A[0] 1020 2388 931 931 NOR2_X1 $T=34630 31800 0 180 $X=33945 $Y=30285
X17248 976 A[0] 399 1739 931 931 NOR2_X1 $T=34630 62600 1 180 $X=33945 $Y=62485
X17249 399 A[0] 1011 390 931 931 NOR2_X1 $T=35010 23400 0 180 $X=34325 $Y=21885
X17250 399 A[0] 995 2051 931 931 NOR2_X1 $T=34440 79400 1 0 $X=34325 $Y=77885
X17251 506 A[0] 989 371 931 931 NOR2_X1 $T=34630 48600 1 0 $X=34515 $Y=47085
X17252 664 A[0] 980 388 931 931 NOR2_X1 $T=34820 65400 0 0 $X=34705 $Y=65285
X17253 392 A[0] 1056 1319 931 931 NOR2_X1 $T=35010 23400 1 0 $X=34895 $Y=21885
X17254 655 A[0] 1022 2054 931 931 NOR2_X1 $T=35200 48600 0 0 $X=35085 $Y=48485
X17255 660 A[0] 1014 1740 931 931 NOR2_X1 $T=35200 73800 0 0 $X=35085 $Y=73685
X17256 319 A[0] 986 2062 931 931 NOR2_X1 $T=35390 76600 1 0 $X=35275 $Y=75085
X17257 404 A[0] 981 2460 931 931 NOR2_X1 $T=36530 48600 0 0 $X=36415 $Y=48485
X17258 985 A[0] 995 1327 931 931 NOR2_X1 $T=36530 62600 0 0 $X=36415 $Y=62485
X17259 399 A[0] 1015 2065 931 931 NOR2_X1 $T=37480 71000 0 180 $X=36795 $Y=69485
X17260 1025 A[0] 1009 393 931 931 NOR2_X1 $T=37670 48600 1 180 $X=36985 $Y=48485
X17261 338 A[0] 399 395 931 931 NOR2_X1 $T=37290 59800 1 0 $X=37175 $Y=58285
X17262 1022 A[0] 1014 1749 931 931 NOR2_X1 $T=38240 76600 0 180 $X=37555 $Y=75085
X17263 501 A[0] 788 402 931 931 NOR2_X1 $T=37860 3800 0 0 $X=37745 $Y=3685
X17264 660 A[0] 1020 1336 931 931 NOR2_X1 $T=38430 37400 0 180 $X=37745 $Y=35885
X17265 1022 A[0] 986 1353 931 931 NOR2_X1 $T=38240 76600 1 0 $X=38125 $Y=75085
X17266 1000 A[0] 338 401 931 931 NOR2_X1 $T=38620 48600 1 0 $X=38505 $Y=47085
X17267 399 A[0] 989 400 931 931 NOR2_X1 $T=38620 71000 1 0 $X=38505 $Y=69485
X17268 1080 A[0] 338 1756 931 931 NOR2_X1 $T=39570 12200 1 180 $X=38885 $Y=12085
X17269 744 A[0] 164 2285 931 931 NOR2_X1 $T=40140 6600 0 180 $X=39455 $Y=5085
X17270 1024 A[0] 338 427 931 931 NOR2_X1 $T=40140 20600 0 180 $X=39455 $Y=19085
X17271 1080 A[0] 655 1346 931 931 NOR2_X1 $T=40520 17800 0 180 $X=39835 $Y=16285
X17272 506 A[0] 1009 1023 931 931 NOR2_X1 $T=40520 51400 1 180 $X=39835 $Y=51285
X17273 1007 A[0] 981 1350 931 931 NOR2_X1 $T=40520 71000 0 180 $X=39835 $Y=69485
X17274 1033 A[0] 995 1348 931 931 NOR2_X1 $T=40710 54200 0 180 $X=40025 $Y=52685
X17275 501 A[0] 975 1352 931 931 NOR2_X1 $T=40900 48600 0 180 $X=40215 $Y=47085
X17276 392 A[0] 1015 1354 931 931 NOR2_X1 $T=41090 71000 0 180 $X=40405 $Y=69485
X17277 985 A[0] 986 1360 931 931 NOR2_X1 $T=40900 59800 0 0 $X=40785 $Y=59685
X17278 501 A[0] 1029 A[0] 931 931 NOR2_X1 $T=41280 20600 0 0 $X=41165 $Y=20485
X17279 985 A[0] 655 1364 931 931 NOR2_X1 $T=41850 45800 0 180 $X=41165 $Y=44285
X17280 392 A[0] 995 2080 931 931 NOR2_X1 $T=41850 79400 0 180 $X=41165 $Y=77885
X17281 1033 A[0] 976 1365 931 931 NOR2_X1 $T=42040 45800 1 180 $X=41355 $Y=45685
X17282 1000 A[0] 1014 2081 931 931 NOR2_X1 $T=42040 59800 1 180 $X=41355 $Y=59685
X17283 973 A[0] 503 417 931 931 NOR2_X1 $T=42230 68200 1 180 $X=41545 $Y=68085
X17284 660 A[0] 1015 1363 931 931 NOR2_X1 $T=42610 65400 0 180 $X=41925 $Y=63885
X17285 399 A[0] 788 1368 931 931 NOR2_X1 $T=42800 26200 0 180 $X=42115 $Y=24685
X17286 931 A[0] 1014 2082 931 931 NOR2_X1 $T=42800 29000 0 180 $X=42115 $Y=27485
X17287 664 A[0] 164 2075 931 931 NOR2_X1 $T=42800 43000 1 180 $X=42115 $Y=42885
X17288 660 A[0] 986 1361 931 931 NOR2_X1 $T=42800 68200 1 180 $X=42115 $Y=68085
X17289 1007 A[0] 319 1369 931 931 NOR2_X1 $T=42800 79400 1 180 $X=42115 $Y=79285
X17290 448 A[0] 1014 2294 931 931 NOR2_X1 $T=43370 68200 1 180 $X=42685 $Y=68085
X17291 1000 A[0] 983 2508 931 931 NOR2_X1 $T=43370 15000 1 0 $X=43255 $Y=13485
X17292 660 A[0] 989 447 931 931 NOR2_X1 $T=43940 62600 0 0 $X=43825 $Y=62485
X17293 664 A[0] 981 2303 931 931 NOR2_X1 $T=45080 62600 1 180 $X=44395 $Y=62485
X17294 501 A[0] 976 1782 931 931 NOR2_X1 $T=45270 23400 1 180 $X=44585 $Y=23285
X17295 980 A[0] 660 461 931 931 NOR2_X1 $T=45650 68200 1 0 $X=45535 $Y=66685
X17296 501 A[0] 983 463 931 931 NOR2_X1 $T=46600 3800 0 180 $X=45915 $Y=2285
X17297 258 A[0] 503 460 931 931 NOR2_X1 $T=46030 34600 1 0 $X=45915 $Y=33085
X17298 1080 A[0] 995 1387 931 931 NOR2_X1 $T=46790 37400 0 180 $X=46105 $Y=35885
X17299 1024 A[0] 1009 2102 931 931 NOR2_X1 $T=47170 37400 1 180 $X=46485 $Y=37285
X17300 399 A[0] 655 2306 931 931 NOR2_X1 $T=46790 48600 1 0 $X=46675 $Y=47085
X17301 931 A[0] 164 2103 931 931 NOR2_X1 $T=46790 51400 1 0 $X=46675 $Y=49885
X17302 1080 A[0] 164 1401 931 931 NOR2_X1 $T=47930 15000 0 0 $X=47815 $Y=14885
X17303 392 A[0] 1012 476 931 931 NOR2_X1 $T=48500 23400 1 180 $X=47815 $Y=23285
X17304 1024 A[0] 655 2113 931 931 NOR2_X1 $T=48310 12200 0 0 $X=48195 $Y=12085
X17305 501 A[0] 989 496 931 931 NOR2_X1 $T=48310 37400 1 0 $X=48195 $Y=35885
X17306 506 A[0] 788 1403 931 931 NOR2_X1 $T=49260 3800 0 180 $X=48575 $Y=2285
X17307 973 A[0] 976 2314 931 931 NOR2_X1 $T=49260 62600 0 0 $X=49145 $Y=62485
X17308 448 A[0] 319 1042 931 931 NOR2_X1 $T=50210 68200 1 180 $X=49525 $Y=68085
X17309 973 A[0] 1020 2311 931 931 NOR2_X1 $T=49830 23400 1 0 $X=49715 $Y=21885
X17310 1007 A[0] 1014 1410 931 931 NOR2_X1 $T=50400 76600 0 180 $X=49715 $Y=75085
X17311 1036 A[0] 976 1411 931 931 NOR2_X1 $T=50780 17800 0 180 $X=50095 $Y=16285
X17312 989 A[0] 1022 2474 931 931 NOR2_X1 $T=50400 65400 1 0 $X=50285 $Y=63885
X17313 664 A[0] 997 517 931 2528 NOR2_X1 $T=50780 1000 0 0 $X=50665 $Y=885
X17314 1048 A[0] 1052 1807 931 931 NOR2_X1 $T=50780 9400 0 0 $X=50665 $Y=9285
X17315 1007 A[0] 975 1412 931 931 NOR2_X1 $T=50780 59800 0 0 $X=50665 $Y=59685
X17316 1007 A[0] 980 529 931 931 NOR2_X1 $T=51920 79400 0 0 $X=51805 $Y=79285
X17317 744 A[0] 1020 1817 931 931 NOR2_X1 $T=52110 6600 0 0 $X=51995 $Y=6485
X17318 258 A[0] 1009 2312 931 931 NOR2_X1 $T=52680 57000 0 180 $X=51995 $Y=55485
X17319 319 A[0] 1015 1417 931 931 NOR2_X1 $T=52110 71000 1 0 $X=51995 $Y=69485
X17320 501 A[0] 1056 505 931 931 NOR2_X1 $T=52300 17800 0 0 $X=52185 $Y=17685
X17321 1080 A[0] 1025 1053 931 931 NOR2_X1 $T=52870 23400 0 180 $X=52185 $Y=21885
X17322 660 A[0] 164 1414 931 931 NOR2_X1 $T=52490 26200 1 0 $X=52375 $Y=24685
X17323 931 A[0] 1015 2120 931 931 NOR2_X1 $T=53060 65400 0 180 $X=52375 $Y=63885
X17324 399 A[0] 981 2124 931 931 NOR2_X1 $T=53630 68200 0 180 $X=52945 $Y=66685
X17325 985 A[0] 1011 1421 931 931 NOR2_X1 $T=53440 3800 1 0 $X=53325 $Y=2285
X17326 506 A[0] 1029 1058 931 931 NOR2_X1 $T=54200 20600 0 180 $X=53515 $Y=19085
X17327 399 A[0] 986 1423 931 931 NOR2_X1 $T=54960 79400 0 180 $X=54275 $Y=77885
X17328 1000 A[0] 976 2131 931 931 NOR2_X1 $T=54580 29000 1 0 $X=54465 $Y=27485
X17329 1022 A[0] 1020 2317 931 931 NOR2_X1 $T=54580 43000 1 0 $X=54465 $Y=41485
X17330 1000 A[0] 503 531 931 931 NOR2_X1 $T=54960 62600 1 0 $X=54845 $Y=61085
X17331 392 A[0] 1014 1430 931 931 NOR2_X1 $T=55530 79400 0 180 $X=54845 $Y=77885
X17332 258 A[0] 995 1446 931 931 NOR2_X1 $T=56290 54200 1 0 $X=56175 $Y=52685
X17333 448 A[0] 989 535 931 931 NOR2_X1 $T=56480 62600 0 0 $X=56365 $Y=62485
X17334 1009 A[0] 1020 2320 931 931 NOR2_X1 $T=57430 43000 0 180 $X=56745 $Y=41485
X17335 1000 A[0] 1011 1445 931 931 NOR2_X1 $T=57050 3800 1 0 $X=56935 $Y=2285
X17336 501 A[0] 986 2437 931 931 NOR2_X1 $T=57240 59800 0 0 $X=57125 $Y=59685
X17337 1007 A[0] 1020 2141 931 931 NOR2_X1 $T=57430 23400 0 0 $X=57315 $Y=23285
X17338 991 A[0] 338 1459 931 931 NOR2_X1 $T=58380 17800 1 0 $X=58265 $Y=16285
X17339 1036 A[0] 975 1842 931 931 NOR2_X1 $T=58380 17800 0 0 $X=58265 $Y=17685
X17340 1009 A[0] 983 566 931 931 NOR2_X1 $T=58380 26200 0 0 $X=58265 $Y=26085
X17341 985 A[0] 981 2146 931 931 NOR2_X1 $T=59140 62600 1 180 $X=58455 $Y=62485
X17342 664 A[0] 1015 1451 931 931 NOR2_X1 $T=59520 65400 0 180 $X=58835 $Y=63885
X17343 501 A[0] 1011 572 931 931 NOR2_X1 $T=59710 3800 0 180 $X=59025 $Y=2285
X17344 931 A[0] 1009 1458 931 931 NOR2_X1 $T=59710 43000 0 180 $X=59025 $Y=41485
X17345 1022 A[0] 788 2321 931 931 NOR2_X1 $T=59710 29000 0 0 $X=59595 $Y=28885
X17346 1033 A[0] 503 570 931 931 NOR2_X1 $T=59900 48600 1 0 $X=59785 $Y=47085
X17347 1033 A[0] 1056 2163 931 931 NOR2_X1 $T=60090 3800 0 0 $X=59975 $Y=3685
X17348 1022 A[0] 1012 607 931 931 NOR2_X1 $T=60660 37400 1 0 $X=60545 $Y=35885
X17349 931 A[0] 965 601 931 931 NOR2_X1 $T=61420 6600 0 0 $X=61305 $Y=6485
X17350 1000 A[0] 989 593 931 931 NOR2_X1 $T=61420 29000 1 0 $X=61305 $Y=27485
X17351 506 A[0] 983 1480 931 931 NOR2_X1 $T=62940 3800 0 180 $X=62255 $Y=2285
X17352 991 A[0] 655 1468 931 931 NOR2_X1 $T=62940 15000 0 180 $X=62255 $Y=13485
X17353 501 A[0] 997 2491 931 931 NOR2_X1 $T=63130 26200 0 0 $X=63015 $Y=26085
X17354 1036 A[0] 338 2164 931 931 NOR2_X1 $T=64080 15000 0 180 $X=63395 $Y=13485
X17355 392 A[0] 1020 1490 931 931 NOR2_X1 $T=64840 34600 1 180 $X=64155 $Y=34485
X17356 392 A[0] 1025 632 931 931 NOR2_X1 $T=64650 37400 0 0 $X=64535 $Y=37285
X17357 931 A[0] 1012 604 931 931 NOR2_X1 $T=65980 17800 0 180 $X=65295 $Y=16285
X17358 506 A[0] 1056 2326 931 931 NOR2_X1 $T=66170 26200 1 180 $X=65485 $Y=26085
X17359 258 A[0] 1029 640 931 931 NOR2_X1 $T=65980 3800 0 0 $X=65865 $Y=3685
X17360 448 A[0] 976 2412 931 931 NOR2_X1 $T=66550 54200 0 180 $X=65865 $Y=52685
X17361 448 A[0] 338 656 931 931 NOR2_X1 $T=66550 29000 0 0 $X=66435 $Y=28885
X17362 973 A[0] 164 1508 931 931 NOR2_X1 $T=67120 37400 0 180 $X=66435 $Y=35885
X17363 1024 A[0] 1020 1510 931 931 NOR2_X1 $T=67500 17800 0 180 $X=66815 $Y=16285
X17364 664 A[0] 976 2182 931 931 NOR2_X1 $T=67880 43000 0 180 $X=67195 $Y=41485
X17365 973 A[0] 655 661 931 931 NOR2_X1 $T=68260 37400 1 180 $X=67575 $Y=37285
X17366 931 A[0] 788 631 931 931 NOR2_X1 $T=68450 23400 1 180 $X=67765 $Y=23285
X17367 1007 A[0] 164 2187 931 931 NOR2_X1 $T=68830 37400 1 180 $X=68145 $Y=37285
X17368 1036 A[0] 164 2339 931 931 NOR2_X1 $T=69210 23400 1 0 $X=69095 $Y=21885
X17369 1532 A[0] 736 1888 931 931 NOR2_X1 $T=71110 73800 0 180 $X=70425 $Y=72285
X17370 258 A[0] 997 724 931 931 NOR2_X1 $T=72250 12200 1 180 $X=71565 $Y=12085
X17371 744 A[0] 983 2345 931 931 NOR2_X1 $T=72630 29000 0 0 $X=72515 $Y=28885
X17372 404 A[0] 997 784 931 931 NOR2_X1 $T=73200 3800 0 0 $X=73085 $Y=3685
X17373 737 A[0] reset 709 931 931 NOR2_X1 $T=74340 71000 0 180 $X=73655 $Y=69485
X17374 1080 A[0] 1029 1549 931 931 NOR2_X1 $T=75480 17800 0 180 $X=74795 $Y=16285
X17375 1024 A[0] 788 2489 931 931 NOR2_X1 $T=75670 15000 0 0 $X=75555 $Y=14885
X17376 744 A[0] 1011 2199 931 931 NOR2_X1 $T=76240 3800 1 0 $X=76125 $Y=2285
X17377 991 A[0] 1011 1560 931 931 NOR2_X1 $T=77760 26200 1 180 $X=77075 $Y=26085
X17378 1036 A[0] 1056 821 931 931 NOR2_X1 $T=78900 26200 0 180 $X=78215 $Y=24685
X17379 1024 A[0] 983 2204 931 931 NOR2_X1 $T=79280 3800 0 180 $X=78595 $Y=2285
X17380 1024 A[0] 1011 1568 931 931 NOR2_X1 $T=79470 26200 0 180 $X=78785 $Y=24685
X17381 1101 A[0] 840 1575 931 931 NOR2_X1 $T=80040 68200 0 0 $X=79925 $Y=68085
X17382 1024 A[0] 1056 1920 931 931 NOR2_X1 $T=80230 15000 0 0 $X=80115 $Y=14885
X17383 931 A[0] 1056 920 931 931 NOR2_X1 $T=80420 3800 0 0 $X=80305 $Y=3685
X17384 1024 A[0] 997 864 931 931 NOR2_X1 $T=81370 26200 1 0 $X=81255 $Y=24685
X17385 1080 A[0] 983 1591 931 931 NOR2_X1 $T=82320 3800 1 0 $X=82205 $Y=2285
X17386 1592 A[0] 1589 1582 931 931 NOR2_X1 $T=82890 15000 0 180 $X=82205 $Y=13485
X17387 931 A[0] 1139 1145 941 ICV_23 $T=5370 31800 1 0 $X=5255 $Y=30285
X17388 931 A[0] 1186 137 949 ICV_23 $T=11260 45800 1 0 $X=11145 $Y=44285
X17389 931 A[0] 501 965 168 ICV_23 $T=11450 3800 1 0 $X=11335 $Y=2285
X17390 931 A[0] 1033 1025 1192 ICV_23 $T=13160 6600 1 0 $X=13045 $Y=5085
X17391 931 A[0] 744 655 1998 ICV_23 $T=19050 9400 0 0 $X=18935 $Y=9285
X17392 931 A[0] 506 975 1225 ICV_23 $T=20190 51400 1 0 $X=20075 $Y=49885
X17393 931 A[0] 1080 989 2005 ICV_23 $T=22280 20600 0 0 $X=22165 $Y=20485
X17394 931 A[0] 660 503 284 ICV_23 $T=23230 65400 0 0 $X=23115 $Y=65285
X17395 931 A[0] 655 1009 1261 ICV_23 $T=23800 51400 1 0 $X=23685 $Y=49885
X17396 931 A[0] 931 503 2381 ICV_23 $T=24370 43000 0 0 $X=24255 $Y=42885
X17397 931 A[0] 1000 788 1287 ICV_23 $T=27410 3800 1 0 $X=27295 $Y=2285
X17398 931 A[0] 501 338 316 ICV_23 $T=28360 45800 0 0 $X=28245 $Y=45685
X17399 931 A[0] 1024 980 330 ICV_23 $T=28930 37400 1 0 $X=28815 $Y=35885
X17400 931 A[0] 399 983 361 ICV_23 $T=31210 26200 1 0 $X=31095 $Y=24685
X17401 931 A[0] 975 399 2386 ICV_23 $T=31970 48600 0 0 $X=31855 $Y=48485
X17402 931 A[0] 1009 997 391 ICV_23 $T=35010 26200 1 0 $X=34895 $Y=24685
X17403 931 A[0] 991 989 1018 ICV_23 $T=35200 17800 0 0 $X=35085 $Y=17685
X17404 931 A[0] 973 989 426 ICV_23 $T=39190 62600 0 0 $X=39075 $Y=62485
X17405 931 A[0] 404 503 409 ICV_23 $T=39380 29000 1 0 $X=39265 $Y=27485
X17406 931 A[0] 664 1011 A[0] ICV_23 $T=41090 15000 1 0 $X=40975 $Y=13485
X17407 931 A[0] 985 983 2084 ICV_23 $T=43180 3800 1 0 $X=43065 $Y=2285
X17408 931 A[0] 1022 1025 464 ICV_23 $T=44130 48600 0 0 $X=44015 $Y=48485
X17409 931 A[0] 660 1025 474 ICV_23 $T=47170 23400 0 0 $X=47055 $Y=23285
X17410 931 A[0] 501 503 519 ICV_23 $T=50590 40200 0 0 $X=50475 $Y=40085
X17411 931 A[0] 501 1014 1057 ICV_23 $T=52680 59800 0 0 $X=52565 $Y=59685
X17412 931 A[0] 392 965 1450 ICV_23 $T=55720 26200 1 0 $X=55605 $Y=24685
X17413 931 A[0] 1007 338 575 ICV_23 $T=58190 57000 1 0 $X=58075 $Y=55485
X17414 931 A[0] 1009 1029 1456 ICV_23 $T=58950 29000 0 0 $X=58835 $Y=28885
X17415 931 A[0] 404 1029 2428 ICV_23 $T=59140 23400 0 0 $X=59025 $Y=23285
X17416 931 A[0] 1080 965 1492 ICV_23 $T=66550 17800 0 0 $X=66435 $Y=17685
X17417 931 A[0] 448 975 2179 ICV_23 $T=66550 43000 1 0 $X=66435 $Y=41485
X17418 931 A[0] 428 1020 650 ICV_23 $T=67500 20600 0 0 $X=67385 $Y=20485
X17419 931 A[0] 1080 1012 1509 ICV_23 $T=70730 26200 1 0 $X=70615 $Y=24685
X17420 931 A[0] 991 1020 2418 ICV_23 $T=71110 17800 0 0 $X=70995 $Y=17685
X17421 931 A[0] 1036 1020 1091 ICV_23 $T=71110 20600 1 0 $X=70995 $Y=19085
X17422 931 A[0] 1080 788 1544 ICV_23 $T=73580 23400 0 0 $X=73465 $Y=23285
X17423 931 A[0] 404 983 2480 ICV_23 $T=74150 26200 1 0 $X=74035 $Y=24685
X17424 931 A[0] 991 1029 1576 ICV_23 $T=77380 15000 1 0 $X=77265 $Y=13485
X17425 931 A[0] 1024 981 1691 ICV_24 $T=22280 17800 1 0 $X=22165 $Y=16285
X17426 931 A[0] 982 1256 203 ICV_24 $T=23040 15000 1 0 $X=22925 $Y=13485
X17427 931 A[0] 338 931 362 ICV_24 $T=29500 48600 1 0 $X=29385 $Y=47085
X17428 931 A[0] 664 986 1311 ICV_24 $T=31590 51400 0 0 $X=31475 $Y=51285
X17429 931 A[0] 991 1015 1314 ICV_24 $T=32160 15000 0 0 $X=32045 $Y=14885
X17430 931 A[0] 931 1011 2270 ICV_24 $T=33300 23400 1 0 $X=33185 $Y=21885
X17431 931 A[0] 985 1015 1476 ICV_24 $T=60850 54200 0 0 $X=60735 $Y=54085
X17432 931 A[0] 399 1025 610 ICV_24 $T=62750 48600 1 0 $X=62635 $Y=47085
X17433 931 A[0] 1000 1015 1495 ICV_24 $T=63320 43000 0 0 $X=63205 $Y=42885
X17434 931 A[0] 1080 997 2212 ICV_24 $T=82320 26200 1 0 $X=82205 $Y=24685
X17435 1599 1941 7 931 A[0] 1950 HA_X1 $T=1000 54200 0 0 $X=885 $Y=54085
X17436 1109 1950 29 931 A[0] 47 HA_X1 $T=2330 57000 0 0 $X=2215 $Y=56885
X17437 933 1616 37 931 A[0] 38 HA_X1 $T=3280 31800 0 0 $X=3165 $Y=31685
X17438 1124 1621 44 931 A[0] 1148 HA_X1 $T=3850 76600 0 0 $X=3735 $Y=76485
X17439 1144 1134 43 931 A[0] 1139 HA_X1 $T=5940 23400 0 180 $X=3925 $Y=21885
X17440 1145 1605 1947 931 A[0] 1112 HA_X1 $T=4040 26200 0 0 $X=3925 $Y=26085
X17441 1604 47 49 931 A[0] 1141 HA_X1 $T=4230 57000 0 0 $X=4115 $Y=56885
X17442 1121 1133 52 931 A[0] 1621 HA_X1 $T=4230 76600 1 0 $X=4115 $Y=75085
X17443 1609 1138 55 931 A[0] 1961 HA_X1 $T=4610 59800 1 0 $X=4495 $Y=58285
X17444 1158 1140 932 931 A[0] 13 HA_X1 $T=4990 37400 1 0 $X=4875 $Y=35885
X17445 1129 1141 62 931 A[0] 1138 HA_X1 $T=4990 57000 1 0 $X=4875 $Y=55485
X17446 1613 1961 63 931 A[0] 1153 HA_X1 $T=4990 59800 0 0 $X=4875 $Y=59685
X17447 1120 1148 67 931 A[0] 1159 HA_X1 $T=5180 79400 1 0 $X=5065 $Y=77885
X17448 1607 1153 76 931 A[0] 1628 HA_X1 $T=5750 62600 1 0 $X=5635 $Y=61085
X17449 1620 1628 79 931 A[0] 1156 HA_X1 $T=8030 62600 1 180 $X=6015 $Y=62485
X17450 1608 1156 81 931 A[0] 944 HA_X1 $T=6130 65400 1 0 $X=6015 $Y=63885
X17451 1634 1648 83 931 A[0] 1133 HA_X1 $T=8220 73800 1 180 $X=6205 $Y=73685
X17452 1154 1159 92 931 A[0] 1969 HA_X1 $T=7080 79400 1 0 $X=6965 $Y=77885
X17453 1629 944 106 931 A[0] 1169 HA_X1 $T=8220 65400 0 0 $X=8105 $Y=65285
X17454 1631 1168 107 931 A[0] 1638 HA_X1 $T=8220 71000 1 0 $X=8105 $Y=69485
X17455 1165 1169 1627 931 A[0] 1972 HA_X1 $T=8410 68200 1 0 $X=8295 $Y=66685
X17456 1171 1969 114 931 A[0] 1181 HA_X1 $T=8980 79400 1 0 $X=8865 $Y=77885
X17457 1962 1972 116 931 A[0] 1168 HA_X1 $T=11260 68200 1 180 $X=9245 $Y=68085
X17458 99 1638 124 931 A[0] 1977 HA_X1 $T=9930 71000 0 0 $X=9815 $Y=70885
X17459 1642 1977 135 931 A[0] 1648 HA_X1 $T=10690 73800 0 0 $X=10575 $Y=73685
X17460 1643 1181 141 931 A[0] 1656 HA_X1 $T=10880 79400 1 0 $X=10765 $Y=77885
X17461 1197 952 182 931 A[0] 959 HA_X1 $T=14490 9400 0 0 $X=14375 $Y=9285
X17462 1199 959 210 931 A[0] 945 HA_X1 $T=16390 12200 0 0 $X=16275 $Y=12085
X17463 1256 1719 323 931 A[0] 2259 HA_X1 $T=27030 12200 0 0 $X=26915 $Y=12085
X17464 969 2033 335 931 A[0] 982 HA_X1 $T=28930 12200 0 0 $X=28815 $Y=12085
X17465 1048 1415 511 931 A[0] 2033 HA_X1 $T=51160 9400 1 0 $X=51045 $Y=7885
X17466 509 1834 520 931 A[0] 1415 HA_X1 $T=53440 9400 0 0 $X=53325 $Y=9285
X17467 512 1440 539 931 A[0] 1834 HA_X1 $T=58000 9400 0 180 $X=55985 $Y=7885
X17468 1847 2167 554 931 A[0] 1440 HA_X1 $T=59900 9400 0 180 $X=57885 $Y=7885
X17469 1452 2148 557 931 A[0] 591 HA_X1 $T=58190 76600 0 0 $X=58075 $Y=76485
X17470 1078 2410 612 931 A[0] 2167 HA_X1 $T=64270 6600 1 180 $X=62255 $Y=6485
X17471 649 1498 636 931 A[0] 2410 HA_X1 $T=66550 6600 0 180 $X=64535 $Y=5085
X17472 663 2184 682 931 A[0] 636 HA_X1 $T=68450 6600 1 0 $X=68335 $Y=5085
X17473 1889 776 690 931 A[0] 2336 HA_X1 $T=71110 76600 0 180 $X=69095 $Y=75085
X17474 1890 778 691 931 A[0] 1882 HA_X1 $T=71110 76600 1 180 $X=69095 $Y=76485
X17475 1525 2192 711 931 A[0] 682 HA_X1 $T=70540 6600 0 0 $X=70425 $Y=6485
X17476 1898 769 718 931 A[0] 1503 HA_X1 $T=73200 73800 1 180 $X=71185 $Y=73685
X17477 1088 786 756 931 A[0] 670 HA_X1 $T=73390 79400 1 180 $X=71375 $Y=79285
X17478 1900 1540 722 931 A[0] 2343 HA_X1 $T=73580 82200 0 180 $X=71565 $Y=80685
X17479 1906 787 734 931 A[0] 2330 HA_X1 $T=74720 79400 0 180 $X=72705 $Y=77885
X17480 1533 1547 753 931 A[0] 711 HA_X1 $T=74340 9400 1 0 $X=74225 $Y=7885
X17481 861 1566 797 931 A[0] 781 HA_X1 $T=79470 6600 0 180 $X=77455 $Y=5085
X17482 1559 1560 821 931 A[0] 1573 HA_X1 $T=78330 26200 0 0 $X=78215 $Y=26085
X17483 799 1573 864 931 A[0] 826 HA_X1 $T=80230 26200 0 0 $X=80115 $Y=26085
X17484 2427 2425 904 931 A[0] 903 HA_X1 $T=82320 12200 1 0 $X=82205 $Y=10685
X17485 1592 2216 905 931 A[0] 904 HA_X1 $T=82320 15000 0 0 $X=82205 $Y=14885
X17486 829 1594 906 931 A[0] 2216 HA_X1 $T=82320 20600 1 0 $X=82205 $Y=19085
X17498 931 A[0] 104 141 257 ICV_26 $T=20000 82200 0 0 $X=19885 $Y=82085
X17499 931 A[0] 1436 1465 582 ICV_26 $T=60090 65400 1 0 $X=59975 $Y=63885
X17500 931 A[0] 1436 1453 583 ICV_26 $T=60090 65400 0 0 $X=59975 $Y=65285
X17501 931 A[0] 883 547 585 ICV_26 $T=60090 73800 0 0 $X=59975 $Y=73685
X17502 931 A[0] 883 551 586 ICV_26 $T=60090 76600 0 0 $X=59975 $Y=76485
X17503 931 A[0] 1005 Res[25] 587 ICV_26 $T=60090 82200 0 0 $X=59975 $Y=82085
X17504 931 A[0] 1436 2352 848 ICV_26 $T=80040 29000 0 0 $X=79925 $Y=28885
X17505 931 A[0] 1436 1577 850 ICV_26 $T=80040 34600 0 0 $X=79925 $Y=34485
X17506 931 A[0] 883 827 851 ICV_26 $T=80040 40200 1 0 $X=79925 $Y=38685
X17507 931 A[0] 883 785 852 ICV_26 $T=80040 43000 1 0 $X=79925 $Y=41485
X17508 931 A[0] 883 755 854 ICV_26 $T=80040 54200 1 0 $X=79925 $Y=52685
X17509 931 A[0] 883 760 856 ICV_26 $T=80040 57000 0 0 $X=79925 $Y=56885
X17510 931 A[0] 883 721 857 ICV_26 $T=80040 62600 1 0 $X=79925 $Y=61085
X17511 931 A[0] 883 710 858 ICV_26 $T=80040 73800 1 0 $X=79925 $Y=72285
X17512 931 A[0] 883 690 859 ICV_26 $T=80040 76600 0 0 $X=79925 $Y=76485
X17513 931 A[0] 1436 2361 896 ICV_26 $T=82130 31800 0 0 $X=82015 $Y=31685
X17514 931 A[0] 883 907 897 ICV_26 $T=82130 37400 1 0 $X=82015 $Y=35885
X17515 931 A[0] 883 876 898 ICV_26 $T=82130 40200 0 0 $X=82015 $Y=40085
X17516 931 A[0] 883 1101 899 ICV_26 $T=82130 68200 0 0 $X=82015 $Y=68085
X17517 931 A[0] 883 691 901 ICV_26 $T=82130 79400 1 0 $X=82015 $Y=77885
X17518 931 A[0] 104 7 27 ICV_27 $T=1950 43000 0 0 $X=1835 $Y=42885
X17519 931 A[0] 104 49 28 ICV_27 $T=1950 54200 1 0 $X=1835 $Y=52685
X17520 931 A[0] 1005 Res[5] 31 ICV_27 $T=1950 68200 1 0 $X=1835 $Y=66685
X17521 931 A[0] 1436 1483 615 ICV_27 $T=61990 59800 0 0 $X=61875 $Y=59685
X17522 931 A[0] 1436 1482 617 ICV_27 $T=61990 68200 0 0 $X=61875 $Y=68085
X17523 931 A[0] 883 590 618 ICV_27 $T=61990 73800 1 0 $X=61875 $Y=72285
X17524 931 A[0] 883 886 909 ICV_27 $T=81940 43000 0 0 $X=81825 $Y=42885
X17525 931 A[0] 883 1540 913 ICV_27 $T=81940 82200 1 0 $X=81825 $Y=80685
X17537 1941 56 A[0] 1109 1105 934 931 AOI22_X1 $T=1950 59800 0 0 $X=1835 $Y=59685
X17538 29 56 A[0] 1604 1113 934 931 AOI22_X1 $T=2330 62600 1 0 $X=2215 $Y=61085
X17539 83 56 A[0] 1121 1954 934 931 AOI22_X1 $T=2900 73800 0 0 $X=2785 $Y=73685
X17540 44 56 A[0] 1120 1110 934 931 AOI22_X1 $T=3280 79400 0 0 $X=3165 $Y=79285
X17541 63 56 A[0] 1607 1115 934 931 AOI22_X1 $T=3470 71000 1 0 $X=3355 $Y=69485
X17542 49 56 A[0] 1129 2224 934 931 AOI22_X1 $T=4040 59800 0 0 $X=3925 $Y=59685
X17543 106 56 A[0] 1165 2222 934 931 AOI22_X1 $T=4230 68200 1 0 $X=4115 $Y=66685
X17544 79 56 A[0] 1608 1116 934 931 AOI22_X1 $T=5180 71000 1 180 $X=4115 $Y=70885
X17545 52 56 A[0] 1124 1130 934 931 AOI22_X1 $T=5180 79400 1 180 $X=4115 $Y=79285
X17546 62 56 A[0] 1609 1957 934 931 AOI22_X1 $T=4420 62600 1 0 $X=4305 $Y=61085
X17547 55 56 A[0] 1613 1618 934 931 AOI22_X1 $T=6130 65400 0 180 $X=5065 $Y=63885
X17548 76 56 A[0] 1620 1619 934 931 AOI22_X1 $T=5370 73800 0 0 $X=5255 $Y=73685
X17549 67 56 A[0] 1154 1623 934 931 AOI22_X1 $T=5940 79400 0 0 $X=5825 $Y=79285
X17550 1627 56 A[0] 1962 1152 934 931 AOI22_X1 $T=7460 68200 0 180 $X=6395 $Y=66685
X17551 116 56 A[0] 1631 82 934 931 AOI22_X1 $T=7270 71000 1 0 $X=7155 $Y=69485
X17552 81 56 A[0] 1629 2230 934 931 AOI22_X1 $T=7460 68200 1 0 $X=7345 $Y=66685
X17553 135 56 A[0] 1634 1166 934 931 AOI22_X1 $T=9170 73800 1 180 $X=8105 $Y=73685
X17554 107 56 A[0] 99 1635 934 931 AOI22_X1 $T=9550 73800 0 180 $X=8485 $Y=72285
X17555 92 56 A[0] 1171 1172 934 931 AOI22_X1 $T=8790 79400 0 0 $X=8675 $Y=79285
X17556 124 56 A[0] 1642 1639 934 931 AOI22_X1 $T=10690 76600 1 0 $X=10575 $Y=75085
X17557 114 56 A[0] 1643 1190 934 931 AOI22_X1 $T=10880 82200 1 0 $X=10765 $Y=80685
X17558 141 56 A[0] 1654 1201 934 931 AOI22_X1 $T=13350 79400 0 0 $X=13235 $Y=79285
X17559 1599 543 A[0] 157 704 7 931 AOI22_X1 $T=23230 68200 1 0 $X=23115 $Y=66685
X17560 982 1256 A[0] 967 971 969 931 AOI22_X1 $T=23990 12200 0 0 $X=23875 $Y=12085
X17561 290 2018 A[0] 1703 287 297 931 AOI22_X1 $T=24180 79400 1 0 $X=24065 $Y=77885
X17562 509 507 A[0] 1052 493 1048 931 AOI22_X1 $T=51160 12200 0 180 $X=50095 $Y=10685
X17563 512 1422 A[0] 504 1823 1847 931 AOI22_X1 $T=53440 12200 0 0 $X=53325 $Y=12085
X17564 663 1519 A[0] 1887 1884 1525 931 AOI22_X1 $T=69400 9400 1 0 $X=69285 $Y=7885
X17565 861 1923 A[0] 1904 686 1533 931 AOI22_X1 $T=73390 9400 1 0 $X=73275 $Y=7885
X17566 1560 1563 A[0] 1562 2203 1559 931 AOI22_X1 $T=78140 29000 1 0 $X=78025 $Y=27485
X17567 2427 1587 A[0] 1589 1584 1592 931 AOI22_X1 $T=81940 12200 0 0 $X=81825 $Y=12085
X17637 1598 1 1951 1659 A[0] 931 1117 2528 FA_X1 $T=1000 1000 0 0 $X=885 $Y=885
X17638 1953 1636 1114 1601 A[0] 931 1118 931 FA_X1 $T=1000 23400 1 0 $X=885 $Y=21885
X17639 37 2 1953 1968 A[0] 931 1605 931 FA_X1 $T=1000 26200 0 0 $X=885 $Y=26085
X17640 1956 41 1111 947 A[0] 931 2 931 FA_X1 $T=5370 26200 0 180 $X=2215 $Y=24685
X17641 932 22 1956 1664 A[0] 931 1616 931 FA_X1 $T=2330 29000 0 0 $X=2215 $Y=28885
X17642 34 33 1960 1641 A[0] 931 1140 931 FA_X1 $T=3090 37400 0 0 $X=2975 $Y=37285
X17643 1606 40 1150 1626 A[0] 931 87 931 FA_X1 $T=4040 9400 1 0 $X=3925 $Y=7885
X17644 43 87 1143 1655 A[0] 931 176 931 FA_X1 $T=8410 12200 0 180 $X=5255 $Y=10685
X17645 1960 88 2444 2228 A[0] 931 22 931 FA_X1 $T=8410 29000 1 180 $X=5255 $Y=28885
X17646 195 70 1161 1205 A[0] 931 2226 931 FA_X1 $T=5940 23400 1 0 $X=5825 $Y=21885
X17647 74 73 1967 1674 A[0] 931 1617 931 FA_X1 $T=6130 37400 0 0 $X=6015 $Y=37285
X17648 78 75 950 1210 A[0] 931 938 931 FA_X1 $T=6130 43000 1 0 $X=6015 $Y=41485
X17649 71 77 1966 961 A[0] 931 1636 931 FA_X1 $T=6320 26200 1 0 $X=6205 $Y=24685
X17650 1625 85 1192 2232 A[0] 931 1637 931 FA_X1 $T=7080 3800 0 0 $X=6965 $Y=3685
X17651 91 90 1622 1174 A[0] 931 948 931 FA_X1 $T=7460 43000 0 0 $X=7345 $Y=42885
X17652 1632 100 1637 1645 A[0] 931 1975 931 FA_X1 $T=8410 6600 0 0 $X=8295 $Y=6485
X17653 73 2370 1180 1704 A[0] 931 1641 931 FA_X1 $T=8410 34600 1 0 $X=8295 $Y=33085
X17654 1952 109 1974 2237 A[0] 931 1645 2528 FA_X1 $T=8980 1000 0 0 $X=8865 $Y=885
X17655 950 128 1173 2234 A[0] 931 1136 931 FA_X1 $T=12210 40200 0 180 $X=9055 $Y=38685
X17656 2225 145 1973 122 A[0] 931 101 931 FA_X1 $T=13350 12200 1 180 $X=10195 $Y=12085
X17657 1655 160 977 1958 A[0] 931 121 931 FA_X1 $T=14490 9400 1 180 $X=11335 $Y=9285
X17658 1951 168 1982 1194 A[0] 931 1647 2528 FA_X1 $T=15060 1000 1 180 $X=11905 $Y=885
X17659 137 146 1196 1787 A[0] 931 94 931 FA_X1 $T=12020 45800 1 0 $X=11905 $Y=44285
X17660 1976 170 1717 1978 A[0] 931 21 931 FA_X1 $T=15250 17800 1 180 $X=12095 $Y=17685
X17661 145 165 2374 1986 A[0] 931 2492 931 FA_X1 $T=13350 12200 0 0 $X=13235 $Y=12085
X17662 151 169 1699 1694 A[0] 931 961 931 FA_X1 $T=13730 26200 0 0 $X=13615 $Y=26085
X17663 1659 187 1672 1209 A[0] 931 1670 2528 FA_X1 $T=15060 1000 0 0 $X=14945 $Y=885
X17664 170 188 1684 2245 A[0] 931 17 931 FA_X1 $T=15250 17800 0 0 $X=15135 $Y=17685
X17665 955 189 978 216 A[0] 931 169 931 FA_X1 $T=15250 23400 0 0 $X=15135 $Y=23285
X17666 2242 217 1204 1765 A[0] 931 1164 931 FA_X1 $T=18480 40200 0 180 $X=15325 $Y=38685
X17667 1131 194 1647 1670 A[0] 931 268 931 FA_X1 $T=15820 3800 0 0 $X=15705 $Y=3685
X17668 1979 196 1669 1676 A[0] 931 184 931 FA_X1 $T=15820 31800 0 0 $X=15705 $Y=31685
X17669 1205 204 1218 2247 A[0] 931 59 931 FA_X1 $T=16200 20600 1 0 $X=16085 $Y=19085
X17670 189 207 1222 1223 A[0] 931 1126 931 FA_X1 $T=16580 23400 1 0 $X=16465 $Y=21885
X17671 1238 232 1234 1685 A[0] 931 2007 931 FA_X1 $T=18670 54200 1 0 $X=18555 $Y=52685
X17672 1170 234 1240 2492 A[0] 931 1689 931 FA_X1 $T=18860 9400 1 0 $X=18745 $Y=7885
X17673 165 259 2015 2248 A[0] 931 277 931 FA_X1 $T=21900 12200 1 180 $X=18745 $Y=12085
X17674 216 2013 1695 1691 A[0] 931 1684 931 FA_X1 $T=18860 17800 0 0 $X=18745 $Y=17685
X17675 1214 237 1235 2254 A[0] 931 142 931 FA_X1 $T=18860 29000 1 0 $X=18745 $Y=27485
X17676 149 260 1692 1677 A[0] 931 242 931 FA_X1 $T=21900 45800 0 180 $X=18745 $Y=44285
X17677 197 242 1690 1224 A[0] 931 2240 931 FA_X1 $T=18860 48600 0 0 $X=18745 $Y=48485
X17678 1244 968 1997 1225 A[0] 931 1224 931 FA_X1 $T=21900 51400 1 180 $X=18745 $Y=51285
X17679 256 243 1237 2007 A[0] 931 1686 931 FA_X1 $T=18860 57000 1 0 $X=18745 $Y=55485
X17680 1207 261 1707 2249 A[0] 931 221 931 FA_X1 $T=21900 59800 0 180 $X=18745 $Y=58285
X17681 212 245 2006 1687 A[0] 931 1213 931 FA_X1 $T=18860 62600 0 0 $X=18745 $Y=62485
X17682 1229 256 1246 1726 A[0] 931 245 931 FA_X1 $T=20190 68200 1 0 $X=20075 $Y=66685
X17683 1232 264 2378 2257 A[0] 931 1696 931 FA_X1 $T=20760 34600 1 0 $X=20645 $Y=33085
X17684 2006 267 1252 1770 A[0] 931 244 931 FA_X1 $T=21330 62600 1 0 $X=21215 $Y=61085
X17685 978 269 1254 1263 A[0] 931 188 931 FA_X1 $T=21520 26200 1 0 $X=21405 $Y=24685
X17686 234 277 1682 A[0] A[0] 931 1269 931 FA_X1 $T=22280 9400 0 0 $X=22165 $Y=9285
X17687 207 278 1260 1267 A[0] 931 1178 931 FA_X1 $T=22280 23400 1 0 $X=22165 $Y=21885
X17688 1250 988 1270 2021 A[0] 931 1711 931 FA_X1 $T=23040 48600 1 0 $X=22925 $Y=47085
X17689 1235 309 2016 2258 A[0] 931 1694 931 FA_X1 $T=26460 26200 1 180 $X=23305 $Y=26085
X17690 299 291 2454 2024 A[0] 931 120 931 FA_X1 $T=23420 34600 0 0 $X=23305 $Y=34485
X17691 303 293 992 2261 A[0] 931 1714 931 FA_X1 $T=23990 17800 0 0 $X=23875 $Y=17685
X17692 324 2453 2022 1289 A[0] 931 1277 931 FA_X1 $T=23990 65400 0 0 $X=23875 $Y=65285
X17693 1698 294 2023 1322 A[0] 931 1715 931 FA_X1 $T=23990 71000 0 0 $X=23875 $Y=70885
X17694 2023 296 1277 1721 A[0] 931 1246 931 FA_X1 $T=24180 68200 1 0 $X=24065 $Y=66685
X17695 2453 2025 2433 1723 A[0] 931 232 931 FA_X1 $T=24370 54200 0 0 $X=24255 $Y=54085
X17696 1701 1727 1278 1295 A[0] 931 1252 931 FA_X1 $T=24370 62600 1 0 $X=24255 $Y=61085
X17697 2233 298 1279 1725 A[0] 931 1253 931 FA_X1 $T=24560 15000 1 0 $X=24445 $Y=13485
X17698 1264 300 1280 2262 A[0] 931 994 931 FA_X1 $T=24560 40200 1 0 $X=24445 $Y=38685
X17699 282 2383 1281 2263 A[0] 931 1309 931 FA_X1 $T=24560 51400 1 0 $X=24445 $Y=49885
X17700 2380 303 1718 1294 A[0] 931 1717 931 FA_X1 $T=24750 20600 0 0 $X=24635 $Y=20485
X17701 1237 317 1301 2019 A[0] 931 1268 931 FA_X1 $T=27790 51400 1 180 $X=24635 $Y=51285
X17702 2254 308 2027 2264 A[0] 931 60 931 FA_X1 $T=25130 23400 0 0 $X=25015 $Y=23285
X17703 1721 321 2020 1305 A[0] 931 1278 931 FA_X1 $T=28360 62600 1 180 $X=25205 $Y=62485
X17704 290 314 1722 2266 A[0] 931 302 931 FA_X1 $T=25700 76600 0 0 $X=25585 $Y=76485
X17705 15 326 2457 2260 A[0] 931 1712 931 FA_X1 $T=29120 6600 0 180 $X=25965 $Y=5085
X17706 2454 322 1297 1720 A[0] 931 1003 931 FA_X1 $T=27220 26200 1 0 $X=27105 $Y=24685
X17707 1718 327 1300 2269 A[0] 931 16 931 FA_X1 $T=27980 20600 1 0 $X=27865 $Y=19085
X17708 1720 2461 2035 2270 A[0] 931 220 931 FA_X1 $T=28170 23400 0 0 $X=28055 $Y=23285
X17709 1280 330 2037 2043 A[0] 931 1729 931 FA_X1 $T=28360 37400 0 0 $X=28245 $Y=37285
X17710 314 336 1733 2274 A[0] 931 1732 931 FA_X1 $T=29500 79400 0 0 $X=29385 $Y=79285
X17711 453 339 994 2452 A[0] 931 348 931 FA_X1 $T=29690 40200 0 0 $X=29575 $Y=40085
X17712 2047 350 1306 1328 A[0] 931 1726 931 FA_X1 $T=33490 71000 0 180 $X=30335 $Y=69485
X17713 2048 351 1008 2456 A[0] 931 1006 931 FA_X1 $T=33680 29000 0 180 $X=30525 $Y=27485
X17714 1727 341 1738 2275 A[0] 931 283 931 FA_X1 $T=30640 59800 0 0 $X=30525 $Y=59685
X17715 1008 343 1310 2388 A[0] 931 1315 931 FA_X1 $T=31020 31800 1 0 $X=30905 $Y=30285
X17716 2039 344 1311 2049 A[0] 931 340 931 FA_X1 $T=31020 54200 1 0 $X=30905 $Y=52685
X17717 1305 345 2041 1739 A[0] 931 1738 931 FA_X1 $T=31020 62600 0 0 $X=30905 $Y=62485
X17718 1016 362 2386 2044 A[0] 931 1734 931 FA_X1 $T=34630 48600 0 180 $X=31475 $Y=47085
X17719 1308 353 1017 1737 A[0] 931 354 931 FA_X1 $T=32540 9400 0 0 $X=32425 $Y=9285
X17720 1733 355 2051 1744 A[0] 931 360 931 FA_X1 $T=32540 79400 0 0 $X=32425 $Y=79285
X17721 2055 368 2046 1316 A[0] 931 326 931 FA_X1 $T=35770 6600 1 180 $X=32615 $Y=6485
X17722 2298 358 1743 2050 A[0] 931 1322 931 FA_X1 $T=32730 71000 0 0 $X=32615 $Y=70885
X17723 292 359 1732 1730 A[0] 931 1741 931 FA_X1 $T=32730 82200 0 0 $X=32615 $Y=82085
X17724 359 360 1320 2283 A[0] 931 386 931 FA_X1 $T=32920 82200 1 0 $X=32805 $Y=80685
X17725 1019 376 1774 1735 A[0] 931 1737 931 FA_X1 $T=36910 12200 0 180 $X=33755 $Y=10685
X17726 1298 369 2061 1333 A[0] 931 350 931 FA_X1 $T=34440 68200 0 0 $X=34325 $Y=68085
X17727 2461 390 1319 2281 A[0] 931 1157 931 FA_X1 $T=37670 20600 1 180 $X=34515 $Y=20485
X17728 2457 372 1750 1355 A[0] 931 1747 2528 FA_X1 $T=35010 1000 0 0 $X=34895 $Y=885
X17729 1317 374 1018 2059 A[0] 931 1021 931 FA_X1 $T=35200 15000 0 0 $X=35085 $Y=14885
X17730 367 375 1332 1336 A[0] 931 380 931 FA_X1 $T=35200 34600 0 0 $X=35085 $Y=34485
X17731 347 2391 2394 1777 A[0] 931 1751 931 FA_X1 $T=35390 20600 1 0 $X=35275 $Y=19085
X17732 372 379 2067 2285 A[0] 931 1339 931 FA_X1 $T=35770 6600 0 0 $X=35655 $Y=6485
X17733 1333 400 1354 1350 A[0] 931 1351 931 FA_X1 $T=37480 68200 0 0 $X=37365 $Y=68085
X17734 1748 401 1352 1365 A[0] 931 1344 931 FA_X1 $T=37860 45800 0 0 $X=37745 $Y=45685
X17735 1750 402 2392 1349 A[0] 931 2495 2528 FA_X1 $T=38050 1000 0 0 $X=37935 $Y=885
X17736 2393 421 1763 1773 A[0] 931 438 931 FA_X1 $T=38810 12200 1 0 $X=38695 $Y=10685
X17737 2462 409 1028 2082 A[0] 931 2085 931 FA_X1 $T=38810 29000 0 0 $X=38695 $Y=28885
X17738 2074 412 1264 2488 A[0] 931 1765 931 FA_X1 $T=38810 37400 0 0 $X=38695 $Y=37285
X17739 2287 413 1357 1515 A[0] 931 1766 931 FA_X1 $T=38810 40200 1 0 $X=38695 $Y=38685
X17740 382 414 1358 1786 A[0] 931 1174 931 FA_X1 $T=38810 43000 1 0 $X=38695 $Y=41485
X17741 1342 415 2075 1364 A[0] 931 1767 931 FA_X1 $T=38810 43000 0 0 $X=38695 $Y=42885
X17742 172 1383 2076 429 A[0] 931 931 931 FA_X1 $T=38810 48600 0 0 $X=38695 $Y=48485
X17743 1338 423 1359 1831 A[0] 931 1768 931 FA_X1 $T=38810 57000 1 0 $X=38695 $Y=55485
X17744 406 A[0] 1372 2508 A[0] 931 2089 931 FA_X1 $T=41280 12200 0 0 $X=41165 $Y=12085
X17745 2295 435 1373 1782 A[0] 931 449 931 FA_X1 $T=41850 23400 1 0 $X=41735 $Y=21885
X17746 365 454 1768 1769 A[0] 931 1776 931 FA_X1 $T=45080 54200 1 180 $X=41925 $Y=54085
X17747 2293 440 2079 1784 A[0] 931 217 931 FA_X1 $T=42230 34600 1 0 $X=42115 $Y=33085
X17748 1030 441 2091 1406 A[0] 931 1375 931 FA_X1 $T=42230 34600 0 0 $X=42115 $Y=34485
X17749 2396 458 1031 2112 A[0] 931 418 931 FA_X1 $T=45270 71000 0 180 $X=42115 $Y=69485
X17750 1233 459 2466 2296 A[0] 931 274 931 FA_X1 $T=45270 76600 1 180 $X=42115 $Y=76485
X17751 2096 2098 2467 2472 A[0] 931 420 931 FA_X1 $T=45270 82200 1 180 $X=42115 $Y=82085
X17752 444 450 2094 1850 A[0] 931 1795 931 FA_X1 $T=42800 43000 0 0 $X=42685 $Y=42885
X17753 2467 451 2092 2304 A[0] 931 466 931 FA_X1 $T=42800 79400 0 0 $X=42685 $Y=79285
X17754 462 2395 1836 1402 A[0] 931 458 931 FA_X1 $T=46410 68200 1 180 $X=43255 $Y=68085
X17755 2302 462 1793 2305 A[0] 931 2105 931 FA_X1 $T=44510 73800 0 0 $X=44395 $Y=73685
X17756 2093 464 2103 2306 A[0] 931 486 931 FA_X1 $T=44890 48600 0 0 $X=44775 $Y=48485
X17757 1384 465 2104 2307 A[0] 931 1397 931 FA_X1 $T=45080 54200 0 0 $X=44965 $Y=54085
X17758 1797 480 1385 1815 A[0] 931 1791 931 FA_X1 $T=48120 62600 1 180 $X=44965 $Y=62485
X17759 2097 471 1809 1791 A[0] 931 1034 931 FA_X1 $T=45270 57000 0 0 $X=45155 $Y=56885
X17760 1793 472 1041 1042 A[0] 931 2112 931 FA_X1 $T=45270 71000 1 0 $X=45155 $Y=69485
X17761 2098 2136 1811 2116 A[0] 931 1379 931 FA_X1 $T=45270 82200 0 0 $X=45155 $Y=82085
X17762 1374 475 2109 1783 A[0] 931 484 931 FA_X1 $T=45650 9400 0 0 $X=45535 $Y=9285
X17763 1388 479 2115 1817 A[0] 931 495 931 FA_X1 $T=46600 6600 0 0 $X=46485 $Y=6485
X17764 2299 481 1046 1806 A[0] 931 500 931 FA_X1 $T=46980 17800 0 0 $X=46865 $Y=17685
X17765 2472 492 2107 2117 A[0] 931 1390 931 FA_X1 $T=50020 79400 1 180 $X=46865 $Y=79285
X17766 470 499 2114 2168 A[0] 931 1408 931 FA_X1 $T=50970 48600 1 180 $X=47815 $Y=48485
X17767 465 485 2118 1050 A[0] 931 1809 931 FA_X1 $T=48120 54200 0 0 $X=48005 $Y=54085
X17768 2307 486 1049 1457 A[0] 931 1810 931 FA_X1 $T=48310 51400 0 0 $X=48195 $Y=51285
X17769 1393 487 2119 2312 A[0] 931 1050 931 FA_X1 $T=48310 57000 0 0 $X=48195 $Y=56885
X17770 1391 500 1407 1804 A[0] 931 1801 931 FA_X1 $T=51540 15000 1 180 $X=48385 $Y=14885
X17771 1043 491 1047 1839 A[0] 931 1337 931 FA_X1 $T=48690 40200 1 0 $X=48575 $Y=38685
X17772 1405 495 1038 2505 A[0] 931 530 931 FA_X1 $T=49070 3800 0 0 $X=48955 $Y=3685
X17773 1406 496 2121 1409 A[0] 931 1816 931 FA_X1 $T=49070 34600 0 0 $X=48955 $Y=34485
X17774 446 1821 1825 1824 A[0] 931 2291 931 FA_X1 $T=50590 76600 0 0 $X=50475 $Y=76485
X17775 514 513 1424 1827 A[0] 931 491 931 FA_X1 $T=51730 34600 1 0 $X=51615 $Y=33085
X17776 1814 514 1466 1828 A[0] 931 450 931 FA_X1 $T=51730 40200 1 0 $X=51615 $Y=38685
X17777 2123 2485 1428 2319 A[0] 931 1829 931 FA_X1 $T=52680 45800 1 0 $X=52565 $Y=44285
X17778 2118 1837 2123 2316 A[0] 931 1419 931 FA_X1 $T=55910 45800 1 180 $X=52755 $Y=45685
X17779 1049 527 2126 2317 A[0] 931 2438 931 FA_X1 $T=56290 40200 1 180 $X=53135 $Y=40085
X17780 2136 529 2128 2127 A[0] 931 1821 931 FA_X1 $T=56290 82200 1 180 $X=53135 $Y=82085
X17781 1836 536 1429 1427 A[0] 931 1426 931 FA_X1 $T=57240 68200 1 180 $X=54085 $Y=68085
X17782 1831 532 592 2320 A[0] 931 537 931 FA_X1 $T=55720 54200 0 0 $X=55605 $Y=54085
X17783 1844 552 1830 1445 A[0] 931 1832 2528 FA_X1 $T=59140 1000 1 180 $X=55985 $Y=885
X17784 527 540 2145 555 A[0] 931 549 931 FA_X1 $T=56290 34600 0 0 $X=56175 $Y=34485
X17785 2104 553 2138 537 A[0] 931 471 931 FA_X1 $T=59330 57000 1 180 $X=56175 $Y=56885
X17786 2402 542 1832 1846 A[0] 931 561 931 FA_X1 $T=56480 15000 0 0 $X=56365 $Y=14885
X17787 1463 556 1446 2135 A[0] 931 1820 931 FA_X1 $T=59900 54200 0 180 $X=56745 $Y=52685
X17788 1434 2404 1479 2322 A[0] 931 1848 931 FA_X1 $T=57050 3800 0 0 $X=56935 $Y=3685
X17789 1066 2133 1450 2141 A[0] 931 1838 931 FA_X1 $T=60470 26200 0 180 $X=57315 $Y=24685
X17790 1833 1441 1459 1842 A[0] 931 546 931 FA_X1 $T=61990 17800 0 180 $X=58835 $Y=16285
X17791 2147 569 1448 1458 A[0] 931 1856 931 FA_X1 $T=58950 40200 0 0 $X=58835 $Y=40085
X17792 592 588 1461 2151 A[0] 931 1845 931 FA_X1 $T=61990 51400 0 180 $X=58835 $Y=49885
X17793 931 591 1906 2140 A[0] 931 1462 931 FA_X1 $T=61990 79400 1 180 $X=58835 $Y=79285
X17794 552 572 2163 1480 A[0] 931 1475 2528 FA_X1 $T=59140 1000 0 0 $X=59025 $Y=885
X17795 1464 574 1472 2154 A[0] 931 568 931 FA_X1 $T=59330 34600 1 0 $X=59215 $Y=33085
X17796 532 575 2165 594 A[0] 931 2506 931 FA_X1 $T=59330 57000 0 0 $X=59215 $Y=56885
X17797 2174 624 1880 1475 A[0] 931 581 2528 FA_X1 $T=65220 1000 1 180 $X=62065 $Y=885
X17798 1479 601 1487 2170 A[0] 931 624 931 FA_X1 $T=62370 3800 0 0 $X=62255 $Y=3685
X17799 560 602 1491 2327 A[0] 931 643 931 FA_X1 $T=62370 9400 1 0 $X=62255 $Y=7885
X17800 2327 2434 1076 1075 A[0] 931 603 931 FA_X1 $T=65410 12200 1 180 $X=62255 $Y=12085
X17801 1472 2172 1489 1490 A[0] 931 1870 931 FA_X1 $T=62370 34600 1 0 $X=62255 $Y=33085
X17802 1069 610 2173 1499 A[0] 931 1872 931 FA_X1 $T=62370 48600 0 0 $X=62255 $Y=48485
X17803 2411 637 1862 1868 A[0] 931 1861 931 FA_X1 $T=66170 15000 1 180 $X=63015 $Y=14885
X17804 1073 632 2187 661 A[0] 931 1514 931 FA_X1 $T=64650 40200 1 0 $X=64535 $Y=38685
X17805 574 638 1508 2180 A[0] 931 1081 931 FA_X1 $T=64840 34600 0 0 $X=64725 $Y=34485
X17806 2322 640 1507 2338 A[0] 931 1880 2528 FA_X1 $T=65220 1000 0 0 $X=65105 $Y=885
X17807 630 2413 1889 1882 A[0] 931 1526 931 FA_X1 $T=66170 76600 0 0 $X=66055 $Y=76485
X17808 637 1520 1527 2421 A[0] 931 2188 931 FA_X1 $T=66550 15000 0 0 $X=66435 $Y=14885
X17809 2185 679 1909 2341 A[0] 931 673 2528 FA_X1 $T=68260 1000 0 0 $X=68145 $Y=885
X17810 2434 701 2188 1881 A[0] 931 644 931 FA_X1 $T=71680 12200 1 180 $X=68525 $Y=12085
X17811 1076 692 1087 1876 A[0] 931 1894 931 FA_X1 $T=69590 26200 0 0 $X=69475 $Y=26085
X17812 628 713 1543 2345 A[0] 931 2507 931 FA_X1 $T=71110 29000 1 0 $X=70995 $Y=27485
X17813 701 714 2507 2479 A[0] 931 2191 931 FA_X1 $T=71300 20600 0 0 $X=71185 $Y=20485
X17814 2193 724 1090 1550 A[0] 931 1548 931 FA_X1 $T=72250 12200 0 0 $X=72135 $Y=12085
X17815 2421 763 1544 2419 A[0] 931 714 931 FA_X1 $T=76620 23400 0 180 $X=73465 $Y=21885
X17816 2479 742 2200 1091 A[0] 931 1556 931 FA_X1 $T=74150 17800 0 0 $X=74035 $Y=17685
X17817 2192 781 1546 1908 A[0] 931 1904 931 FA_X1 $T=77570 6600 0 180 $X=74415 $Y=5085
X17818 1546 770 1930 1917 A[0] 931 797 931 FA_X1 $T=75860 6600 0 0 $X=75745 $Y=6485
X17819 906 771 2481 1555 A[0] 931 820 931 FA_X1 $T=75860 20600 0 0 $X=75745 $Y=20485
X17820 1093 782 1095 2350 A[0] 931 1567 931 FA_X1 $T=76240 9400 1 0 $X=76125 $Y=7885
X17821 862 804 1576 1558 A[0] 931 905 931 FA_X1 $T=78140 15000 1 0 $X=78025 $Y=13485
X17822 1917 824 1561 2424 A[0] 931 2213 931 FA_X1 $T=78900 6600 0 0 $X=78785 $Y=6485
X17823 1930 862 2207 2202 A[0] 931 902 931 FA_X1 $T=81940 12200 1 180 $X=78785 $Y=12085
X17824 2423 826 2212 1568 A[0] 931 1594 931 FA_X1 $T=78900 23400 0 0 $X=78785 $Y=23285
X17825 1566 902 2213 1924 A[0] 931 1587 931 FA_X1 $T=84030 3800 1 180 $X=80875 $Y=3685
X17826 753 903 1567 1926 A[0] 931 1923 931 FA_X1 $T=84030 9400 0 180 $X=80875 $Y=7885
X17827 1939 920 1591 1581 A[0] 931 1926 2528 FA_X1 $T=84410 1000 1 180 $X=81255 $Y=885
X17843 573 A[0] 590 547 551 1852 931 NOR4_X1 $T=60090 71000 0 0 $X=59975 $Y=70885
X17844 579 A[0] 625 635 629 1874 931 NOR4_X1 $T=65980 65400 1 180 $X=64915 $Y=65285
X17845 706 A[0] 687 598 708 1891 931 NOR4_X1 $T=70730 62600 0 0 $X=70615 $Y=62485
X17846 681 A[0] 683 717 716 1892 931 NOR4_X1 $T=70920 45800 1 0 $X=70805 $Y=44285
X17847 672 A[0] 665 703 654 1897 931 NOR4_X1 $T=72060 54200 0 0 $X=71945 $Y=54085
X17848 700 A[0] 695 728 694 1541 931 NOR4_X1 $T=73580 62600 0 180 $X=72515 $Y=61085
X17849 699 A[0] 684 719 732 1893 931 NOR4_X1 $T=73960 48600 0 180 $X=72895 $Y=47085
X17850 738 A[0] 715 785 774 1899 931 NOR4_X1 $T=75480 40200 0 0 $X=75365 $Y=40085
X17851 693 A[0] 721 761 760 1092 931 NOR4_X1 $T=76620 59800 0 180 $X=75555 $Y=58285
X17852 1912 A[0] 1903 739 reset 1913 931 NOR4_X1 $T=75860 68200 1 0 $X=75745 $Y=66685
X17853 907 A[0] 844 886 876 1895 931 NOR4_X1 $T=82130 37400 0 180 $X=81065 $Y=35885
X17854 1158 38 2487 64 931 A[0] AOI21_X1 $T=4040 34600 0 0 $X=3925 $Y=34485
X17855 1162 53 1107 941 931 A[0] AOI21_X1 $T=5940 31800 1 180 $X=5065 $Y=31685
X17856 1132 24 2445 942 931 A[0] AOI21_X1 $T=6510 45800 1 0 $X=6395 $Y=44285
X17857 94 91 2227 1167 931 A[0] AOI21_X1 $T=7650 48600 1 0 $X=7535 $Y=47085
X17858 1667 129 1176 1189 931 A[0] AOI21_X1 $T=11070 51400 0 0 $X=10955 $Y=51285
X17859 1644 133 2239 949 931 A[0] AOI21_X1 $T=12210 45800 1 180 $X=11335 $Y=45685
X17860 155 148 1185 102 931 A[0] AOI21_X1 $T=13350 34600 0 180 $X=12475 $Y=33085
X17861 1652 152 954 201 931 A[0] AOI21_X1 $T=13540 59800 1 180 $X=12665 $Y=59685
X17862 1219 154 1651 1995 931 A[0] AOI21_X1 $T=13730 57000 1 180 $X=12855 $Y=56885
X17863 2373 199 1212 1999 931 A[0] AOI21_X1 $T=16010 71000 1 0 $X=15895 $Y=69485
X17864 206 208 2244 218 931 A[0] AOI21_X1 $T=16770 68200 0 0 $X=16655 $Y=68085
X17865 221 224 2449 201 931 A[0] AOI21_X1 $T=18100 59800 1 0 $X=17985 $Y=58285
X17866 2002 227 231 254 931 A[0] AOI21_X1 $T=18290 76600 1 0 $X=18175 $Y=75085
X17867 1697 230 2450 1999 931 A[0] AOI21_X1 $T=18670 71000 1 0 $X=18555 $Y=69485
X17868 1703 290 2379 1251 931 A[0] AOI21_X1 $T=24180 79400 0 180 $X=23305 $Y=77885
X17869 2018 297 2026 2379 931 A[0] AOI21_X1 $T=24370 79400 0 0 $X=24255 $Y=79285
X17870 1078 643 648 1879 931 A[0] AOI21_X1 $T=67310 9400 1 0 $X=67195 $Y=7885
X17871 1934 674 2337 reset 931 A[0] AOI21_X1 $T=68450 76600 1 0 $X=68335 $Y=75085
X17872 2342 709 1433 1913 931 A[0] AOI21_X1 $T=70920 68200 0 0 $X=70805 $Y=68085
X17873 829 869 874 2435 931 A[0] AOI21_X1 $T=81940 20600 1 180 $X=81065 $Y=20485
X17874 936 13 1602 24 931 A[0] OAI21_X1 $T=2330 45800 1 0 $X=2215 $Y=44285
X17875 1123 35 1122 1137 931 A[0] OAI21_X1 $T=3470 45800 0 0 $X=3355 $Y=45685
X17876 935 48 1612 940 931 A[0] OAI21_X1 $T=4800 48600 1 0 $X=4685 $Y=47085
X17877 1943 64 1146 1624 931 A[0] OAI21_X1 $T=5750 34600 0 0 $X=5635 $Y=34485
X17878 1155 68 1624 939 931 A[0] OAI21_X1 $T=6890 34600 0 180 $X=6015 $Y=33085
X17879 953 68 1162 1163 931 A[0] OAI21_X1 $T=8030 31800 0 0 $X=7915 $Y=31685
X17880 946 102 2231 1177 931 A[0] OAI21_X1 $T=9550 34600 1 180 $X=8675 $Y=34485
X17881 2235 111 1971 133 931 A[0] OAI21_X1 $T=10310 45800 1 180 $X=9435 $Y=45685
X17882 1185 136 1644 1175 931 A[0] OAI21_X1 $T=11450 43000 1 0 $X=11335 $Y=41485
X17883 1186 137 115 1187 931 A[0] OAI21_X1 $T=11450 48600 1 0 $X=11335 $Y=47085
X17884 129 138 2500 1188 931 A[0] OAI21_X1 $T=11450 51400 1 0 $X=11335 $Y=49885
X17885 1189 143 144 1191 931 A[0] OAI21_X1 $T=12020 54200 1 0 $X=11905 $Y=52685
X17886 1202 172 2447 1191 931 A[0] OAI21_X1 $T=14110 51400 0 0 $X=13995 $Y=51285
X17887 1202 172 143 1188 931 A[0] OAI21_X1 $T=14870 51400 0 0 $X=14755 $Y=51285
X17888 1688 212 1666 206 931 A[0] OAI21_X1 $T=16960 65400 0 0 $X=16845 $Y=65285
X17889 1215 223 1673 1219 931 A[0] OAI21_X1 $T=18100 57000 1 0 $X=17985 $Y=55485
X17890 1221 231 2432 1226 931 A[0] OAI21_X1 $T=18670 79400 1 0 $X=18555 $Y=77885
X17891 2009 274 1228 2002 931 A[0] OAI21_X1 $T=22280 73800 0 0 $X=22165 $Y=73685
X17892 302 292 1266 1226 931 A[0] OAI21_X1 $T=24940 76600 1 180 $X=24065 $Y=76485
X17893 1285 319 307 993 931 A[0] OAI21_X1 $T=27790 79400 1 180 $X=26915 $Y=79285
X17894 1285 319 320 2030 931 A[0] OAI21_X1 $T=28550 79400 1 180 $X=27675 $Y=79285
X17895 1431 528 544 1433 931 A[0] OAI21_X1 $T=55150 82200 1 0 $X=55035 $Y=80685
X17896 2149 528 558 1433 931 A[0] OAI21_X1 $T=58570 82200 1 0 $X=58455 $Y=80685
X17897 1470 528 587 1433 931 A[0] OAI21_X1 $T=61610 82200 0 180 $X=60735 $Y=80685
X17898 1082 528 619 1433 931 A[0] OAI21_X1 $T=66170 76600 1 180 $X=65295 $Y=76485
X17899 1501 528 642 1433 931 A[0] OAI21_X1 $T=65980 82200 1 0 $X=65865 $Y=80685
X17900 1518 528 662 1433 931 A[0] OAI21_X1 $T=68830 73800 1 0 $X=68715 $Y=72285
X17901 1523 528 671 1433 931 A[0] OAI21_X1 $T=69970 82200 0 180 $X=69095 $Y=80685
X17902 1531 528 688 1433 931 A[0] OAI21_X1 $T=71680 82200 0 180 $X=70805 $Y=80685
X17903 1545 730 766 1542 931 A[0] OAI21_X1 $T=73770 68200 0 180 $X=72895 $Y=66685
X17904 1582 874 868 1584 931 A[0] OAI21_X1 $T=81180 15000 1 0 $X=81065 $Y=13485
X17905 931 A[0] 1 233 2003 1993 194 ICV_35 $T=18860 3800 0 0 $X=18745 $Y=3685
X17906 931 A[0] 1676 238 1696 263 1198 ICV_35 $T=18860 31800 0 0 $X=18745 $Y=31685
X17907 931 A[0] 270 239 1232 2255 1992 ICV_35 $T=18860 37400 1 0 $X=18745 $Y=35885
X17908 931 A[0] 171 240 348 2056 1173 ICV_35 $T=18860 40200 0 0 $X=18745 $Y=40085
X17909 931 A[0] 1216 244 262 1686 177 ICV_35 $T=18860 59800 0 0 $X=18745 $Y=59685
X17910 931 A[0] 2070 406 1032 2292 1761 ICV_35 $T=38810 6600 0 0 $X=38695 $Y=6485
X17911 931 A[0] 1340 1021 2073 1339 1762 ICV_35 $T=38810 9400 0 0 $X=38695 $Y=9285
X17912 931 A[0] 2300 408 1026 1368 363 ICV_35 $T=38810 26200 1 0 $X=38695 $Y=24685
X17913 931 A[0] 2009 425 1362 2110 301 ICV_35 $T=38810 76600 1 0 $X=38695 $Y=75085
X17914 931 A[0] 1437 561 1849 2406 554 ICV_35 $T=58950 12200 0 0 $X=58835 $Y=12085
X17915 931 A[0] 2404 562 1468 2164 1853 ICV_35 $T=58950 15000 1 0 $X=58835 $Y=13485
X17916 931 A[0] 1065 563 2407 2323 1473 ICV_35 $T=58950 17800 0 0 $X=58835 $Y=17685
X17917 931 A[0] 564 565 2428 1471 606 ICV_35 $T=58950 23400 1 0 $X=58835 $Y=21885
X17918 931 A[0] 2476 566 2160 2324 2166 ICV_35 $T=58950 26200 0 0 $X=58835 $Y=26085
X17919 931 A[0] 482 568 1855 1856 1474 ICV_35 $T=58950 37400 0 0 $X=58835 $Y=37285
X17920 931 A[0] 1457 571 2162 1069 502 ICV_35 $T=58950 51400 0 0 $X=58835 $Y=51285
X17921 931 A[0] 2425 875 2423 2365 1589 ICV_35 $T=80990 17800 0 0 $X=80875 $Y=17685
X17957 1105 931 A[0] 25 INV_X1 $T=1570 62600 1 0 $X=1455 $Y=61085
X17958 1943 931 A[0] 1108 INV_X1 $T=1760 31800 0 0 $X=1645 $Y=31685
X17959 1954 931 A[0] 32 INV_X1 $T=2330 76600 0 0 $X=2215 $Y=76485
X17960 1110 931 A[0] 45 INV_X1 $T=2710 82200 1 0 $X=2595 $Y=80685
X17961 1113 931 A[0] 8 INV_X1 $T=3280 65400 0 180 $X=2785 $Y=63885
X17962 2222 931 A[0] 3 INV_X1 $T=3280 68200 1 180 $X=2785 $Y=68085
X17963 1115 931 A[0] 26 INV_X1 $T=3470 71000 0 180 $X=2975 $Y=69485
X17964 1116 931 A[0] 4 INV_X1 $T=3470 73800 0 180 $X=2975 $Y=72285
X17965 1619 931 A[0] 9 INV_X1 $T=3850 76600 1 180 $X=3355 $Y=76485
X17966 1618 931 A[0] 31 INV_X1 $T=4230 65400 1 180 $X=3735 $Y=65285
X17967 2224 931 A[0] 30 INV_X1 $T=4610 59800 0 180 $X=4115 $Y=58285
X17968 1122 931 A[0] 935 INV_X1 $T=4420 48600 1 0 $X=4305 $Y=47085
X17969 1130 931 A[0] 72 INV_X1 $T=4610 82200 1 0 $X=4495 $Y=80685
X17970 1132 931 A[0] 35 INV_X1 $T=5180 45800 0 180 $X=4685 $Y=44285
X17971 1128 931 A[0] 1137 INV_X1 $T=5180 45800 1 0 $X=5065 $Y=44285
X17972 1957 931 A[0] 50 INV_X1 $T=5750 62600 0 180 $X=5255 $Y=61085
X17973 1144 931 A[0] 1149 INV_X1 $T=5940 26200 1 0 $X=5825 $Y=24685
X17974 1151 931 A[0] 940 INV_X1 $T=6510 48600 0 180 $X=6015 $Y=47085
X17975 1152 931 A[0] 51 INV_X1 $T=6510 68200 0 180 $X=6015 $Y=66685
X17976 1635 931 A[0] 39 INV_X1 $T=6700 71000 1 180 $X=6205 $Y=70885
X17977 53 931 A[0] 1155 INV_X1 $T=6890 31800 1 180 $X=6395 $Y=31685
X17978 82 931 A[0] 66 INV_X1 $T=7270 71000 0 180 $X=6775 $Y=69485
X17979 1623 931 A[0] 84 INV_X1 $T=6890 79400 0 0 $X=6775 $Y=79285
X17980 2230 931 A[0] 69 INV_X1 $T=8030 71000 1 180 $X=7535 $Y=70885
X17981 1166 931 A[0] 98 INV_X1 $T=8600 76600 1 0 $X=8485 $Y=75085
X17982 1167 931 A[0] 61 INV_X1 $T=8980 48600 1 0 $X=8865 $Y=47085
X17983 945 931 A[0] 1160 INV_X1 $T=9170 20600 1 0 $X=9055 $Y=19085
X17984 1172 931 A[0] 108 INV_X1 $T=9740 82200 0 180 $X=9245 $Y=80685
X17985 953 931 A[0] 946 INV_X1 $T=9930 34600 1 180 $X=9435 $Y=34485
X17986 1175 931 A[0] 111 INV_X1 $T=10500 45800 0 180 $X=10005 $Y=44285
X17987 1176 931 A[0] 97 INV_X1 $T=10500 54200 0 180 $X=10005 $Y=52685
X17988 1177 931 A[0] 136 INV_X1 $T=10500 37400 1 0 $X=10385 $Y=35885
X17989 1183 931 A[0] 129 INV_X1 $T=11070 51400 1 0 $X=10955 $Y=49885
X17990 1639 931 A[0] 140 INV_X1 $T=11640 76600 1 0 $X=11525 $Y=75085
X17991 1190 931 A[0] 131 INV_X1 $T=12210 82200 0 180 $X=11715 $Y=80685
X17992 1187 931 A[0] 1182 INV_X1 $T=12970 48600 1 0 $X=12855 $Y=47085
X17993 543 931 A[0] 157 INV_X1 $T=13160 71000 0 0 $X=13045 $Y=70885
X17994 1651 931 A[0] 1652 INV_X1 $T=13920 59800 1 180 $X=13425 $Y=59685
X17995 1197 931 A[0] 1657 INV_X1 $T=14490 12200 1 0 $X=14375 $Y=10685
X17996 1200 931 A[0] 154 INV_X1 $T=14870 57000 0 180 $X=14375 $Y=55485
X17997 1201 931 A[0] 202 INV_X1 $T=14680 82200 1 0 $X=14565 $Y=80685
X17998 1662 931 A[0] 1663 INV_X1 $T=16010 62600 1 180 $X=15515 $Y=62485
X17999 957 931 A[0] 1188 INV_X1 $T=16200 51400 0 180 $X=15705 $Y=49885
X18000 2244 931 A[0] 2373 INV_X1 $T=16770 68200 1 180 $X=16275 $Y=68085
X18001 2095 931 A[0] 960 INV_X1 $T=16960 54200 1 180 $X=16465 $Y=54085
X18002 211 931 A[0] 1668 INV_X1 $T=16960 62600 1 180 $X=16465 $Y=62485
X18003 1367 931 A[0] 1989 INV_X1 $T=17340 54200 1 180 $X=16845 $Y=54085
X18004 1220 931 A[0] 1990 INV_X1 $T=18860 73800 0 180 $X=18365 $Y=72285
X18005 971 931 A[0] 175 INV_X1 $T=19050 15000 1 0 $X=18935 $Y=13485
X18006 2040 931 A[0] 2251 INV_X1 $T=19620 82200 0 0 $X=19505 $Y=82085
X18007 2252 931 A[0] 1221 INV_X1 $T=20570 76600 1 180 $X=20075 $Y=76485
X18008 2000 931 A[0] 286 INV_X1 $T=22280 76600 1 0 $X=22165 $Y=75085
X18009 1710 931 A[0] 275 INV_X1 $T=23610 76600 0 180 $X=23115 $Y=75085
X18010 1703 931 A[0] 2018 INV_X1 $T=23990 79400 0 0 $X=23875 $Y=79285
X18011 2259 931 A[0] 1661 INV_X1 $T=24180 15000 1 0 $X=24065 $Y=13485
X18012 290 931 A[0] 297 INV_X1 $T=26650 79400 0 180 $X=26155 $Y=77885
X18013 1283 931 A[0] 1285 INV_X1 $T=27030 79400 1 0 $X=26915 $Y=77885
X18014 reset 931 A[0] 93 INV_X1 $T=44130 65400 0 0 $X=44015 $Y=65285
X18015 1416 931 A[0] 1413 INV_X1 $T=51920 12200 0 0 $X=51805 $Y=12085
X18016 1835 931 A[0] 524 INV_X1 $T=54390 65400 0 0 $X=54275 $Y=65285
X18017 1452 931 A[0] 1431 INV_X1 $T=55720 79400 1 180 $X=55225 $Y=79285
X18018 1462 931 A[0] 2149 INV_X1 $T=59710 82200 0 180 $X=59215 $Y=80685
X18019 1478 931 A[0] 1470 INV_X1 $T=62370 82200 0 180 $X=61875 $Y=80685
X18020 1511 931 A[0] 1501 INV_X1 $T=67120 79400 1 0 $X=67005 $Y=77885
X18021 2183 931 A[0] 1082 INV_X1 $T=67500 73800 0 0 $X=67385 $Y=73685
X18022 enable 931 A[0] 1084 INV_X1 $T=69590 68200 1 180 $X=69095 $Y=68085
X18023 1526 931 A[0] 1523 INV_X1 $T=70350 82200 0 180 $X=69855 $Y=80685
X18024 1528 931 A[0] 1531 INV_X1 $T=70540 82200 1 0 $X=70425 $Y=80685
X18025 1530 931 A[0] 730 INV_X1 $T=72630 68200 1 0 $X=72515 $Y=66685
X18026 1913 931 A[0] 1542 INV_X1 $T=73390 68200 0 0 $X=73275 $Y=68085
X18027 2198 931 A[0] 1912 INV_X1 $T=75480 68200 0 0 $X=75365 $Y=68085
X18028 1559 931 A[0] 2348 INV_X1 $T=77570 26200 0 180 $X=77075 $Y=24685
X18029 reset 931 A[0] 783 INV_X1 $T=79660 65400 1 180 $X=79165 $Y=65285
X18030 1572 931 A[0] 2435 INV_X1 $T=80800 20600 0 0 $X=80685 $Y=20485
X18031 1989 960 931 167 166 A[0] 1191 1200 OAI221_X1 $T=13540 54200 0 0 $X=13425 $Y=54085
X18032 1662 205 931 211 214 A[0] 958 1203 OAI221_X1 $T=16960 59800 1 0 $X=16845 $Y=58285
X18033 2040 1265 931 275 286 A[0] 1266 1251 OAI221_X1 $T=22280 76600 0 0 $X=22165 $Y=76485
X18034 1823 1416 931 488 493 A[0] 1807 966 OAI221_X1 $T=48880 12200 0 0 $X=48765 $Y=12085
X18035 751 769 931 736 735 A[0] 718 2194 OAI221_X1 $T=74530 71000 1 180 $X=73275 $Y=70885
X18036 1903 1552 931 709 739 A[0] 1551 1545 OAI221_X1 $T=73770 68200 0 0 $X=73655 $Y=68085
X18037 2427 1587 931 868 861 A[0] 1923 1097 OAI221_X1 $T=81940 12200 0 180 $X=80685 $Y=10685
X18038 1097 686 1529 931 641 1879 A[0] AOI211_X1 $T=69400 9400 0 0 $X=69285 $Y=9285
X18039 2348 428 2203 931 997 1094 A[0] AOI211_X1 $T=77190 23400 0 0 $X=77075 $Y=23285
X18040 1101 840 1575 931 reset 792 A[0] AOI211_X1 $T=81560 68200 1 180 $X=80495 $Y=68085
X18349 931 A[0] 1990 247 1208 931 ICV_47 $T=17340 71000 0 0 $X=17225 $Y=70885
X18350 931 A[0] 1033 965 963 931 ICV_47 $T=17530 9400 1 0 $X=17415 $Y=7885
X18351 931 A[0] 985 788 1672 2528 ICV_47 $T=18100 1000 0 0 $X=17985 $Y=885
X18352 931 A[0] 1242 1221 1996 931 ICV_47 $T=18670 76600 0 0 $X=18555 $Y=76485
X18353 931 A[0] 985 980 272 931 ICV_47 $T=22280 51400 0 0 $X=22165 $Y=51285
X18354 931 A[0] 1036 503 990 931 ICV_47 $T=26270 23400 1 0 $X=26155 $Y=21885
X18355 931 A[0] 1007 989 2383 931 ICV_47 $T=28170 48600 1 0 $X=28055 $Y=47085
X18356 931 A[0] 973 1012 343 931 ICV_47 $T=32160 31800 0 0 $X=32045 $Y=31685
X18357 931 A[0] 931 980 355 931 ICV_47 $T=33110 79400 1 0 $X=32995 $Y=77885
X18358 931 A[0] 1007 788 2284 931 ICV_47 $T=33680 26200 1 0 $X=33565 $Y=24685
X18359 931 A[0] 1007 983 2281 931 ICV_47 $T=35580 23400 1 0 $X=35465 $Y=21885
X18360 931 A[0] 1009 1056 2057 931 ICV_47 $T=35580 29000 0 0 $X=35465 $Y=28885
X18361 931 A[0] 744 1025 2071 931 ICV_47 $T=39950 20600 0 0 $X=39835 $Y=20485
X18362 931 A[0] 319 981 2116 931 ICV_47 $T=49260 76600 0 0 $X=49145 $Y=76485
X18363 931 A[0] 995 660 1041 931 ICV_47 $T=50780 71000 1 0 $X=50665 $Y=69485
X18364 931 A[0] 1033 980 487 931 ICV_47 $T=51350 59800 0 0 $X=51235 $Y=59685
X18365 931 A[0] 258 983 565 931 ICV_47 $T=59900 23400 0 0 $X=59785 $Y=23285
X18366 931 A[0] 428 1025 589 931 ICV_47 $T=62370 20600 0 0 $X=62255 $Y=20485
X18367 931 A[0] 399 965 1489 931 ICV_47 $T=64270 31800 1 0 $X=64155 $Y=30285
X18368 931 A[0] 258 1056 772 931 ICV_47 $T=72630 26200 0 0 $X=72515 $Y=26085
X18369 931 A[0] 404 1056 1543 931 ICV_47 $T=73200 29000 0 0 $X=73085 $Y=28885
X18370 931 A[0] 973 788 264 ICV_48 $T=22280 31800 0 0 $X=22165 $Y=31685
X18371 931 A[0] 991 995 2028 ICV_48 $T=27220 37400 1 0 $X=27105 $Y=35885
X18372 931 A[0] 931 995 1010 ICV_48 $T=31590 73800 0 0 $X=31475 $Y=73685
X18373 931 A[0] 448 1056 2273 ICV_48 $T=32920 3800 0 0 $X=32805 $Y=3685
X18374 931 A[0] 1036 981 2277 ICV_48 $T=33490 17800 0 0 $X=33375 $Y=17685
X18375 931 A[0] 404 1025 2067 ICV_48 $T=37860 6600 1 0 $X=37745 $Y=5085
X18376 931 A[0] 501 980 398 ICV_48 $T=38240 51400 0 0 $X=38125 $Y=51285
X18377 931 A[0] 448 981 2083 ICV_48 $T=42230 62600 0 0 $X=42115 $Y=62485
X18378 931 A[0] 1033 1015 2121 ICV_48 $T=50020 34600 1 0 $X=49905 $Y=33085
X18379 931 A[0] 503 392 536 ICV_48 $T=52680 71000 1 0 $X=52565 $Y=69485
X18380 931 A[0] 258 986 2139 ICV_48 $T=57240 29000 0 0 $X=57125 $Y=28885
X18381 931 A[0] 931 1025 588 ICV_48 $T=57240 48600 0 0 $X=57125 $Y=48485
X18382 931 A[0] 744 995 1448 ICV_48 $T=57430 43000 1 0 $X=57315 $Y=41485
X18383 931 A[0] 506 997 1537 ICV_48 $T=70350 12200 1 0 $X=70235 $Y=10685
X18384 931 A[0] 931 1029 763 ICV_48 $T=71870 23400 0 0 $X=71755 $Y=23285
X18385 931 A[0] 1024 1012 2419 ICV_48 $T=74340 23400 0 0 $X=74225 $Y=23285
X18386 931 A[0] 744 1056 1550 ICV_48 $T=75290 12200 0 0 $X=75175 $Y=12085
X18387 931 A[0] 428 788 782 ICV_48 $T=77190 9400 0 0 $X=77075 $Y=9285
X18388 931 A[0] 428 1029 824 ICV_48 $T=79280 9400 1 0 $X=79165 $Y=7885
X18389 931 A[0] 931 997 825 ICV_48 $T=79280 17800 0 0 $X=79165 $Y=17685
X18390 931 A[0] 948 78 1151 ICV_49 $T=4800 43000 0 0 $X=4685 $Y=42885
X18391 931 A[0] 448 983 1316 ICV_49 $T=32730 9400 1 0 $X=32615 $Y=7885
X18392 931 A[0] 428 976 374 ICV_49 $T=33300 15000 0 0 $X=33185 $Y=14885
X18393 931 A[0] 164 1009 2052 ICV_49 $T=33300 48600 0 0 $X=33185 $Y=48485
X18394 931 A[0] 744 986 1028 ICV_49 $T=39190 31800 1 0 $X=39075 $Y=30285
X18395 931 A[0] 1033 989 2087 ICV_49 $T=42800 29000 1 0 $X=42685 $Y=27485
X18396 931 A[0] 931 965 1494 ICV_49 $T=62370 34600 0 0 $X=62255 $Y=34485
X18397 931 A[0] 973 338 620 ICV_49 $T=62370 51400 0 0 $X=62255 $Y=51285
X18398 931 A[0] 1024 1029 1581 ICV_49 $T=79280 3800 1 0 $X=79165 $Y=2285
X18399 931 A[0] 104 107 139 ICV_50 $T=10690 65400 1 0 $X=10575 $Y=63885
X18400 931 A[0] 104 83 158 ICV_50 $T=12210 73800 1 0 $X=12095 $Y=72285
X18401 931 A[0] 883 573 584 ICV_50 $T=59900 73800 1 0 $X=59785 $Y=72285
X18402 931 A[0] 1436 2417 712 ICV_50 $T=70350 34600 1 0 $X=70235 $Y=33085
X18403 931 A[0] 1436 2478 725 ICV_50 $T=71870 40200 0 0 $X=71755 $Y=40085
X18404 931 A[0] 883 700 765 ICV_50 $T=74720 62600 1 0 $X=74605 $Y=61085
X18405 931 A[0] 883 684 767 ICV_50 $T=75100 48600 0 0 $X=74985 $Y=48485
X18406 931 A[0] 883 717 805 ICV_50 $T=77570 45800 1 0 $X=77455 $Y=44285
X18407 931 A[0] 883 775 808 ICV_50 $T=77760 51400 0 0 $X=77645 $Y=51285
X18408 931 A[0] 883 728 815 ICV_50 $T=77950 57000 0 0 $X=77835 $Y=56885
X18409 931 A[0] 883 718 818 ICV_50 $T=77950 71000 1 0 $X=77835 $Y=69485
X18410 931 A[0] 883 1534 822 ICV_50 $T=78140 71000 0 0 $X=78025 $Y=70885
X18411 931 A[0] 883 732 836 ICV_50 $T=79090 48600 0 0 $X=78975 $Y=48485
X18412 931 A[0] 883 786 839 ICV_50 $T=79090 79400 0 0 $X=78975 $Y=79285
X18468 931 A[0] 931 655 387 ICV_52 $T=36910 12200 1 0 $X=36795 $Y=10685
X18469 931 A[0] 931 1056 1329 ICV_52 $T=36910 26200 1 0 $X=36795 $Y=24685
X18470 931 A[0] 506 1014 1051 ICV_52 $T=51350 40200 0 0 $X=51235 $Y=40085
X18471 931 A[0] 744 980 522 ICV_52 $T=52110 34600 0 0 $X=51995 $Y=34485
X18472 931 A[0] 258 788 533 ICV_52 $T=54960 23400 1 0 $X=54845 $Y=21885
X18473 931 A[0] 392 164 2173 ICV_52 $T=63890 48600 1 0 $X=63775 $Y=47085
X18474 931 A[0] 744 997 2202 ICV_52 $T=77000 12200 0 0 $X=76885 $Y=12085
X18475 931 A[0] 1080 1056 2210 ICV_52 $T=78520 3800 0 0 $X=78405 $Y=3685
X18476 931 A[0] 1036 1029 2357 ICV_52 $T=78900 20600 0 0 $X=78785 $Y=20485
X18477 931 A[0] 1033 1020 1982 ICV_53 $T=13350 3800 1 180 $X=12665 $Y=3685
X18478 931 A[0] 506 655 1983 ICV_53 $T=15250 17800 0 180 $X=14565 $Y=16285
X18479 931 A[0] 506 338 1988 ICV_53 $T=16770 20600 1 180 $X=16085 $Y=20485
X18480 931 A[0] 744 1015 2010 ICV_53 $T=22850 45800 1 180 $X=22165 $Y=45685
X18481 931 A[0] 428 1015 987 ICV_53 $T=25700 17800 0 180 $X=25015 $Y=16285
X18482 931 A[0] 976 1022 1289 ICV_53 $T=28360 65400 1 180 $X=27675 $Y=65285
X18483 931 A[0] 1033 975 1293 ICV_53 $T=29690 45800 1 180 $X=29005 $Y=45685
X18484 931 A[0] 1024 989 1299 ICV_53 $T=30450 17800 0 180 $X=29765 $Y=16285
X18485 931 A[0] 319 1014 2274 ICV_53 $T=31210 79400 0 180 $X=30525 $Y=77885
X18486 931 A[0] 1033 1009 2279 ICV_53 $T=35770 59800 0 180 $X=35085 $Y=58285
X18487 931 A[0] 319 392 1744 ICV_53 $T=36150 79400 1 180 $X=35465 $Y=79285
X18488 931 A[0] 1022 1056 1331 ICV_53 $T=37860 29000 0 180 $X=37175 $Y=27485
X18489 931 A[0] 404 986 1399 ICV_53 $T=48500 34600 0 180 $X=47815 $Y=33085
X18490 931 A[0] 258 1012 479 ICV_53 $T=50210 6600 1 180 $X=49525 $Y=6485
X18491 931 A[0] 404 965 2115 ICV_53 $T=51540 6600 0 180 $X=50855 $Y=5085
X18492 931 A[0] 989 319 525 ICV_53 $T=52870 71000 1 180 $X=52185 $Y=70885
X18493 931 A[0] 448 655 1055 ICV_53 $T=53250 23400 1 180 $X=52565 $Y=23285
X18494 931 A[0] 1024 164 2313 ICV_53 $T=53440 23400 0 180 $X=52755 $Y=21885
X18495 931 A[0] 931 1020 555 ICV_53 $T=59900 34600 1 180 $X=59215 $Y=34485
X18496 931 A[0] 664 975 1516 ICV_53 $T=69020 31800 1 180 $X=68335 $Y=31685
X18497 931 A[0] 1007 1025 638 ICV_53 $T=69020 34600 1 180 $X=68335 $Y=34485
X18498 931 A[0] 258 1011 713 ICV_53 $T=71110 29000 1 180 $X=70425 $Y=28885
X18499 931 A[0] 991 965 2200 ICV_53 $T=75290 20600 0 180 $X=74605 $Y=19085
X18500 931 A[0] 428 1056 807 ICV_53 $T=77760 17800 1 180 $X=77075 $Y=17685
X18501 931 A[0] 1036 1012 2424 ICV_53 $T=79470 9400 1 180 $X=78785 $Y=9285
X18527 1048 1052 931 507 509 512 A[0] 1422 1416 OAI222_X1 $T=51160 12200 1 0 $X=51045 $Y=10685
X18528 1078 643 931 659 649 663 A[0] 1519 641 OAI222_X1 $T=66550 6600 0 0 $X=66435 $Y=6485
X18529 1094 2205 931 820 799 829 A[0] 869 1572 OAI222_X1 $T=78710 23400 1 0 $X=78595 $Y=21885
X18551 1005 Res[4] 50 931 A[0] Res[1] 25 ICV_55 $T=4230 62600 1 180 $X=2215 $Y=62485
X18552 104 79 80 931 A[0] 62 46 ICV_55 $T=6130 54200 0 180 $X=4115 $Y=52685
X18553 104 81 112 931 A[0] 76 89 ICV_55 $T=8790 57000 0 180 $X=6775 $Y=55485
X18554 1005 Res[21] 131 931 A[0] Res[20] 108 ICV_55 $T=10500 82200 1 180 $X=8485 $Y=82085
X18555 104 44 213 931 A[0] 52 181 ICV_55 $T=16390 76600 0 180 $X=14375 $Y=75085
X18556 1005 Res[24] 558 931 A[0] Res[23] 544 ICV_55 $T=58190 82200 1 180 $X=56175 $Y=82085
X18557 1436 1488 633 931 A[0] 1863 613 ICV_55 $T=64270 57000 1 180 $X=62255 $Y=56885
X18558 1005 Res[28] 671 931 A[0] Res[26] 642 ICV_55 $T=66930 82200 1 180 $X=64915 $Y=82085
X18559 1436 1538 729 931 A[0] 1083 705 ICV_55 $T=72250 57000 1 180 $X=70235 $Y=56885
X18560 883 695 777 931 A[0] 687 741 ICV_55 $T=75670 62600 1 180 $X=73655 $Y=62485
X18561 1436 1563 800 931 A[0] 2346 773 ICV_55 $T=77570 31800 0 180 $X=75555 $Y=30285
X18562 883 665 837 931 A[0] 672 795 ICV_55 $T=79280 57000 0 180 $X=77265 $Y=55485
X18563 883 761 867 931 A[0] 693 816 ICV_55 $T=80230 59800 1 180 $X=78215 $Y=59685
X18597 985 A[0] 965 1179 931 1640 132 1195 1983 58 ICV_57 $T=10500 17800 1 0 $X=10385 $Y=16285
X18598 258 A[0] 655 236 931 1223 236 1679 2001 100 ICV_57 $T=18290 23400 0 0 $X=18175 $Y=23285
X18599 1036 A[0] 995 2017 931 2243 299 1794 2088 2234 ICV_57 $T=23990 31800 0 0 $X=23875 $Y=31685
X18600 428 A[0] 1014 228 931 2255 304 1282 2031 263 ICV_57 $T=24180 31800 1 0 $X=24065 $Y=30285
X18601 1036 A[0] 1009 2029 931 351 2493 2036 2042 2032 ICV_57 $T=27600 31800 0 0 $X=27485 $Y=31685
X18602 995 A[0] 319 1284 931 2266 332 1010 2384 1730 ICV_57 $T=27980 76600 1 0 $X=27865 $Y=75085
X18603 1036 A[0] 1015 2059 931 2391 396 1346 427 1757 ICV_57 $T=36340 17800 1 0 $X=36225 $Y=16285
X18604 1024 A[0] 975 2289 931 2271 422 1027 1751 1763 ICV_57 $T=38240 15000 0 0 $X=38125 $Y=14885
X18605 1080 A[0] 980 410 931 1341 411 2074 2293 414 ICV_57 $T=38240 34600 0 0 $X=38125 $Y=34485
X18606 975 A[0] 392 2068 931 2288 1759 2077 1775 1769 ICV_57 $T=38240 57000 0 0 $X=38125 $Y=56885
X18607 664 A[0] 503 424 931 397 424 1360 2081 2077 ICV_57 $T=38240 62600 1 0 $X=38125 $Y=61085
X18608 1033 A[0] 1012 2392 931 1343 2495 1778 1761 1773 ICV_57 $T=38430 3800 0 0 $X=38315 $Y=3685
X18609 664 A[0] 1056 431 931 434 2468 1418 2111 455 ICV_57 $T=42040 3800 0 0 $X=41925 $Y=3685
X18610 1007 A[0] 995 2092 931 2296 466 1390 2122 2110 ICV_57 $T=44510 79400 1 0 $X=44395 $Y=77885
X18611 1000 A[0] 975 1373 931 2469 474 1395 2398 1382 ICV_57 $T=44890 23400 1 0 $X=44775 $Y=21885
X18612 931 A[0] 1025 477 931 2099 477 1401 2113 1804 ICV_57 $T=45650 15000 1 0 $X=45535 $Y=13485
X18613 1080 A[0] 1009 2125 931 2315 522 1059 2125 526 ICV_57 $T=53440 37400 1 0 $X=53325 $Y=35885
X18614 931 A[0] 981 2130 931 510 525 1439 2130 1378 ICV_57 $T=54010 73800 1 0 $X=53895 $Y=72285
X18615 1009 A[0] 1012 540 931 2114 549 1464 2405 1466 ICV_57 $T=57050 37400 1 0 $X=56935 $Y=35885
X18616 428 A[0] 164 562 931 2406 1854 1473 1853 1491 ICV_57 $T=59520 15000 0 0 $X=59405 $Y=14885
X18617 1000 A[0] 997 2153 931 2407 589 1481 1864 1862 ICV_57 $T=60090 20600 1 0 $X=59975 $Y=19085
X18618 985 A[0] 976 2340 931 1502 656 1516 2340 645 ICV_57 $T=65600 31800 1 0 $X=65485 $Y=30285
X18619 1036 A[0] 1025 2344 931 1527 1885 2418 2344 2341 ICV_57 $T=69780 17800 1 0 $X=69665 $Y=16285
X18620 991 A[0] 983 1578 931 2365 807 1578 2357 869 ICV_57 $T=77760 20600 1 0 $X=77645 $Y=19085
X18621 1080 A[0] 1011 863 931 2207 825 863 1920 875 ICV_57 $T=78330 17800 1 0 $X=78215 $Y=16285
X18622 506 A[0] 164 2232 931 506 1025 1194 ICV_58 $T=14490 6600 0 180 $X=13805 $Y=5085
X18623 664 A[0] 1029 187 931 664 788 109 ICV_58 $T=19240 3800 0 180 $X=18555 $Y=2285
X18624 258 A[0] 975 308 931 931 1015 309 ICV_58 $T=26650 26200 0 180 $X=25965 $Y=24685
X18625 1022 A[0] 980 332 931 1022 319 2034 ICV_58 $T=30070 73800 1 180 $X=29385 $Y=73685
X18626 399 A[0] 980 419 931 931 1014 2484 ICV_58 $T=39570 76600 1 180 $X=38885 $Y=76485
X18627 991 A[0] 976 2100 931 428 975 456 ICV_58 $T=45840 20600 0 180 $X=45155 $Y=19085
X18628 1033 A[0] 1029 1802 931 448 997 2111 ICV_58 $T=48500 3800 1 180 $X=47815 $Y=3685
X18629 503 A[0] 399 473 931 503 1022 492 ICV_58 $T=49260 76600 0 180 $X=48575 $Y=75085
X18630 973 A[0] 1025 497 931 931 1020 489 ICV_58 $T=50970 23400 0 180 $X=50285 $Y=21885
X18631 744 A[0] 965 1064 931 404 1012 1442 ICV_58 $T=57430 23400 0 180 $X=56745 $Y=21885
X18632 931 A[0] 788 2324 931 1022 1029 2160 ICV_58 $T=61040 26200 0 180 $X=60355 $Y=24685
X18633 660 A[0] 975 1074 931 1007 655 1499 ICV_58 $T=65980 51400 0 180 $X=65295 $Y=49885
X18634 991 A[0] 1056 2481 931 428 1011 771 ICV_58 $T=76620 23400 1 180 $X=75935 $Y=23285
X18635 428 A[0] 983 804 931 1036 788 1558 ICV_58 $T=77760 17800 0 180 $X=77075 $Y=16285
X18636 991 A[0] 1012 1095 931 991 788 1561 ICV_58 $T=77950 12200 0 180 $X=77265 $Y=10685
X18637 722 756 734 747 931 A[0] 1907 OR4_X1 $T=75670 79400 1 180 $X=74415 $Y=79285
X18638 735 751 752 759 931 A[0] 1536 OR4_X1 $T=74910 73800 0 0 $X=74795 $Y=73685
X18639 1907 752 690 691 931 A[0] 2196 OR4_X1 $T=74910 76600 1 0 $X=74795 $Y=75085
X18640 1564 759 776 778 931 A[0] 1914 OR4_X1 $T=76050 73800 0 0 $X=75935 $Y=73685
X18641 1540 786 787 557 931 A[0] 1564 OR4_X1 $T=77000 76600 0 0 $X=76885 $Y=76485
X18659 931 A[0] 501 1025 132 ICV_61 $T=12590 15000 0 0 $X=12475 $Y=14885
X18660 931 A[0] 404 338 1679 ICV_61 $T=19620 23400 1 0 $X=19505 $Y=21885
X18661 931 A[0] 973 983 293 ICV_61 $T=25320 20600 1 0 $X=25205 $Y=19085
X18662 931 A[0] 664 1025 2493 ICV_61 $T=29120 34600 1 0 $X=29005 $Y=33085
X18663 931 A[0] 985 319 2272 ICV_61 $T=32920 65400 1 0 $X=32805 $Y=63885
X18664 931 A[0] 258 1020 379 ICV_61 $T=36150 9400 1 0 $X=36035 $Y=7885
X18665 931 A[0] 1000 319 2066 ICV_61 $T=37100 62600 0 0 $X=36985 $Y=62485
X18666 931 A[0] 985 338 435 ICV_61 $T=42230 23400 0 0 $X=42115 $Y=23285
X18667 931 A[0] 986 392 1394 ICV_61 $T=49830 71000 0 0 $X=49715 $Y=70885
X18668 931 A[0] 1033 986 2475 ICV_61 $T=52490 43000 1 0 $X=52375 $Y=41485
X18669 931 A[0] 973 995 2128 ICV_61 $T=53060 82200 1 0 $X=52945 $Y=80685
X18670 931 A[0] 660 319 2127 ICV_61 $T=53630 76600 0 0 $X=53515 $Y=76485
X18671 931 A[0] 1000 1056 2318 ICV_61 $T=54390 3800 0 0 $X=54275 $Y=3685
X18672 931 A[0] 399 1012 2133 ICV_61 $T=55340 23400 0 0 $X=55225 $Y=23285
X18673 931 A[0] 404 1009 2135 ICV_61 $T=55910 51400 0 0 $X=55795 $Y=51285
X18674 931 A[0] 404 980 569 ICV_61 $T=56290 40200 0 0 $X=56175 $Y=40085
X18675 931 A[0] 664 989 576 ICV_61 $T=58760 54200 0 0 $X=58645 $Y=54085
X18676 931 A[0] 1033 997 1505 ICV_61 $T=66930 26200 0 0 $X=66815 $Y=26085
X18677 931 A[0] 660 655 2180 ICV_61 $T=67120 37400 1 0 $X=67005 $Y=35885
X18678 931 A[0] 1534 710 1532 ICV_61 $T=70920 71000 0 0 $X=70805 $Y=70885
X18679 931 A[0] 744 1029 2420 ICV_61 $T=74910 26200 1 0 $X=74795 $Y=24685
X18680 931 A[0] 1036 983 1555 ICV_61 $T=76620 23400 1 0 $X=76505 $Y=21885
X18681 clk 931 A[0] 674 CLKBUF_X3 $T=2900 82200 0 0 $X=2785 $Y=82085
X18682 524 931 A[0] 319 CLKBUF_X3 $T=54770 65400 0 0 $X=54655 $Y=65285
X18683 93 931 A[0] 538 CLKBUF_X3 $T=57620 68200 0 180 $X=56555 $Y=66685
X18684 1085 931 A[0] 883 CLKBUF_X3 $T=75480 59800 0 0 $X=75365 $Y=59685
X18685 783 931 A[0] 870 CLKBUF_X3 $T=77190 65400 0 180 $X=76125 $Y=63885
X18686 957 138 931 A[0] 1667 OR2_X1 $T=15820 51400 0 0 $X=15705 $Y=51285
X18687 248 273 931 A[0] 1248 OR2_X1 $T=22280 73800 1 0 $X=22165 $Y=72285
X18688 747 543 931 A[0] 2140 OR2_X1 $T=56860 79400 0 0 $X=56745 $Y=79285
X18689 710 718 931 A[0] 752 OR2_X1 $T=74910 73800 1 180 $X=74035 $Y=73685
X18690 1534 769 931 A[0] 759 OR2_X1 $T=76050 73800 1 0 $X=75935 $Y=72285
X18691 2239 A[0] 138 1182 931 161 NOR3_X1 $T=12970 48600 0 0 $X=12855 $Y=48485
X18692 1661 A[0] 1987 1657 931 183 NOR3_X1 $T=15630 15000 0 0 $X=15515 $Y=14885
X18693 1999 A[0] 247 248 931 972 NOR3_X1 $T=19240 71000 0 0 $X=19125 $Y=70885
X18694 775 A[0] 755 758 931 746 NOR3_X1 $T=76620 51400 1 180 $X=75745 $Y=51285
X18695 749 A[0] 827 740 931 2201 NOR3_X1 $T=76050 37400 1 0 $X=75935 $Y=35885
X18708 786 787 1901 931 A[0] 751 AND3_X1 $T=73390 76600 0 0 $X=73275 $Y=76485
X18709 756 734 1553 931 A[0] 735 AND3_X1 $T=75860 79400 1 0 $X=75745 $Y=77885
X18775 1137 931 940 61 A[0] 942 NAND3_X1 $T=5560 45800 0 0 $X=5445 $Y=45685
X18776 2194 931 1551 1552 A[0] 2342 NAND3_X1 $T=72250 71000 1 0 $X=72135 $Y=69485
X18777 2195 931 2201 1892 A[0] 1903 NAND3_X1 $T=73960 45800 0 0 $X=73845 $Y=45685
X18778 769 931 751 1534 A[0] 1551 NAND3_X1 $T=74530 71000 0 0 $X=74415 $Y=70885
X18779 1089 931 746 1092 A[0] 739 NAND3_X1 $T=74720 59800 0 0 $X=74605 $Y=59685
X18780 718 931 735 710 A[0] 1552 NAND3_X1 $T=75290 73800 1 0 $X=75175 $Y=72285
X18781 1107 1108 931 23 933 1112 A[0] OAI22_X1 $T=2330 34600 1 0 $X=2215 $Y=33085
X18782 1971 1182 931 1183 137 1186 A[0] OAI22_X1 $T=10880 48600 0 0 $X=10765 $Y=48485
X18783 954 1663 931 163 1207 177 A[0] OAI22_X1 $T=14300 62600 1 0 $X=14185 $Y=61085
X18784 960 1989 931 1649 1367 2095 A[0] OAI22_X1 $T=16200 54200 1 0 $X=16085 $Y=52685
X18785 1212 1990 931 1211 1994 1241 A[0] OAI22_X1 $T=17340 73800 0 180 $X=16275 $Y=72285
X18786 231 1221 931 249 1233 1239 A[0] OAI22_X1 $T=19430 79400 0 0 $X=19315 $Y=79285
X18787 1533 1904 931 1529 1887 1525 A[0] OAI22_X1 $T=71300 9400 0 180 $X=70235 $Y=7885
X18788 739 1914 931 737 2196 1903 A[0] OAI22_X1 $T=75290 71000 0 180 $X=74225 $Y=69485
X18789 2196 1551 931 2198 1552 1914 A[0] OAI22_X1 $T=75290 71000 0 0 $X=75175 $Y=70885
X18822 1945 16 2382 1598 A[0] 931 57 1959 57 1964 1632 1125 931 ICV_66 $T=2330 6600 0 0 $X=2215 $Y=6485
X18823 1947 1118 1127 1606 A[0] 931 1134 2442 59 1157 2229 77 931 ICV_66 $T=2330 20600 1 0 $X=2215 $Y=19085
X18824 1147 34 1136 1617 A[0] 931 936 1622 74 1164 1781 75 931 ICV_66 $T=3090 40200 1 0 $X=2975 $Y=38685
X18825 42 58 1965 1714 A[0] 931 1630 1633 1646 1179 2371 1965 931 ICV_66 $T=5370 15000 0 0 $X=5255 $Y=14885
X18826 1626 86 1170 2233 A[0] 931 160 210 121 974 1981 952 931 ICV_66 $T=7080 9400 1 0 $X=6965 $Y=7885
X18827 1180 1705 1184 1106 A[0] 931 2228 1184 142 955 1236 147 931 ICV_66 $T=8410 29000 0 0 $X=8295 $Y=28885
X18828 2370 2446 1003 999 A[0] 931 88 159 147 1198 2240 41 931 ICV_66 $T=9170 31800 1 0 $X=9055 $Y=30285
X18829 1967 120 1979 984 A[0] 931 153 2241 159 1985 184 1664 931 ICV_66 $T=9930 34600 0 0 $X=9815 $Y=34485
X18830 128 153 1984 2241 A[0] 931 33 1204 193 1991 2246 1674 931 ICV_66 $T=12590 37400 0 0 $X=12475 $Y=37285
X18831 1196 156 1766 2242 A[0] 931 90 1665 197 1992 1660 1985 931 ICV_66 $T=12780 43000 0 0 $X=12665 $Y=42885
X18832 964 228 1693 2017 A[0] 931 1236 237 266 1702 1255 1699 931 ICV_66 $T=18290 29000 0 0 $X=18175 $Y=28885
X18833 2246 229 1729 1724 A[0] 931 1683 2452 270 1980 1709 291 931 ICV_66 $T=18480 40200 1 0 $X=18365 $Y=38685
X18834 2223 252 2008 1243 A[0] 931 253 289 1262 1275 1287 315 2528 ICV_66 $T=19620 1000 0 0 $X=19505 $Y=885
X18835 1964 253 1245 1249 A[0] 931 150 1249 289 1272 305 1240 931 ICV_66 $T=20000 6600 1 0 $X=19885 $Y=5085
X18836 974 1290 1291 1689 A[0] 931 310 2382 2055 1001 1302 1245 931 ICV_66 $T=22280 6600 0 0 $X=22165 $Y=6485
X18837 193 279 1006 1706 A[0] 931 1704 1709 311 2028 2029 280 931 ICV_66 $T=22280 37400 0 0 $X=22165 $Y=37285
X18838 281 2381 1274 1716 A[0] 931 1713 2262 996 1292 1013 1724 931 ICV_66 $T=23420 43000 1 0 $X=23305 $Y=41485
X18839 1973 987 1286 990 A[0] 931 1279 122 1296 1728 1299 1725 931 ICV_66 $T=23610 15000 0 0 $X=23495 $Y=14885
X18840 182 310 1700 1308 A[0] 931 1719 1291 329 1269 2271 1307 931 ICV_66 $T=25320 9400 0 0 $X=25205 $Y=9285
X18841 2265 315 1731 2070 A[0] 931 329 1272 334 1313 2273 1731 2528 ICV_66 $T=26270 1000 0 0 $X=26155 $Y=885
X18842 1295 333 2385 2039 A[0] 931 255 2385 349 1321 2279 378 931 ICV_66 $T=29120 59800 1 0 $X=29005 $Y=58285
X18843 1301 340 1309 1734 A[0] 931 1736 2275 1326 2052 2054 1325 931 ICV_66 $T=30450 51400 1 0 $X=30335 $Y=49885
X18844 224 342 2045 2276 A[0] 931 1215 2249 365 1752 1384 342 931 ICV_66 $T=30830 54200 0 0 $X=30715 $Y=54085
X18845 192 346 1742 1795 A[0] 931 1186 383 371 2060 2460 394 931 ICV_66 $T=31780 45800 0 0 $X=31665 $Y=45685
X18846 1357 356 1318 2282 A[0] 931 1206 1323 381 1324 2286 1318 931 ICV_66 $T=32730 40200 1 0 $X=32615 $Y=38685
X18847 2456 361 2053 2284 A[0] 931 322 2459 389 2063 1331 1755 931 ICV_66 $T=33110 26200 0 0 $X=32995 $Y=26085
X18848 1312 364 2058 378 A[0] 931 352 2390 395 2068 2290 423 931 ICV_66 $T=33680 59800 0 0 $X=33565 $Y=59685
X18849 317 1325 1366 1746 A[0] 931 384 1746 398 1348 1023 1759 931 ICV_66 $T=34060 54200 1 0 $X=33945 $Y=52685
X18850 357 380 1335 1755 A[0] 931 984 2286 410 1347 1758 433 931 ICV_66 $T=35770 34600 1 0 $X=35655 $Y=33085
X18851 1743 385 2065 1330 A[0] 931 296 405 418 1792 1796 265 931 ICV_66 $T=35770 71000 0 0 $X=35655 $Y=70885
X18852 2038 386 1754 2096 A[0] 931 1239 1754 420 1772 1760 459 931 ICV_66 $T=35770 82200 0 0 $X=35655 $Y=82085
X18853 369 388 1327 2066 A[0] 931 416 1345 426 1363 2083 1775 931 ICV_66 $T=35960 65400 1 0 $X=35845 $Y=63885
X18854 1271 405 2072 2291 A[0] 931 1994 1362 2396 2086 2105 2072 931 ICV_66 $T=38430 73800 0 0 $X=38315 $Y=73685
X18855 2463 2462 2078 2295 A[0] 931 412 1037 2469 2090 2300 1784 931 ICV_66 $T=39190 26200 0 0 $X=39075 $Y=26085
X18856 1027 430 1757 1764 A[0] 931 467 1370 456 2100 1389 430 931 ICV_66 $T=40900 17800 0 0 $X=40785 $Y=17685
X18857 2079 433 2085 1785 A[0] 931 2088 2091 460 1399 2397 490 931 ICV_66 $T=41470 31800 0 0 $X=41355 $Y=31685
X18858 2076 2464 1396 1043 A[0] 931 346 1788 1873 1044 482 1396 931 ICV_66 $T=42040 45800 0 0 $X=41925 $Y=45685
X18859 2078 2087 1035 2301 A[0] 931 1785 1047 468 2106 2308 413 931 ICV_66 $T=42230 29000 0 0 $X=42115 $Y=28885
X18860 2464 1040 1341 1474 A[0] 931 1787 2094 1497 1392 2309 1040 931 ICV_66 $T=42230 43000 1 0 $X=42115 $Y=41485
X18861 1367 1798 2465 1034 A[0] 931 1202 1376 469 1799 2129 1798 931 ICV_66 $T=42230 51400 0 0 $X=42115 $Y=51285
X18862 2280 1797 1377 1800 A[0] 931 1790 2058 1045 1393 2310 1800 931 ICV_66 $T=42230 59800 1 0 $X=42115 $Y=58285
X18863 2086 445 1378 2298 A[0] 931 1792 2305 473 1394 1410 445 931 ICV_66 $T=42230 73800 1 0 $X=42115 $Y=72285
X18864 440 449 1382 1803 A[0] 931 1794 2090 476 1398 2311 1803 931 ICV_66 $T=42800 26200 1 0 $X=42685 $Y=24685
X18865 469 483 1408 1814 A[0] 931 429 2473 502 1419 1820 483 931 ICV_66 $T=47360 51400 1 0 $X=47245 $Y=49885
X18866 2399 494 1412 2314 A[0] 931 1815 2310 515 1425 1057 480 931 ICV_66 $T=48880 62600 1 0 $X=48765 $Y=61085
X18867 1819 516 2471 1066 A[0] 931 443 2106 1818 1838 2166 436 931 ICV_66 $T=52300 26200 0 0 $X=52185 $Y=26085
X18868 1045 1463 2401 2134 A[0] 931 485 2138 545 1455 2506 2137 931 ICV_66 $T=53630 59800 1 0 $X=53515 $Y=58285
X18869 2132 530 1801 1841 A[0] 931 521 1841 2174 1848 1065 2157 931 ICV_66 $T=55340 6600 0 0 $X=55225 $Y=6485
X18870 1046 533 1442 1064 A[0] 931 1843 1846 564 2159 2153 1854 931 ICV_66 $T=55910 20600 0 0 $X=55795 $Y=20485
X18871 567 534 2139 1454 A[0] 931 1443 2405 567 2497 1502 1855 931 ICV_66 $T=55910 31800 1 0 $X=55795 $Y=30285
X18872 553 1845 2438 1070 A[0] 931 523 1460 570 2142 2155 609 931 ICV_66 $T=55910 45800 0 0 $X=55795 $Y=45685
X18873 571 576 1476 2325 A[0] 931 611 2162 620 1074 2412 1496 931 ICV_66 $T=59900 54200 1 0 $X=59785 $Y=52685
X18874 2159 2491 1486 2326 A[0] 931 1866 1493 631 1509 2190 692 931 ICV_66 $T=61610 26200 1 0 $X=61495 $Y=24685
X18875 612 603 1869 1861 A[0] 931 659 1498 644 1894 2185 1519 931 ICV_66 $T=62370 9400 0 0 $X=62255 $Y=9285
X18876 1070 608 1073 2329 A[0] 931 2150 608 646 2179 2182 2186 931 ICV_66 $T=62370 40200 0 0 $X=62255 $Y=40085
X18877 680 1859 1900 670 A[0] 931 1511 2413 680 1890 2343 1528 931 ICV_66 $T=65410 79400 0 0 $X=65295 $Y=79285
X18878 1520 1539 2193 1537 A[0] 931 679 1539 727 1549 2489 1911 931 ICV_66 $T=69590 15000 0 0 $X=69475 $Y=14885
X18879 1909 762 1093 1939 A[0] 931 1908 757 806 2210 2204 1924 2528 ICV_66 $T=75290 1000 0 0 $X=75175 $Y=885
X18880 1000 A[0] 1025 2238 931 1161 119 2436 2238 1650 931 ICV_67 $T=9930 23400 1 0 $X=9815 $Y=21885
X18881 501 A[0] 164 127 931 70 127 1658 1988 1653 931 ICV_67 $T=10880 20600 0 0 $X=10765 $Y=20485
X18882 506 A[0] 1020 1675 931 1986 191 963 1675 A[0] 931 ICV_67 $T=15440 6600 0 0 $X=15325 $Y=6485
X18883 404 A[0] 164 1230 931 2374 222 1230 1998 1682 931 ICV_67 $T=17910 12200 1 0 $X=17795 $Y=10685
X18884 931 A[0] 981 260 931 240 241 1683 1665 1984 931 ICV_67 $T=18860 43000 0 0 $X=18745 $Y=42885
X18885 404 A[0] 989 1247 931 1678 251 1247 2010 1690 931 ICV_67 $T=19430 48600 1 0 $X=19315 $Y=47085
X18886 501 A[0] 995 1321 931 2387 352 1736 2280 2276 931 ICV_67 $T=32350 57000 0 0 $X=32235 $Y=56885
X18887 392 A[0] 788 1753 931 2458 377 1334 1753 1335 931 ICV_67 $T=35580 31800 1 0 $X=35465 $Y=30285
X18888 1000 A[0] 1029 452 931 1355 431 2084 452 1778 2528 ICV_67 $T=41090 1000 0 0 $X=40975 $Y=885
X18889 448 A[0] 1015 1381 931 437 447 1381 2303 1385 931 ICV_67 $T=42610 65400 1 0 $X=42495 $Y=63885
X18890 991 A[0] 975 1404 931 2470 2101 1404 1411 1407 931 ICV_67 $T=46600 17800 1 0 $X=46485 $Y=16285
X18891 1033 A[0] 983 518 931 1806 505 518 1058 542 931 ICV_67 $T=50780 17800 1 0 $X=50665 $Y=16285
X18892 1022 A[0] 981 1826 931 2122 510 1417 1826 1824 931 ICV_67 $T=51350 73800 0 0 $X=51235 $Y=73685
X18893 1033 A[0] 1014 1840 931 2401 531 2437 1840 545 931 ICV_67 $T=55530 62600 1 0 $X=55415 $Y=61085
X18894 931 A[0] 1011 806 931 762 757 784 2199 770 931 ICV_67 $T=74910 3800 0 0 $X=74795 $Y=3685
X18895 1897 1852 1893 1895 931 A[0] 2195 AND4_X1 $T=71870 48600 1 0 $X=71755 $Y=47085
X18896 1891 1874 1541 1899 931 A[0] 1089 AND4_X1 $T=72820 59800 0 0 $X=72705 $Y=59685
X18897 776 778 1540 557 931 A[0] 1901 AND4_X1 $T=74910 76600 0 180 $X=73655 $Y=75085
X18898 690 691 722 747 931 A[0] 1553 AND4_X1 $T=74720 79400 1 0 $X=74605 $Y=77885
X18945 931 A[0] 744 976 2004 ICV_69 $T=20950 15000 0 0 $X=20835 $Y=14885
X18946 931 A[0] 428 981 278 ICV_69 $T=22280 23400 0 0 $X=22165 $Y=23285
X18947 931 A[0] 448 986 1259 ICV_69 $T=23800 65400 1 0 $X=23685 $Y=63885
X18948 931 A[0] 404 1015 1270 ICV_69 $T=26080 48600 1 0 $X=25965 $Y=47085
X18949 931 A[0] 428 989 373 ICV_69 $T=31970 17800 0 0 $X=31855 $Y=17685
X18950 931 A[0] 1007 503 366 ICV_69 $T=33300 73800 0 0 $X=33185 $Y=73685
X18951 931 A[0] 931 983 727 ICV_69 $T=73390 17800 1 0 $X=73275 $Y=16285
X18952 931 A[0] 428 1012 742 ICV_69 $T=74340 20600 0 0 $X=74225 $Y=20485
X18953 104 63 96 931 A[0] ICV_70 $T=7650 51400 1 0 $X=7535 $Y=49885
X18954 104 116 105 931 A[0] ICV_70 $T=8030 62600 0 0 $X=7915 $Y=62485
X18955 104 1627 117 931 A[0] ICV_70 $T=9360 59800 0 0 $X=9245 $Y=59685
X18956 104 135 126 931 A[0] ICV_70 $T=10310 68200 1 0 $X=10195 $Y=66685
X18957 1436 1835 538 931 A[0] ICV_70 $T=55720 65400 0 0 $X=55605 $Y=65285
X18958 1436 1504 657 931 A[0] ICV_70 $T=65980 62600 0 0 $X=65865 $Y=62485
X18959 883 716 743 931 A[0] ICV_70 $T=73770 45800 1 0 $X=73655 $Y=44285
X18960 1436 1905 748 931 A[0] ICV_70 $T=74150 29000 1 0 $X=74035 $Y=27485
X18961 931 A[0] 2446 151 1976 1680 947 ICV_71 $T=10500 26200 0 0 $X=10385 $Y=26085
X18962 931 A[0] 1150 173 150 1975 1981 ICV_71 $T=12210 6600 0 0 $X=12095 $Y=6485
X18963 931 A[0] 239 2448 2451 1227 238 ICV_71 $T=18670 34600 0 0 $X=18555 $Y=34485
X18964 931 A[0] 323 354 1307 2393 967 ICV_71 $T=30640 12200 1 0 $X=30525 $Y=10685
X18965 931 A[0] 2260 373 1314 2277 1735 ICV_71 $T=33110 17800 1 0 $X=32995 $Y=16285
X18966 931 A[0] 333 397 1345 2390 364 ICV_71 $T=35010 62600 1 0 $X=34895 $Y=61085
X18967 931 A[0] 353 1762 1779 1780 2297 ICV_71 $T=38620 9400 1 0 $X=38505 $Y=7885
X18968 931 A[0] 2316 519 2475 1051 1808 ICV_71 $T=50780 43000 0 0 $X=50665 $Y=42885
X18969 931 A[0] 2109 548 2402 1061 1435 ICV_71 $T=55720 15000 1 0 $X=55605 $Y=13485
X18970 931 A[0] 2161 2476 1456 2321 2144 ICV_71 $T=58190 29000 1 0 $X=58075 $Y=27485
X18971 931 A[0] 1867 772 2480 2420 1087 ICV_71 $T=73960 26200 0 0 $X=73845 $Y=26085
X18986 93 95 931 A[0] 80 ICV_72 $T=8790 54200 0 180 $X=7915 $Y=52685
X18987 93 174 931 A[0] 126 ICV_72 $T=15060 68200 0 180 $X=14185 $Y=66685
X18988 93 219 931 A[0] 200 ICV_72 $T=18100 79400 1 180 $X=17225 $Y=79285
X18989 1077 B[21] 931 A[0] 2152 ICV_72 $T=60850 79400 0 180 $X=59975 $Y=77885
X18990 1077 A[21] 931 A[0] 1875 ICV_72 $T=66360 73800 0 180 $X=65485 $Y=72285
X18991 538 654 931 A[0] 578 ICV_72 $T=66930 57000 1 180 $X=66055 $Y=56885
X18992 538 683 931 A[0] 667 ICV_72 $T=69780 45800 0 180 $X=68905 $Y=44285
X18993 538 732 931 A[0] 720 ICV_72 $T=73960 48600 1 180 $X=73085 $Y=48485
X18994 931 A[0] 931 997 1294 ICV_73 $T=27790 20600 0 0 $X=27675 $Y=20485
X18995 931 A[0] 399 1056 304 ICV_73 $T=29120 29000 0 0 $X=29005 $Y=28885
X18996 931 A[0] 660 1011 1313 ICV_73 $T=32730 3800 1 0 $X=32615 $Y=2285
X18997 931 A[0] 506 965 1349 ICV_73 $T=38810 3800 1 0 $X=38695 $Y=2285
X18998 931 A[0] 428 338 2101 ICV_73 $T=45270 15000 0 0 $X=45155 $Y=14885
X18999 931 A[0] 392 338 494 ICV_73 $T=46600 59800 0 0 $X=46485 $Y=59685
X19000 931 A[0] 506 981 1409 ICV_73 $T=48880 37400 1 0 $X=48765 $Y=35885
X19001 931 A[0] 428 655 1441 ICV_73 $T=55910 17800 0 0 $X=55795 $Y=17685
X19002 931 A[0] 399 1020 2328 ICV_73 $T=62370 37400 0 0 $X=62255 $Y=37285
X19003 931 A[0] 660 338 646 ICV_73 $T=64460 43000 0 0 $X=64345 $Y=42885
X19004 931 A[0] 404 1011 1090 ICV_73 $T=73200 15000 1 0 $X=73085 $Y=13485
X19005 1863 989 931 A[0] INV_X8 $T=64270 59800 0 180 $X=62445 $Y=58285
X19006 1500 1015 931 A[0] INV_X8 $T=65410 54200 1 180 $X=63585 $Y=54085
X19007 2415 1024 931 A[0] INV_X8 $T=71110 31800 0 0 $X=70995 $Y=31685
X19008 2417 744 931 A[0] INV_X8 $T=71110 34600 0 0 $X=70995 $Y=34485
X19009 2478 1080 931 A[0] INV_X8 $T=72630 40200 1 0 $X=72515 $Y=38685
X19010 1896 404 931 A[0] INV_X8 $T=72630 51400 1 0 $X=72515 $Y=49885
X19026 404 A[0] 975 1681 931 110 1217 1681 2004 2245 931 ICV_75 $T=17340 15000 0 0 $X=17225 $Y=14885
X19027 744 A[0] 975 2001 931 1669 220 2380 2250 1680 931 ICV_75 $T=17340 26200 1 0 $X=17225 $Y=24685
X19028 1009 A[0] 1011 2063 931 2282 363 2459 2048 1991 931 ICV_75 $T=33680 29000 1 0 $X=33565 $Y=27485
X19029 392 A[0] 981 1330 931 358 366 2389 1740 1328 931 ICV_75 $T=33870 73800 1 0 $X=33755 $Y=72285
X19030 973 A[0] 965 1332 931 381 367 2458 2057 2064 931 ICV_75 $T=34250 37400 1 0 $X=34135 $Y=35885
X19031 319 A[0] 503 403 931 336 370 2062 1749 1320 931 ICV_75 $T=34440 76600 0 0 $X=34325 $Y=76485
X19032 448 A[0] 1025 415 931 1745 394 1344 1767 241 931 ICV_75 $T=36720 45800 1 0 $X=36605 $Y=44285
X19033 448 A[0] 995 2108 931 2395 461 2108 1400 478 931 ICV_75 $T=44510 65400 0 0 $X=44395 $Y=65285
X19034 1009 A[0] 965 2126 931 498 1819 1030 2315 2309 931 ICV_75 $T=50780 37400 0 0 $X=50665 $Y=37285
X19035 985 A[0] 997 1830 931 1418 517 1421 2318 2505 2528 ICV_75 $T=52490 1000 0 0 $X=52375 $Y=885
X19036 506 A[0] 503 534 931 516 1420 2490 2131 1432 931 ICV_75 $T=52870 29000 0 0 $X=52755 $Y=28885
X19037 1022 A[0] 965 2145 931 1827 526 1443 1072 411 931 ICV_75 $T=54770 34600 1 0 $X=54655 $Y=33085
X19038 258 A[0] 1014 2155 931 1837 2147 1460 1858 1851 931 ICV_75 $T=57240 45800 1 0 $X=57125 $Y=44285
X19039 1036 A[0] 965 2350 931 1086 1556 1911 1548 1547 931 ICV_75 $T=72060 12200 1 0 $X=71945 $Y=10685
X19051 1112 931 933 1943 A[0] NAND2_X1 $T=2140 31800 0 0 $X=2025 $Y=31685
X19052 936 931 13 24 A[0] NAND2_X1 $T=4800 43000 1 180 $X=4115 $Y=42885
X19053 938 931 1147 1132 A[0] NAND2_X1 $T=5560 43000 1 0 $X=5445 $Y=41485
X19054 1139 931 1145 53 A[0] NAND2_X1 $T=7080 31800 0 180 $X=6395 $Y=30285
X19055 939 931 1163 102 A[0] NAND2_X1 $T=7840 34600 1 0 $X=7725 $Y=33085
X19056 1160 931 1149 1163 A[0] NAND2_X1 $T=9170 31800 0 180 $X=8485 $Y=30285
X19057 1186 931 137 1187 A[0] NAND2_X1 $T=13920 48600 0 180 $X=13235 $Y=47085
X19058 172 931 1202 1191 A[0] NAND2_X1 $T=14490 54200 1 0 $X=14375 $Y=52685
X19059 1207 931 177 1662 A[0] NAND2_X1 $T=15440 59800 0 0 $X=15325 $Y=59685
X19060 1216 931 1213 211 A[0] NAND2_X1 $T=18290 62600 0 180 $X=17605 $Y=61085
X19061 212 931 1688 206 A[0] NAND2_X1 $T=17720 65400 0 0 $X=17605 $Y=65285
X19062 2040 931 2432 1671 A[0] NAND2_X1 $T=18100 79400 1 0 $X=17985 $Y=77885
X19063 223 931 1215 1219 A[0] NAND2_X1 $T=19810 54200 1 180 $X=19125 $Y=54085
X19064 224 931 221 152 A[0] NAND2_X1 $T=19620 57000 0 0 $X=19505 $Y=56885
X19065 230 931 1697 199 A[0] NAND2_X1 $T=20000 71000 1 0 $X=19885 $Y=69485
X19066 1233 931 1239 2252 A[0] NAND2_X1 $T=20570 76600 0 0 $X=20455 $Y=76485
X19067 1241 931 1994 1220 A[0] NAND2_X1 $T=21330 73800 1 0 $X=21215 $Y=72285
X19068 2009 931 274 2002 A[0] NAND2_X1 $T=24180 73800 1 180 $X=23495 $Y=73685
X19069 2026 931 993 2030 A[0] NAND2_X1 $T=26460 79400 0 0 $X=26345 $Y=79285
X19070 1285 931 319 993 A[0] NAND2_X1 $T=27410 79400 1 0 $X=27295 $Y=77885
X19071 2038 931 1741 2040 A[0] NAND2_X1 $T=30830 82200 0 0 $X=30715 $Y=82085
X19072 1536 931 2194 2416 A[0] NAND2_X1 $T=71300 71000 0 180 $X=70615 $Y=69485
X19073 1536 931 709 528 A[0] NAND2_X1 $T=71870 71000 0 180 $X=71185 $Y=69485
X19117 208 218 206 A[0] 199 2375 931 OAI211_X1 $T=17340 68200 1 0 $X=17225 $Y=66685
X19118 227 254 2002 A[0] 2252 2000 931 OAI211_X1 $T=20190 76600 1 0 $X=20075 $Y=75085
X19119 1847 504 1413 A[0] 508 488 931 OAI211_X1 $T=50970 12200 0 0 $X=50855 $Y=12085
X19120 1884 641 2175 A[0] 648 508 931 OAI211_X1 $T=65410 9400 1 0 $X=65295 $Y=7885
X19121 1078 643 659 A[0] 649 2175 931 OAI211_X1 $T=65600 6600 0 0 $X=65485 $Y=6485
X19122 2416 704 1552 A[0] 1551 1530 931 OAI211_X1 $T=70540 68200 1 0 $X=70425 $Y=66685
X19137 931 A[0] 1207 177 198 ICV_81 $T=16390 62600 0 180 $X=15705 $Y=61085
X19138 931 A[0] 973 1029 204 ICV_81 $T=19810 20600 0 180 $X=19125 $Y=19085
X19139 931 A[0] 976 931 1723 ICV_81 $T=28930 54200 1 180 $X=28245 $Y=54085
X19140 931 A[0] 1080 976 1728 ICV_81 $T=31400 15000 1 180 $X=30715 $Y=14885
X19141 931 A[0] 1022 997 2035 ICV_81 $T=32540 23400 0 180 $X=31855 $Y=21885
X19142 931 A[0] 664 995 1303 ICV_81 $T=33490 65400 1 180 $X=32805 $Y=65285
X19143 931 A[0] 973 986 2389 ICV_81 $T=36340 73800 1 180 $X=35655 $Y=73685
X19144 931 A[0] 506 1015 1035 ICV_81 $T=46980 31800 0 180 $X=46295 $Y=30285
X19145 931 A[0] 744 1009 2319 ICV_81 $T=56290 45800 0 180 $X=55605 $Y=44285
X19146 931 A[0] 1000 981 2325 ICV_81 $T=62940 54200 1 180 $X=62255 $Y=54085
X19147 931 A[0] 428 965 1885 ICV_81 $T=70350 17800 1 180 $X=69665 $Y=17685
X19148 931 A[0] 991 1014 1702 ICV_82 $T=24370 29000 0 0 $X=24255 $Y=28885
X19149 931 A[0] 392 997 1001 ICV_82 $T=29690 17800 0 0 $X=29575 $Y=17685
X19150 931 A[0] 2038 1741 1231 ICV_82 $T=30260 82200 1 0 $X=30145 $Y=80685
X19151 931 A[0] 1007 1012 375 ICV_82 $T=32920 34600 0 0 $X=32805 $Y=34485
X19152 931 A[0] 258 1015 2060 ICV_82 $T=36340 48600 1 0 $X=36225 $Y=47085
X19153 931 A[0] 258 965 407 ICV_82 $T=37670 20600 0 0 $X=37555 $Y=20485
X19154 931 A[0] 931 980 442 ICV_82 $T=43750 37400 1 0 $X=43635 $Y=35885
X19155 931 A[0] 931 995 1059 ICV_82 $T=54010 34600 0 0 $X=53895 $Y=34485
X19156 931 A[0] 506 980 556 ICV_82 $T=54010 54200 1 0 $X=53895 $Y=52685
X19157 931 A[0] 1015 1022 1439 ICV_82 $T=54390 71000 0 0 $X=54275 $Y=70885
X19158 931 A[0] 506 986 2142 ICV_82 $T=57430 48600 1 0 $X=57315 $Y=47085
X19159 931 A[0] 506 1011 2334 ICV_82 $T=68260 29000 0 0 $X=68145 $Y=28885
X19160 931 A[0] 1024 965 2190 ICV_82 $T=69590 23400 0 0 $X=69475 $Y=23285
X19161 931 A[0] 931 989 2013 ICV_83 $T=22660 17800 0 0 $X=22545 $Y=17685
X19162 931 A[0] 428 503 269 ICV_83 $T=22660 26200 0 0 $X=22545 $Y=26085
X19163 931 A[0] 991 503 1260 ICV_83 $T=23800 23400 0 0 $X=23685 $Y=23285
X19164 931 A[0] 664 983 1262 ICV_83 $T=23990 3800 1 0 $X=23875 $Y=2285
X19165 931 A[0] 1024 1014 1716 ICV_83 $T=26650 43000 0 0 $X=26535 $Y=42885
X19166 931 A[0] 319 980 313 ICV_83 $T=28170 71000 0 0 $X=28055 $Y=70885
X19167 931 A[0] 1007 1056 2269 ICV_83 $T=30450 20600 0 0 $X=30335 $Y=20485
X19168 931 A[0] 1000 655 2042 ICV_83 $T=31590 34600 1 0 $X=31475 $Y=33085
X19169 931 A[0] 660 965 1310 ICV_83 $T=33490 31800 0 0 $X=33375 $Y=31685
X19170 931 A[0] 989 931 385 ICV_83 $T=36150 71000 1 0 $X=36035 $Y=69485
X19171 931 A[0] 976 1007 2290 ICV_83 $T=39000 59800 1 0 $X=38885 $Y=58285
X19172 931 A[0] 660 997 1032 ICV_83 $T=43180 6600 1 0 $X=43065 $Y=5085
X19173 931 A[0] 980 392 451 ICV_83 $T=43750 79400 1 0 $X=43635 $Y=77885
X19174 931 A[0] 258 981 2301 ICV_83 $T=45650 31800 1 0 $X=45535 $Y=30285
X19175 931 A[0] 973 319 2304 ICV_83 $T=46220 79400 0 0 $X=46105 $Y=79285
X19176 931 A[0] 664 655 2398 ICV_83 $T=48120 20600 1 0 $X=48005 $Y=19085
X19177 931 A[0] 506 995 2119 ICV_83 $T=51730 54200 1 0 $X=51615 $Y=52685
X19178 931 A[0] 744 788 1471 ICV_83 $T=61230 23400 0 0 $X=61115 $Y=23285
X19179 931 A[0] 1036 655 1864 ICV_83 $T=63700 20600 0 0 $X=63585 $Y=20485
X19180 931 A[0] 1033 1011 1486 ICV_83 $T=64840 26200 0 0 $X=64725 $Y=26085
X19181 931 A[0] 991 1025 2414 ICV_83 $T=68450 23400 1 0 $X=68335 $Y=21885
X19212 931 2487 12 23 A[0] XNOR2_X1 $T=3470 34600 1 180 $X=2215 $Y=34485
X19213 931 2227 54 1612 A[0] XNOR2_X1 $T=4610 51400 1 0 $X=4495 $Y=49885
X19214 931 1971 103 115 A[0] XNOR2_X1 $T=10500 48600 0 180 $X=9245 $Y=47085
X19215 931 1649 130 144 A[0] XNOR2_X1 $T=12970 54200 1 180 $X=11715 $Y=54085
X19216 931 1193 134 163 A[0] XNOR2_X1 $T=14300 62600 1 180 $X=13045 $Y=62485
X19217 931 250 225 249 A[0] XNOR2_X1 $T=20190 82200 0 180 $X=18935 $Y=80685
X19218 931 1251 271 287 A[0] XNOR2_X1 $T=23420 79400 1 180 $X=22165 $Y=79285
X19219 931 2026 295 307 A[0] XNOR2_X1 $T=26080 82200 0 180 $X=24825 $Y=80685
X19220 931 747 2148 543 A[0] XNOR2_X1 $T=57050 76600 0 0 $X=56935 $Y=76485
X19221 931 1503 2477 653 A[0] XNOR2_X1 $T=65980 73800 0 0 $X=65865 $Y=73685
X19222 931 1888 1518 2477 A[0] XNOR2_X1 $T=67690 73800 1 0 $X=67575 $Y=72285
X19223 931 A[0] 2444 71 1615 1946 1968 ICV_86 $T=5940 26200 0 0 $X=5825 $Y=26085
X19224 931 A[0] 1685 272 1257 1258 2011 ICV_86 $T=21710 54200 1 0 $X=21595 $Y=52685
X19225 931 A[0] 306 313 1288 1304 1722 ICV_86 $T=25510 73800 1 0 $X=25395 $Y=72285
X19226 931 A[0] 1366 437 2399 2093 1377 ICV_86 $T=42040 59800 0 0 $X=41925 $Y=59685
X19227 931 A[0] 421 467 1391 1405 1039 ICV_86 $T=45270 12200 1 0 $X=45155 $Y=10685
X19228 931 A[0] 2497 593 1484 2171 1072 ICV_86 $T=61230 29000 0 0 $X=61115 $Y=28885
X19229 931 A[0] 1424 645 1081 1870 1515 ICV_86 $T=65410 34600 1 0 $X=65295 $Y=33085
X19230 931 A[0] 2184 673 2191 1086 1887 ICV_86 $T=67690 3800 0 0 $X=67575 $Y=3685
X19231 448 A[0] 1012 2247 931 258 338 1217 ICV_87 $T=17720 17800 1 0 $X=17605 $Y=16285
X19232 448 A[0] 965 2257 931 660 1012 2378 ICV_87 $T=22280 34600 0 0 $X=22165 $Y=34485
X19233 1024 A[0] 986 1677 931 1080 503 1692 ICV_87 $T=22280 43000 1 0 $X=22165 $Y=41485
X19234 1080 A[0] 981 2016 931 1024 503 2258 ICV_87 $T=26650 29000 0 0 $X=26535 $Y=28885
X19235 975 A[0] 931 2041 931 1000 980 349 ICV_87 $T=31590 62600 1 0 $X=31475 $Y=61085
X19236 931 A[0] 983 377 931 399 1029 1334 ICV_87 $T=36910 29000 0 0 $X=36795 $Y=28885
X19237 164 A[0] 1022 2482 931 655 931 2483 ICV_87 $T=37670 48600 0 0 $X=37555 $Y=48485
X19238 931 A[0] 164 396 931 404 1020 1356 ICV_87 $T=38430 20600 1 0 $X=38315 $Y=19085
X19239 1024 A[0] 995 1347 931 428 1009 1758 ICV_87 $T=39190 31800 0 0 $X=39075 $Y=31685
X19240 1022 A[0] 983 408 931 931 1029 1026 ICV_87 $T=39380 23400 0 0 $X=39265 $Y=23285
X19241 1033 A[0] 788 457 931 506 1012 1380 ICV_87 $T=43940 20600 0 0 $X=43825 $Y=20485
X19242 399 A[0] 1014 2117 931 986 931 2107 ICV_87 $T=49640 79400 1 0 $X=49525 $Y=77885
X19243 985 A[0] 503 515 931 1000 986 1425 ICV_87 $T=52300 62600 0 0 $X=52185 $Y=62485
X19244 664 A[0] 338 1420 931 985 975 2490 ICV_87 $T=53060 31800 1 0 $X=52945 $Y=30285
X19245 258 A[0] 980 2485 931 404 995 1428 ICV_87 $T=54010 43000 0 0 $X=53895 $Y=42885
X19246 973 A[0] 1014 1427 931 1007 986 1429 ICV_87 $T=54390 71000 1 0 $X=54275 $Y=69485
X19247 399 A[0] 164 1461 931 392 655 2151 ICV_87 $T=58950 48600 0 0 $X=58835 $Y=48485
X19248 660 A[0] 976 594 931 973 975 2165 ICV_87 $T=60470 57000 1 0 $X=60355 $Y=55485
X19249 501 A[0] 1015 1484 931 931 1012 2172 ICV_87 $T=63130 31800 1 0 $X=63015 $Y=30285
X19250 985 A[0] 989 2408 931 501 981 2409 ICV_87 $T=63130 45800 0 0 $X=63015 $Y=45685
X19251 1024 A[0] 1025 2170 931 1080 1020 1487 ICV_87 $T=63510 6600 1 0 $X=63395 $Y=5085
X19252 404 A[0] 788 1507 931 744 1012 2338 ICV_87 $T=66550 3800 0 0 $X=66435 $Y=3685
X19253 302 A[0] 292 1265 931 1283 306 1284 2034 1703 ICV_88 $T=24940 76600 0 180 $X=24255 $Y=75085
X19254 744 A[0] 981 2021 931 1276 316 1293 2267 318 ICV_88 $T=26460 45800 0 180 $X=25775 $Y=44285
X19255 975 A[0] 319 2022 931 2020 325 2494 2268 341 ICV_88 $T=27600 65400 0 180 $X=26915 $Y=63885
X19256 448 A[0] 1011 2292 931 1371 2470 2099 1388 1386 ICV_88 $T=43560 6600 1 180 $X=42875 $Y=6485
X19257 448 A[0] 164 1395 931 481 489 1053 2313 559 ICV_88 $T=48690 20600 1 180 $X=48005 $Y=20485
X19258 744 A[0] 1014 2397 931 2308 490 1816 1432 1812 ICV_88 $T=48690 31800 0 180 $X=48005 $Y=30285
X19259 664 A[0] 319 1400 931 1402 2474 2120 2124 1813 ICV_88 $T=48690 65400 1 180 $X=48005 $Y=65285
X19260 1007 A[0] 965 1398 931 2471 497 1414 1055 1818 ICV_88 $T=49450 26200 0 180 $X=48765 $Y=24685
X19261 503 A[0] 931 2400 931 1811 2400 1423 1430 1825 ICV_88 $T=51350 79400 0 180 $X=50665 $Y=77885
X19262 1033 A[0] 981 2171 931 627 628 1505 2334 1876 ICV_88 $T=64270 29000 0 180 $X=63585 $Y=27485
X19263 991 A[0] 164 1481 931 605 650 2414 2339 1881 ICV_88 $T=65790 20600 0 180 $X=65105 $Y=19085
X19279 931 A[0] 2250 110 1640 1633 1978 ICV_90 $T=8980 17800 0 0 $X=8865 $Y=17685
X19280 931 A[0] 229 195 1214 964 196 ICV_90 $T=15630 29000 1 0 $X=15515 $Y=27485
X19281 931 A[0] 1222 235 2005 2253 2236 ICV_90 $T=18670 20600 0 0 $X=18555 $Y=20485
X19282 931 A[0] 285 1701 1238 2256 1687 ICV_90 $T=18670 65400 1 0 $X=18555 $Y=63885
X19283 931 A[0] 230 246 1229 1715 1688 ICV_90 $T=18670 68200 0 0 $X=18555 $Y=68085
X19284 931 A[0] 1241 265 2377 1698 1697 ICV_90 $T=20760 71000 0 0 $X=20645 $Y=70885
X19285 931 A[0] 173 312 1712 2265 1290 ICV_90 $T=25320 3800 0 0 $X=25205 $Y=3685
X19286 931 A[0] 1031 324 1298 2455 294 ICV_90 $T=27220 71000 1 0 $X=27105 $Y=69485
X19287 931 A[0] 2455 331 1303 2272 1306 ICV_90 $T=28360 68200 1 0 $X=28245 $Y=66685
X19288 931 A[0] 298 347 1317 2278 376 ICV_90 $T=31780 15000 1 0 $X=31665 $Y=13485
X19289 931 A[0] 312 1343 1340 1747 1017 ICV_90 $T=34630 3800 0 0 $X=34515 $Y=3685
X19290 931 A[0] 1742 382 1337 2287 146 ICV_90 $T=35580 43000 1 0 $X=35465 $Y=41485
X19291 931 A[0] 1324 383 1748 1342 339 ICV_90 $T=35580 43000 0 0 $X=35465 $Y=42885
X19292 931 A[0] 998 384 1338 2288 1752 ICV_90 $T=35580 57000 1 0 $X=35465 $Y=55485
X19293 931 A[0] 2278 387 1756 2289 2073 ICV_90 $T=35770 12200 0 0 $X=35655 $Y=12085
X19294 931 A[0] 389 391 2069 1329 1297 ICV_90 $T=36150 23400 0 0 $X=36035 $Y=23285
X19295 931 A[0] 370 403 1353 2484 1760 ICV_90 $T=38050 79400 1 0 $X=37935 $Y=77885
X19296 931 A[0] 2394 407 1356 2071 1764 ICV_90 $T=38620 23400 1 0 $X=38505 $Y=21885
X19297 931 A[0] 2256 416 1771 1351 1770 ICV_90 $T=38620 65400 0 0 $X=38505 $Y=65285
X19298 931 A[0] 2061 417 1361 2294 1771 ICV_90 $T=38620 68200 1 0 $X=38505 $Y=66685
X19299 931 A[0] 2283 419 2080 1369 1772 ICV_90 $T=38620 79400 0 0 $X=38505 $Y=79285
X19300 931 A[0] 511 484 1039 2132 507 ICV_90 $T=47930 9400 1 0 $X=47815 $Y=7885
X19301 931 A[0] 499 498 1829 1808 1044 ICV_90 $T=49450 45800 1 0 $X=49335 $Y=44285
X19302 931 A[0] 520 521 1437 1435 1422 ICV_90 $T=53630 12200 1 0 $X=53515 $Y=10685
X19303 931 A[0] 2129 523 2137 1062 1054 ICV_90 $T=54010 48600 0 0 $X=53895 $Y=48485
X19304 931 A[0] 2134 535 1451 2146 1455 ICV_90 $T=55720 65400 1 0 $X=55605 $Y=63885
X19305 931 A[0] 1061 546 559 1843 1849 ICV_90 $T=56860 20600 1 0 $X=56745 $Y=19085
X19306 931 A[0] 1062 2496 2150 1851 1850 ICV_90 $T=57050 43000 0 0 $X=56935 $Y=42885
X19307 931 A[0] 539 560 2158 2157 504 ICV_90 $T=58760 9400 0 0 $X=58645 $Y=9285
X19308 931 A[0] 2158 581 2411 931 602 ICV_90 $T=60280 12200 1 0 $X=60165 $Y=10685
X19309 931 A[0] 653 630 1898 2336 2183 ICV_90 $T=64270 76600 1 0 $X=64155 $Y=75085
X19350 2229 1625 1952 2223 A[0] 931 19 931 ICV_91 $T=1000 3800 0 0 $X=885 $Y=3685
X19351 20 19 1126 2225 A[0] 931 18 931 ICV_91 $T=2330 15000 1 0 $X=2215 $Y=13485
X19352 2369 101 1178 2236 A[0] 931 86 931 ICV_91 $T=8410 12200 1 0 $X=8295 $Y=10685
X19353 156 171 1206 2243 A[0] 931 1210 931 ICV_91 $T=13920 43000 1 0 $X=13805 $Y=41485
X19354 279 280 1713 1711 A[0] 931 1705 931 ICV_91 $T=22280 40200 0 0 $X=22165 $Y=40085
X19355 2024 318 2032 1315 A[0] 931 999 931 ICV_91 $T=26460 34600 0 0 $X=26345 $Y=34485
X19356 1774 434 1371 1370 A[0] 931 1780 931 ICV_91 $T=41850 9400 1 0 $X=41735 $Y=7885
X19357 1358 436 1812 453 A[0] 931 1781 931 ICV_91 $T=41850 40200 0 0 $X=41735 $Y=40085
X19358 2466 446 1379 2302 A[0] 931 425 931 ICV_91 $T=42230 76600 1 0 $X=42115 $Y=75085
X19359 1779 455 1386 1822 A[0] 931 475 931 ICV_91 $T=43940 6600 1 0 $X=43825 $Y=5085
X19360 2468 463 1802 1403 A[0] 931 1038 2528 ICV_91 $T=44700 1000 0 0 $X=44585 $Y=885
X19361 454 470 2473 1810 A[0] 931 1799 931 ICV_91 $T=45270 54200 1 0 $X=45155 $Y=52685
X19362 1796 478 1426 1813 A[0] 931 1805 931 ICV_91 $T=46220 68200 1 0 $X=46105 $Y=66685
X19363 563 605 1493 1867 A[0] 931 1075 931 ICV_91 $T=62370 23400 1 0 $X=62255 $Y=21885
X19364 1858 2408 1495 2409 A[0] 931 1871 931 ICV_91 $T=62370 45800 1 0 $X=62255 $Y=44285
X19365 931 A[0] 1944 15 1131 1117 1958 ICV_92 $T=1950 3800 1 0 $X=1835 $Y=2285
X19366 931 A[0] 1601 17 2369 1944 40 ICV_92 $T=1950 9400 0 0 $X=1835 $Y=9285
X19367 931 A[0] 1114 18 1125 1630 1143 ICV_92 $T=1950 12200 1 0 $X=1835 $Y=10685
X19368 931 A[0] 1946 20 1945 42 1614 ICV_92 $T=1950 15000 0 0 $X=1835 $Y=14885
X19369 931 A[0] 1111 21 1614 1959 1127 ICV_92 $T=1950 17800 1 0 $X=1835 $Y=16285
X19370 931 A[0] 1106 2442 1135 2226 1615 ICV_92 $T=1950 23400 0 0 $X=1835 $Y=23285
X19371 931 A[0] 300 281 1250 1276 1706 ICV_92 $T=21900 45800 1 0 $X=21785 $Y=44285
X19372 931 A[0] 1234 282 1016 1261 2019 ICV_92 $T=21900 48600 0 0 $X=21785 $Y=48485
X19373 931 A[0] 267 283 2014 1312 1707 ICV_92 $T=21900 59800 1 0 $X=21785 $Y=58285
X19374 931 A[0] 321 284 1259 1273 1708 ICV_92 $T=21900 62600 0 0 $X=21785 $Y=62485
X19375 931 A[0] 2377 285 1805 2047 246 ICV_92 $T=21900 68200 0 0 $X=21785 $Y=68085
X19376 931 A[0] 335 438 1374 2297 1052 ICV_92 $T=41850 12200 1 0 $X=41735 $Y=10685
X19377 931 A[0] 422 439 2089 2299 1783 ICV_92 $T=41850 15000 0 0 $X=41735 $Y=14885
X19378 931 A[0] 1777 A[0] 457 1380 439 ICV_92 $T=41850 20600 1 0 $X=41735 $Y=19085
X19379 931 A[0] 441 442 1387 2102 2488 ICV_92 $T=41850 37400 0 0 $X=41735 $Y=37285
X19380 931 A[0] 1392 443 1375 1323 1786 ICV_92 $T=41850 40200 1 0 $X=41735 $Y=38685
X19381 931 A[0] 2465 444 1054 1788 1383 ICV_92 $T=41850 48600 1 0 $X=41735 $Y=47085
X19382 931 A[0] 223 1789 1376 1776 2095 ICV_92 $T=41850 54200 1 0 $X=41735 $Y=52685
X19383 931 A[0] 2045 2097 1397 1790 1789 ICV_92 $T=41850 57000 0 0 $X=41735 $Y=56885
X19384 931 A[0] 2323 604 1492 1510 1868 ICV_92 $T=61990 17800 1 0 $X=61875 $Y=16285
X19385 931 A[0] 931 606 1866 627 1869 ICV_92 $T=61990 23400 0 0 $X=61875 $Y=23285
X19386 931 A[0] 2329 607 1494 2328 1444 ICV_92 $T=61990 37400 1 0 $X=61875 $Y=35885
X19387 931 A[0] 2496 609 1871 2186 1497 ICV_92 $T=61990 43000 1 0 $X=61875 $Y=41485
X19388 931 A[0] 2168 611 1496 1872 1873 ICV_92 $T=61990 51400 1 0 $X=61875 $Y=49885
X19389 931 A[0] 1859 931 1088 2330 1478 ICV_92 $T=61990 79400 0 0 $X=61875 $Y=79285
X19406 931 A[0] 1033 1658 655 ICV_93 $T=15060 20600 1 180 $X=14375 $Y=20485
X19407 931 A[0] 1080 1274 986 ICV_93 $T=27980 43000 1 180 $X=27295 $Y=42885
X19408 931 A[0] 973 2268 981 ICV_93 $T=31780 65400 1 180 $X=31095 $Y=65285
X19409 931 A[0] 1022 2069 1011 ICV_93 $T=37480 23400 0 180 $X=36795 $Y=21885
X19410 931 A[0] 985 1372 1056 ICV_93 $T=44510 15000 0 180 $X=43825 $Y=13485
X19411 931 A[0] 1036 1389 989 ICV_93 $T=46980 20600 0 180 $X=46295 $Y=19085
X19412 931 A[0] 980 472 973 ICV_93 $T=48690 71000 1 180 $X=48005 $Y=70885
X19413 931 A[0] 404 1454 1014 ICV_93 $T=58950 31800 1 180 $X=58265 $Y=31685
X19414 931 A[0] 1009 2154 788 ICV_93 $T=60660 31800 1 180 $X=59975 $Y=31685
X19415 1135 60 1653 1650 A[0] 931 1966 ICV_94 $T=5370 23400 0 0 $X=5255 $Y=23285
X19416 1980 149 1678 1244 A[0] 931 1660 ICV_94 $T=12210 45800 0 0 $X=12095 $Y=45685
X19417 243 255 2011 1708 A[0] 931 2014 ICV_94 $T=20190 57000 0 0 $X=20075 $Y=56885
X19418 977 268 1253 1019 A[0] 931 1700 ICV_94 $T=21520 12200 1 0 $X=21405 $Y=10685
X19419 262 2387 1268 998 A[0] 931 261 ICV_94 $T=26080 57000 1 0 $X=25965 $Y=55485
X19420 356 357 1745 2064 A[0] 931 2056 ICV_94 $T=32730 40200 0 0 $X=32615 $Y=40085
X19421 1326 393 2482 2483 A[0] 931 1359 ICV_94 $T=36530 51400 1 0 $X=36415 $Y=49885
X19422 513 2144 1037 2463 A[0] 931 468 ICV_94 $T=44700 29000 1 0 $X=44585 $Y=27485
X19423 1822 1844 1434 1833 A[0] 931 548 ICV_94 $T=53630 6600 1 0 $X=53515 $Y=5085
X19424 1828 1514 1444 2161 A[0] 931 1839 ICV_94 $T=54770 40200 1 0 $X=54655 $Y=38685
X19429 A[0] 2235 14 1602 931 XOR2_X1 $T=1000 45800 0 0 $X=885 $Y=45685
X19430 A[0] 2447 95 2500 931 XOR2_X1 $T=9170 51400 1 180 $X=7915 $Y=51285
X19431 A[0] 154 125 1673 931 XOR2_X1 $T=12780 57000 1 180 $X=11525 $Y=56885
X19432 A[0] 954 118 2372 931 XOR2_X1 $T=13160 62600 0 180 $X=11905 $Y=61085
X19433 A[0] 1651 123 2449 931 XOR2_X1 $T=13920 59800 0 180 $X=12665 $Y=58285
X19434 A[0] 2012 1654 1656 931 XOR2_X1 $T=15440 79400 1 180 $X=14185 $Y=79285
X19435 A[0] 1248 180 1211 931 XOR2_X1 $T=16770 73800 1 180 $X=15515 $Y=73685
X19436 A[0] 208 186 1666 931 XOR2_X1 $T=17150 65400 0 180 $X=15895 $Y=63885
X19437 A[0] 2244 174 2450 931 XOR2_X1 $T=17340 68200 0 180 $X=16085 $Y=66685
X19438 A[0] 231 178 1996 931 XOR2_X1 $T=18670 76600 1 180 $X=17415 $Y=76485
X19439 A[0] 227 209 1228 931 XOR2_X1 $T=19050 76600 1 0 $X=18935 $Y=75085
X19442 203 A[0] 1987 1657 215 1661 931 AOI211_X2 $T=17340 15000 0 180 $X=15515 $Y=13485
X19443 273 A[0] 2376 972 227 2375 931 AOI211_X2 $T=20380 73800 1 180 $X=18555 $Y=73685
X19444 11 1949 1107 931 A[0] XOR2_X2 $T=1000 37400 1 0 $X=885 $Y=35885
X19445 10 2368 1123 931 A[0] XOR2_X2 $T=4610 51400 0 180 $X=2785 $Y=49885
X19446 65 2443 935 931 A[0] XOR2_X2 $T=4800 48600 0 0 $X=4685 $Y=48485
X19447 179 1208 1212 931 A[0] XOR2_X2 $T=17340 71000 1 180 $X=15515 $Y=70885
X19448 219 276 1671 931 A[0] XOR2_X2 $T=18100 79400 0 180 $X=16275 $Y=77885
X19449 1600 A[0] 24 1123 2235 931 AOI21_X2 $T=2140 45800 0 0 $X=2025 $Y=45685
X19450 1146 A[0] 38 1177 1158 931 AOI21_X2 $T=7080 34600 0 0 $X=6965 $Y=34485
X19451 1203 A[0] 1200 208 185 931 AOI21_X2 $T=14870 57000 1 0 $X=14755 $Y=55485
X19452 1112 937 933 931 A[0] NOR2_X2 $T=1950 34600 0 180 $X=885 $Y=33085
X19453 1147 1128 938 931 A[0] NOR2_X2 $T=4610 43000 1 0 $X=4495 $Y=41485
X19454 38 64 1158 931 A[0] NOR2_X2 $T=4800 34600 0 0 $X=4685 $Y=34485
X19455 176 1987 1199 931 A[0] NOR2_X2 $T=15630 15000 1 180 $X=14565 $Y=14885
X19456 91 94 A[0] 2445 133 61 48 931 AOI221_X2 $T=7460 45800 0 0 $X=7345 $Y=45685
X19457 175 215 A[0] 183 148 176 1199 931 AOI221_X2 $T=15630 15000 0 180 $X=13425 $Y=13485
X19458 528 543 2342 56 A[0] 931 NOR3_X4 $T=15630 68200 1 180 $X=12855 $Y=68085
X19459 157 2342 528 934 A[0] 931 NOR3_X4 $T=12970 71000 1 0 $X=12855 $Y=69485
X19460 93 104 1002 931 A[0] NAND2_X2 $T=7650 82200 0 0 $X=7535 $Y=82085
X19461 155 953 148 931 A[0] NAND2_X2 $T=13920 31800 1 180 $X=12855 $Y=31685
.ENDS
***************************************
