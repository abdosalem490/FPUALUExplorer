/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 16 23:21:39 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 219466199 */

module datapath(A_in, p_0);
   input [31:0]A_in;
   output [31:0]p_0;

   AOI21_X1 i_2 (.A(n_58), .B1(A_in[3]), .B2(n_59), .ZN(p_0[3]));
   AOI21_X1 i_6 (.A(n_55), .B1(A_in[7]), .B2(n_0), .ZN(p_0[7]));
   INV_X1 i_7 (.A(n_1), .ZN(n_0));
   AOI21_X1 i_16 (.A(n_52), .B1(A_in[11]), .B2(n_6), .ZN(p_0[11]));
   INV_X1 i_17 (.A(n_7), .ZN(n_6));
   AOI21_X1 i_23 (.A(n_17), .B1(A_in[12]), .B2(n_51), .ZN(p_0[12]));
   AOI21_X1 i_25 (.A(n_13), .B1(A_in[14]), .B2(n_14), .ZN(p_0[14]));
   AOI21_X1 i_26 (.A(n_49), .B1(A_in[15]), .B2(n_12), .ZN(p_0[15]));
   INV_X1 i_27 (.A(n_13), .ZN(n_12));
   NOR2_X1 i_28 (.A1(n_51), .A2(n_50), .ZN(n_13));
   INV_X1 i_29 (.A(n_15), .ZN(n_14));
   AOI21_X1 i_33 (.A(n_23), .B1(A_in[16]), .B2(n_48), .ZN(p_0[16]));
   AOI21_X1 i_35 (.A(n_19), .B1(A_in[18]), .B2(n_20), .ZN(p_0[18]));
   AOI21_X1 i_36 (.A(n_45), .B1(A_in[19]), .B2(n_18), .ZN(p_0[19]));
   INV_X1 i_37 (.A(n_19), .ZN(n_18));
   NOR2_X1 i_38 (.A1(n_48), .A2(n_46), .ZN(n_19));
   INV_X1 i_39 (.A(n_21), .ZN(n_20));
   AOI21_X1 i_43 (.A(n_25), .B1(A_in[20]), .B2(n_44), .ZN(p_0[20]));
   AOI21_X1 i_44 (.A(n_27), .B1(A_in[21]), .B2(n_24), .ZN(p_0[21]));
   INV_X1 i_45 (.A(n_25), .ZN(n_24));
   NOR2_X1 i_46 (.A1(A_in[20]), .A2(n_44), .ZN(n_25));
   AOI21_X1 i_47 (.A(n_43), .B1(A_in[22]), .B2(n_26), .ZN(p_0[22]));
   INV_X1 i_48 (.A(n_27), .ZN(n_26));
   NOR3_X1 i_49 (.A1(A_in[21]), .A2(A_in[20]), .A3(n_44), .ZN(n_27));
   AOI21_X1 i_50 (.A(n_41), .B1(A_in[23]), .B2(n_42), .ZN(p_0[23]));
   AOI21_X1 i_51 (.A(n_29), .B1(A_in[24]), .B2(n_40), .ZN(p_0[24]));
   AOI21_X1 i_55 (.A(n_32), .B1(A_in[26]), .B2(n_30), .ZN(p_0[26]));
   AOI21_X1 i_57 (.A(n_39), .B1(A_in[27]), .B2(n_31), .ZN(p_0[27]));
   INV_X1 i_58 (.A(n_32), .ZN(n_31));
   NOR2_X1 i_59 (.A1(n_47), .A2(n_40), .ZN(n_32));
   AOI21_X1 i_60 (.A(n_34), .B1(A_in[28]), .B2(n_38), .ZN(p_0[28]));
   AOI21_X1 i_61 (.A(n_36), .B1(A_in[29]), .B2(n_33), .ZN(p_0[29]));
   INV_X1 i_62 (.A(n_34), .ZN(n_33));
   NOR2_X1 i_63 (.A1(A_in[28]), .A2(n_38), .ZN(n_34));
   AOI21_X1 i_64 (.A(n_37), .B1(A_in[30]), .B2(n_35), .ZN(p_0[30]));
   INV_X1 i_65 (.A(n_36), .ZN(n_35));
   NOR3_X1 i_66 (.A1(A_in[29]), .A2(A_in[28]), .A3(n_38), .ZN(n_36));
   XNOR2_X1 i_67 (.A(A_in[31]), .B(n_37), .ZN(p_0[31]));
   NOR4_X1 i_68 (.A1(A_in[29]), .A2(A_in[28]), .A3(A_in[30]), .A4(n_38), 
      .ZN(n_37));
   INV_X1 i_69 (.A(n_39), .ZN(n_38));
   NOR3_X1 i_70 (.A1(A_in[27]), .A2(n_47), .A3(n_40), .ZN(n_39));
   OR3_X1 i_78 (.A1(A_in[26]), .A2(A_in[25]), .A3(A_in[24]), .ZN(n_47));
   NOR2_X1 i_0 (.A1(n_40), .A2(A_in[24]), .ZN(n_29));
   INV_X1 i_1 (.A(n_42), .ZN(n_43));
   NAND2_X1 i_3 (.A1(n_45), .A2(n_10), .ZN(n_42));
   INV_X1 i_4 (.A(n_45), .ZN(n_44));
   NOR2_X1 i_5 (.A1(n_48), .A2(n_22), .ZN(n_45));
   NAND3_X1 i_8 (.A1(n_62), .A2(n_66), .A3(n_63), .ZN(n_50));
   NOR2_X1 i_9 (.A1(n_94), .A2(A_in[13]), .ZN(n_15));
   INV_X1 i_10 (.A(n_94), .ZN(n_17));
   INV_X1 i_12 (.A(n_2), .ZN(p_0[9]));
   NAND2_X1 i_13 (.A1(n_86), .A2(n_3), .ZN(n_2));
   NAND2_X1 i_14 (.A1(n_85), .A2(A_in[9]), .ZN(n_3));
   NOR2_X1 i_15 (.A1(n_4), .A2(n_21), .ZN(p_0[17]));
   NOR2_X1 i_18 (.A1(n_23), .A2(n_54), .ZN(n_4));
   INV_X1 i_19 (.A(n_5), .ZN(n_21));
   NAND2_X1 i_20 (.A1(n_23), .A2(n_54), .ZN(n_5));
   NOR2_X1 i_21 (.A1(n_48), .A2(A_in[16]), .ZN(n_23));
   NOR2_X1 i_22 (.A1(n_9), .A2(n_8), .ZN(p_0[25]));
   INV_X1 i_24 (.A(n_30), .ZN(n_8));
   NAND3_X1 i_30 (.A1(n_41), .A2(n_71), .A3(n_70), .ZN(n_30));
   AOI21_X1 i_31 (.A(n_71), .B1(n_41), .B2(n_70), .ZN(n_9));
   INV_X1 i_32 (.A(n_40), .ZN(n_41));
   NAND4_X1 i_34 (.A1(n_49), .A2(n_69), .A3(n_16), .A4(n_10), .ZN(n_40));
   INV_X1 i_40 (.A(n_11), .ZN(n_10));
   OR3_X1 i_41 (.A1(A_in[20]), .A2(A_in[21]), .A3(A_in[22]), .ZN(n_11));
   INV_X1 i_42 (.A(n_22), .ZN(n_16));
   OR2_X1 i_52 (.A1(n_46), .A2(A_in[19]), .ZN(n_22));
   NAND3_X1 i_53 (.A1(n_54), .A2(n_28), .A3(n_56), .ZN(n_46));
   INV_X1 i_54 (.A(A_in[16]), .ZN(n_28));
   INV_X1 i_56 (.A(A_in[17]), .ZN(n_54));
   INV_X1 i_71 (.A(A_in[18]), .ZN(n_56));
   INV_X1 i_72 (.A(n_48), .ZN(n_49));
   NAND4_X1 i_73 (.A1(n_58), .A2(n_68), .A3(n_53), .A4(n_60), .ZN(n_48));
   INV_X1 i_74 (.A(n_61), .ZN(n_60));
   NAND4_X1 i_75 (.A1(n_62), .A2(n_66), .A3(n_64), .A4(n_63), .ZN(n_61));
   INV_X1 i_76 (.A(A_in[13]), .ZN(n_62));
   INV_X1 i_77 (.A(A_in[14]), .ZN(n_63));
   INV_X1 i_79 (.A(A_in[15]), .ZN(n_64));
   NAND4_X1 i_80 (.A1(n_90), .A2(n_88), .A3(n_67), .A4(n_103), .ZN(n_65));
   INV_X1 i_82 (.A(A_in[11]), .ZN(n_67));
   INV_X1 i_83 (.A(n_96), .ZN(n_68));
   INV_X1 i_84 (.A(n_57), .ZN(n_58));
   INV_X1 i_85 (.A(A_in[23]), .ZN(n_69));
   INV_X1 i_86 (.A(A_in[24]), .ZN(n_70));
   INV_X1 i_87 (.A(A_in[25]), .ZN(n_71));
   NAND3_X1 i_11 (.A1(n_97), .A2(n_99), .A3(n_98), .ZN(n_72));
   INV_X1 i_92 (.A(n_75), .ZN(p_0[2]));
   NAND2_X1 i_93 (.A1(n_76), .A2(n_59), .ZN(n_75));
   NAND2_X1 i_94 (.A1(n_74), .A2(A_in[2]), .ZN(n_76));
   NAND3_X1 i_96 (.A1(n_77), .A2(n_104), .A3(n_84), .ZN(n_59));
   INV_X1 i_97 (.A(n_78), .ZN(p_0[4]));
   XNOR2_X1 i_98 (.A(n_57), .B(A_in[4]), .ZN(n_78));
   NOR2_X1 i_99 (.A1(n_79), .A2(n_80), .ZN(p_0[5]));
   AOI21_X1 i_100 (.A(n_98), .B1(n_82), .B2(n_83), .ZN(n_79));
   INV_X1 i_101 (.A(n_81), .ZN(n_80));
   AOI21_X1 i_102 (.A(n_1), .B1(n_81), .B2(A_in[6]), .ZN(p_0[6]));
   NAND3_X1 i_103 (.A1(n_82), .A2(n_98), .A3(n_83), .ZN(n_81));
   INV_X1 i_104 (.A(n_57), .ZN(n_82));
   INV_X1 i_105 (.A(A_in[4]), .ZN(n_83));
   NOR2_X1 i_106 (.A1(n_57), .A2(n_72), .ZN(n_1));
   INV_X1 i_108 (.A(n_101), .ZN(n_57));
   NAND2_X1 i_109 (.A1(n_55), .A2(n_88), .ZN(n_85));
   INV_X1 i_110 (.A(n_52), .ZN(n_51));
   NOR2_X1 i_111 (.A1(n_92), .A2(n_65), .ZN(n_52));
   XNOR2_X1 i_112 (.A(n_92), .B(n_88), .ZN(p_0[8]));
   AOI21_X1 i_113 (.A(n_7), .B1(A_in[10]), .B2(n_86), .ZN(p_0[10]));
   NAND4_X1 i_114 (.A1(n_101), .A2(n_90), .A3(n_88), .A4(n_95), .ZN(n_86));
   INV_X1 i_117 (.A(n_89), .ZN(n_7));
   NAND2_X1 i_118 (.A1(n_55), .A2(n_87), .ZN(n_89));
   NAND2_X1 i_120 (.A1(n_93), .A2(n_91), .ZN(p_0[13]));
   NAND4_X1 i_121 (.A1(n_55), .A2(A_in[13]), .A3(n_66), .A4(n_53), .ZN(n_91));
   INV_X1 i_122 (.A(n_92), .ZN(n_55));
   NAND2_X1 i_123 (.A1(n_101), .A2(n_95), .ZN(n_92));
   NAND2_X1 i_124 (.A1(n_94), .A2(n_73), .ZN(n_93));
   NAND4_X1 i_125 (.A1(n_53), .A2(n_66), .A3(n_101), .A4(n_95), .ZN(n_94));
   INV_X1 i_81 (.A(n_96), .ZN(n_95));
   NAND4_X1 i_88 (.A1(n_97), .A2(n_100), .A3(n_99), .A4(n_98), .ZN(n_96));
   INV_X1 i_89 (.A(A_in[4]), .ZN(n_97));
   INV_X1 i_90 (.A(A_in[5]), .ZN(n_98));
   INV_X1 i_91 (.A(A_in[6]), .ZN(n_99));
   INV_X1 i_95 (.A(A_in[7]), .ZN(n_100));
   NOR2_X1 i_132 (.A1(n_102), .A2(A_in[0]), .ZN(n_101));
   NAND3_X1 i_133 (.A1(n_105), .A2(n_104), .A3(n_84), .ZN(n_102));
   INV_X1 i_135 (.A(A_in[2]), .ZN(n_104));
   INV_X1 i_136 (.A(A_in[3]), .ZN(n_105));
   INV_X1 i_137 (.A(n_65), .ZN(n_53));
   INV_X1 i_138 (.A(A_in[12]), .ZN(n_66));
   INV_X1 i_139 (.A(A_in[13]), .ZN(n_73));
   AOI22_X1 i_107 (.A1(n_84), .A2(n_77), .B1(A_in[1]), .B2(A_in[0]), .ZN(p_0[1]));
   NAND2_X1 i_115 (.A1(n_84), .A2(n_77), .ZN(n_74));
   INV_X1 i_116 (.A(A_in[0]), .ZN(n_77));
   INV_X1 i_119 (.A(A_in[1]), .ZN(n_84));
   NOR3_X1 i_126 (.A1(A_in[9]), .A2(A_in[8]), .A3(A_in[10]), .ZN(n_87));
   INV_X1 i_127 (.A(A_in[8]), .ZN(n_88));
   INV_X1 i_128 (.A(A_in[9]), .ZN(n_90));
   INV_X1 i_129 (.A(A_in[10]), .ZN(n_103));
endmodule

module datapath__0_0(A_imm, A_imm_2s_complement);
   input [31:0]A_imm;
   output [31:0]A_imm_2s_complement;

   AOI21_X1 i_1 (.A(n_19), .B1(A_imm[2]), .B2(n_13), .ZN(A_imm_2s_complement[2]));
   AOI21_X1 i_6 (.A(n_55), .B1(A_imm[7]), .B2(n_0), .ZN(A_imm_2s_complement[7]));
   INV_X1 i_7 (.A(n_1), .ZN(n_0));
   INV_X1 i_3 (.A(n_23), .ZN(n_55));
   INV_X1 i_5 (.A(n_2), .ZN(A_imm_2s_complement[9]));
   XNOR2_X1 i_8 (.A(n_45), .B(A_imm[9]), .ZN(n_2));
   INV_X1 i_9 (.A(n_3), .ZN(A_imm_2s_complement[10]));
   XNOR2_X1 i_10 (.A(n_43), .B(n_34), .ZN(n_3));
   INV_X1 i_11 (.A(n_4), .ZN(A_imm_2s_complement[12]));
   XNOR2_X1 i_12 (.A(n_5), .B(A_imm[12]), .ZN(n_4));
   NAND3_X1 i_13 (.A1(n_43), .A2(n_33), .A3(n_34), .ZN(n_5));
   INV_X1 i_23 (.A(n_12), .ZN(A_imm_2s_complement[4]));
   XNOR2_X1 i_24 (.A(n_7), .B(n_35), .ZN(n_12));
   INV_X1 i_25 (.A(n_14), .ZN(A_imm_2s_complement[5]));
   OR2_X1 i_26 (.A1(n_57), .A2(n_17), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_8), .B1(n_7), .B2(n_35), .ZN(n_17));
   INV_X1 i_28 (.A(n_18), .ZN(A_imm_2s_complement[6]));
   NAND2_X1 i_29 (.A1(n_24), .A2(n_20), .ZN(n_18));
   NAND2_X1 i_30 (.A1(n_47), .A2(A_imm[6]), .ZN(n_20));
   INV_X1 i_31 (.A(n_21), .ZN(A_imm_2s_complement[8]));
   NAND2_X1 i_32 (.A1(n_22), .A2(n_45), .ZN(n_21));
   NAND2_X1 i_33 (.A1(n_23), .A2(A_imm[8]), .ZN(n_22));
   NAND2_X1 i_34 (.A1(n_1), .A2(n_114), .ZN(n_23));
   INV_X1 i_35 (.A(n_24), .ZN(n_1));
   NAND2_X1 i_36 (.A1(n_57), .A2(n_113), .ZN(n_24));
   INV_X1 i_37 (.A(n_25), .ZN(A_imm_2s_complement[11]));
   NAND2_X1 i_38 (.A1(n_26), .A2(n_28), .ZN(n_25));
   NAND2_X1 i_39 (.A1(n_27), .A2(A_imm[11]), .ZN(n_26));
   NAND3_X1 i_40 (.A1(n_34), .A2(n_30), .A3(n_29), .ZN(n_27));
   NAND4_X1 i_41 (.A1(n_34), .A2(n_30), .A3(n_31), .A4(n_29), .ZN(n_28));
   INV_X1 i_42 (.A(n_45), .ZN(n_29));
   INV_X1 i_43 (.A(A_imm[9]), .ZN(n_30));
   INV_X1 i_44 (.A(A_imm[11]), .ZN(n_31));
   AOI21_X1 i_0 (.A(n_77), .B1(n_32), .B2(A_imm[18]), .ZN(
      A_imm_2s_complement[18]));
   OR2_X1 i_2 (.A1(n_50), .A2(A_imm[17]), .ZN(n_32));
   INV_X1 i_47 (.A(A_imm[11]), .ZN(n_33));
   INV_X1 i_48 (.A(A_imm[10]), .ZN(n_34));
   INV_X1 i_61 (.A(n_57), .ZN(n_47));
   INV_X1 i_4 (.A(n_48), .ZN(A_imm_2s_complement[17]));
   NAND2_X1 i_14 (.A1(n_49), .A2(n_51), .ZN(n_48));
   NAND2_X1 i_15 (.A1(n_50), .A2(A_imm[17]), .ZN(n_49));
   NAND3_X1 i_16 (.A1(n_54), .A2(n_53), .A3(n_52), .ZN(n_50));
   NAND4_X1 i_17 (.A1(n_54), .A2(n_52), .A3(n_56), .A4(n_53), .ZN(n_51));
   INV_X1 i_18 (.A(n_40), .ZN(n_52));
   NOR3_X1 i_19 (.A1(A_imm[14]), .A2(A_imm[16]), .A3(A_imm[15]), .ZN(n_53));
   INV_X1 i_20 (.A(A_imm[13]), .ZN(n_54));
   INV_X1 i_21 (.A(A_imm[17]), .ZN(n_56));
   INV_X1 i_71 (.A(n_63), .ZN(n_57));
   NAND2_X1 i_72 (.A1(n_35), .A2(n_11), .ZN(n_63));
   INV_X1 i_76 (.A(n_65), .ZN(A_imm_2s_complement[13]));
   NAND2_X1 i_77 (.A1(n_38), .A2(n_66), .ZN(n_65));
   NAND2_X1 i_78 (.A1(n_40), .A2(A_imm[13]), .ZN(n_66));
   INV_X1 i_79 (.A(n_67), .ZN(A_imm_2s_complement[14]));
   NAND2_X1 i_80 (.A1(n_68), .A2(n_70), .ZN(n_67));
   NAND2_X1 i_81 (.A1(n_38), .A2(A_imm[14]), .ZN(n_68));
   NAND3_X1 i_83 (.A1(n_39), .A2(n_60), .A3(n_59), .ZN(n_70));
   AOI21_X1 i_87 (.A(n_61), .B1(A_imm[15]), .B2(n_37), .ZN(
      A_imm_2s_complement[15]));
   AOI21_X1 i_22 (.A(n_79), .B1(n_76), .B2(A_imm[21]), .ZN(
      A_imm_2s_complement[21]));
   AOI21_X1 i_45 (.A(n_90), .B1(A_imm[22]), .B2(n_80), .ZN(
      A_imm_2s_complement[22]));
   INV_X1 i_46 (.A(n_82), .ZN(n_90));
   AOI21_X1 i_49 (.A(n_85), .B1(n_82), .B2(A_imm[23]), .ZN(
      A_imm_2s_complement[23]));
   AOI22_X1 i_50 (.A1(n_100), .A2(A_imm[26]), .B1(n_85), .B2(n_97), .ZN(
      A_imm_2s_complement[26]));
   NAND2_X1 i_51 (.A1(n_85), .A2(n_91), .ZN(n_100));
   INV_X1 i_174 (.A(A_imm[10]), .ZN(n_9));
   INV_X1 i_175 (.A(A_imm[11]), .ZN(n_10));
   INV_X1 i_186 (.A(n_6), .ZN(n_11));
   NAND2_X1 i_187 (.A1(n_8), .A2(n_7), .ZN(n_6));
   INV_X1 i_188 (.A(A_imm[4]), .ZN(n_7));
   INV_X1 i_189 (.A(A_imm[5]), .ZN(n_8));
   AOI21_X1 i_52 (.A(n_15), .B1(A_imm[1]), .B2(A_imm[0]), .ZN(
      A_imm_2s_complement[1]));
   INV_X1 i_53 (.A(n_15), .ZN(n_13));
   NOR2_X1 i_54 (.A1(A_imm[1]), .A2(A_imm[0]), .ZN(n_15));
   AOI21_X1 i_55 (.A(n_35), .B1(A_imm[3]), .B2(n_16), .ZN(A_imm_2s_complement[3]));
   INV_X1 i_56 (.A(n_19), .ZN(n_16));
   NOR2_X1 i_57 (.A1(A_imm[2]), .A2(n_13), .ZN(n_19));
   AND2_X1 i_58 (.A1(n_15), .A2(n_36), .ZN(n_35));
   NOR2_X1 i_59 (.A1(A_imm[3]), .A2(A_imm[2]), .ZN(n_36));
   NAND3_X1 i_60 (.A1(n_59), .A2(n_39), .A3(n_60), .ZN(n_37));
   NAND2_X1 i_62 (.A1(n_59), .A2(n_39), .ZN(n_38));
   INV_X1 i_63 (.A(n_40), .ZN(n_39));
   NAND2_X1 i_64 (.A1(n_43), .A2(n_41), .ZN(n_40));
   AND2_X1 i_65 (.A1(n_58), .A2(n_42), .ZN(n_41));
   AND2_X1 i_66 (.A1(n_10), .A2(n_9), .ZN(n_42));
   NOR2_X1 i_67 (.A1(A_imm[9]), .A2(n_45), .ZN(n_43));
   INV_X1 i_68 (.A(n_45), .ZN(n_44));
   NAND4_X1 i_69 (.A1(n_112), .A2(n_15), .A3(n_36), .A4(n_11), .ZN(n_45));
   INV_X1 i_70 (.A(A_imm[9]), .ZN(n_46));
   INV_X1 i_73 (.A(A_imm[12]), .ZN(n_58));
   INV_X1 i_74 (.A(A_imm[13]), .ZN(n_59));
   INV_X1 i_75 (.A(A_imm[14]), .ZN(n_60));
   XNOR2_X1 i_82 (.A(A_imm[16]), .B(n_61), .ZN(A_imm_2s_complement[16]));
   NOR3_X1 i_84 (.A1(A_imm[15]), .A2(A_imm[14]), .A3(n_62), .ZN(n_61));
   NAND3_X1 i_85 (.A1(n_43), .A2(n_59), .A3(n_41), .ZN(n_62));
   INV_X1 i_86 (.A(A_imm[16]), .ZN(n_64));
   XNOR2_X1 i_88 (.A(n_74), .B(n_69), .ZN(A_imm_2s_complement[19]));
   NAND3_X1 i_89 (.A1(n_44), .A2(n_46), .A3(n_71), .ZN(n_69));
   NOR2_X1 i_90 (.A1(n_73), .A2(n_72), .ZN(n_71));
   OR4_X1 i_91 (.A1(A_imm[18]), .A2(A_imm[17]), .A3(A_imm[15]), .A4(A_imm[14]), 
      .ZN(n_72));
   NAND4_X1 i_92 (.A1(n_58), .A2(n_64), .A3(n_59), .A4(n_42), .ZN(n_73));
   INV_X1 i_93 (.A(A_imm[19]), .ZN(n_74));
   AND2_X1 i_94 (.A1(n_76), .A2(n_75), .ZN(A_imm_2s_complement[20]));
   OAI21_X1 i_95 (.A(A_imm[20]), .B1(A_imm[19]), .B2(n_69), .ZN(n_75));
   NAND3_X1 i_96 (.A1(n_77), .A2(n_74), .A3(n_78), .ZN(n_76));
   INV_X1 i_97 (.A(n_69), .ZN(n_77));
   INV_X1 i_98 (.A(A_imm[20]), .ZN(n_78));
   INV_X1 i_99 (.A(n_80), .ZN(n_79));
   NAND3_X1 i_100 (.A1(n_77), .A2(n_74), .A3(n_81), .ZN(n_80));
   NOR2_X1 i_101 (.A1(A_imm[21]), .A2(A_imm[20]), .ZN(n_81));
   NAND4_X1 i_102 (.A1(n_77), .A2(n_78), .A3(n_74), .A4(n_83), .ZN(n_82));
   NOR2_X1 i_103 (.A1(A_imm[22]), .A2(A_imm[21]), .ZN(n_83));
   AOI22_X1 i_104 (.A1(n_89), .A2(n_85), .B1(A_imm[24]), .B2(n_86), .ZN(
      A_imm_2s_complement[24]));
   NAND2_X1 i_105 (.A1(n_89), .A2(n_85), .ZN(n_84));
   INV_X1 i_106 (.A(n_86), .ZN(n_85));
   NAND4_X1 i_107 (.A1(n_44), .A2(n_71), .A3(n_46), .A4(n_87), .ZN(n_86));
   NOR4_X1 i_108 (.A1(A_imm[23]), .A2(A_imm[22]), .A3(n_88), .A4(A_imm[21]), 
      .ZN(n_87));
   NAND2_X1 i_109 (.A1(n_78), .A2(n_74), .ZN(n_88));
   INV_X1 i_110 (.A(A_imm[24]), .ZN(n_89));
   AOI22_X1 i_111 (.A1(A_imm[25]), .A2(n_84), .B1(n_85), .B2(n_91), .ZN(
      A_imm_2s_complement[25]));
   AND2_X1 i_112 (.A1(n_92), .A2(n_89), .ZN(n_91));
   INV_X1 i_113 (.A(A_imm[25]), .ZN(n_92));
   AOI21_X1 i_114 (.A(n_94), .B1(A_imm[27]), .B2(n_93), .ZN(
      A_imm_2s_complement[27]));
   NAND2_X1 i_115 (.A1(n_85), .A2(n_97), .ZN(n_93));
   INV_X1 i_116 (.A(n_95), .ZN(n_94));
   NAND4_X1 i_117 (.A1(n_43), .A2(n_71), .A3(n_87), .A4(n_96), .ZN(n_95));
   NOR2_X1 i_118 (.A1(A_imm[27]), .A2(n_98), .ZN(n_96));
   INV_X1 i_119 (.A(n_98), .ZN(n_97));
   NAND3_X1 i_120 (.A1(n_92), .A2(n_89), .A3(n_99), .ZN(n_98));
   INV_X1 i_121 (.A(A_imm[26]), .ZN(n_99));
   OAI22_X1 i_122 (.A1(A_imm[28]), .A2(n_94), .B1(n_101), .B2(n_95), .ZN(
      A_imm_2s_complement[28]));
   INV_X1 i_123 (.A(A_imm[28]), .ZN(n_101));
   XNOR2_X1 i_124 (.A(A_imm[29]), .B(n_102), .ZN(A_imm_2s_complement[29]));
   NOR2_X1 i_125 (.A1(A_imm[28]), .A2(n_95), .ZN(n_102));
   NOR2_X1 i_126 (.A1(A_imm[30]), .A2(A_imm[29]), .ZN(n_103));
   NAND4_X1 i_127 (.A1(n_103), .A2(n_85), .A3(n_96), .A4(n_101), .ZN(n_104));
   INV_X1 i_128 (.A(A_imm[30]), .ZN(n_105));
   INV_X1 i_129 (.A(A_imm[29]), .ZN(n_106));
   INV_X1 i_130 (.A(n_104), .ZN(n_107));
   NAND3_X1 i_131 (.A1(n_106), .A2(n_101), .A3(n_94), .ZN(n_108));
   AOI21_X1 i_132 (.A(n_107), .B1(A_imm[30]), .B2(n_108), .ZN(
      A_imm_2s_complement[30]));
   AOI21_X1 i_133 (.A(n_109), .B1(A_imm[31]), .B2(n_104), .ZN(
      A_imm_2s_complement[31]));
   NOR3_X1 i_134 (.A1(A_imm[31]), .A2(n_111), .A3(n_110), .ZN(n_109));
   NAND3_X1 i_135 (.A1(n_85), .A2(n_101), .A3(n_96), .ZN(n_110));
   NAND2_X1 i_136 (.A1(n_105), .A2(n_106), .ZN(n_111));
   NOR3_X1 i_137 (.A1(A_imm[8]), .A2(A_imm[6]), .A3(A_imm[7]), .ZN(n_112));
   INV_X1 i_138 (.A(A_imm[6]), .ZN(n_113));
   INV_X1 i_139 (.A(A_imm[7]), .ZN(n_114));
endmodule

module datapath__0_1(B_in, p_0);
   input [31:0]B_in;
   output [31:0]p_0;

   AOI21_X1 i_0 (.A(n_3), .B1(B_in[1]), .B2(B_in[0]), .ZN(p_0[1]));
   AOI21_X1 i_1 (.A(n_37), .B1(B_in[3]), .B2(n_2), .ZN(p_0[3]));
   AOI21_X1 i_2 (.A(n_13), .B1(B_in[5]), .B2(n_15), .ZN(p_0[5]));
   AOI21_X1 i_3 (.A(n_26), .B1(B_in[7]), .B2(n_0), .ZN(p_0[7]));
   INV_X1 i_4 (.A(n_14), .ZN(n_0));
   AOI21_X1 i_5 (.A(n_11), .B1(B_in[8]), .B2(n_25), .ZN(p_0[8]));
   AOI21_X1 i_6 (.A(n_9), .B1(B_in[9]), .B2(n_10), .ZN(p_0[9]));
   AOI21_X1 i_7 (.A(n_24), .B1(B_in[10]), .B2(n_8), .ZN(p_0[10]));
   AOI21_X1 i_8 (.A(n_66), .B1(B_in[11]), .B2(n_19), .ZN(p_0[11]));
   INV_X1 i_9 (.A(n_9), .ZN(n_8));
   NOR2_X1 i_10 (.A1(B_in[9]), .A2(n_10), .ZN(n_9));
   INV_X1 i_11 (.A(n_11), .ZN(n_10));
   NOR2_X1 i_12 (.A1(B_in[8]), .A2(n_25), .ZN(n_11));
   AOI21_X1 i_24 (.A(n_39), .B1(B_in[13]), .B2(n_41), .ZN(p_0[13]));
   AOI21_X1 i_33 (.A(n_23), .B1(B_in[16]), .B2(n_51), .ZN(p_0[16]));
   AOI21_X1 i_34 (.A(n_21), .B1(B_in[17]), .B2(n_22), .ZN(p_0[17]));
   AOI21_X1 i_13 (.A(n_55), .B1(B_in[18]), .B2(n_20), .ZN(p_0[18]));
   INV_X1 i_14 (.A(n_21), .ZN(n_20));
   NOR2_X1 i_15 (.A1(B_in[17]), .A2(n_22), .ZN(n_21));
   INV_X1 i_16 (.A(n_23), .ZN(n_22));
   NOR2_X1 i_17 (.A1(B_in[16]), .A2(n_51), .ZN(n_23));
   AOI21_X1 i_43 (.A(n_61), .B1(B_in[20]), .B2(n_56), .ZN(p_0[20]));
   AOI21_X1 i_18 (.A(n_78), .B1(B_in[23]), .B2(n_63), .ZN(p_0[23]));
   AOI21_X1 i_19 (.A(n_69), .B1(B_in[24]), .B2(n_70), .ZN(p_0[24]));
   NOR2_X1 i_20 (.A1(n_47), .A2(n_48), .ZN(p_0[28]));
   AOI21_X1 i_21 (.A(n_50), .B1(n_78), .B2(n_76), .ZN(n_47));
   INV_X1 i_22 (.A(n_49), .ZN(n_48));
   AOI22_X1 i_23 (.A1(n_49), .A2(B_in[29]), .B1(n_75), .B2(n_79), .ZN(p_0[29]));
   NAND4_X1 i_25 (.A1(n_62), .A2(n_50), .A3(n_71), .A4(n_76), .ZN(n_49));
   INV_X1 i_26 (.A(B_in[28]), .ZN(n_50));
   INV_X1 i_27 (.A(n_1), .ZN(p_0[2]));
   OAI21_X1 i_28 (.A(n_2), .B1(n_4), .B2(n_3), .ZN(n_1));
   NAND2_X1 i_29 (.A1(n_4), .A2(n_3), .ZN(n_2));
   NOR2_X1 i_30 (.A1(B_in[1]), .A2(B_in[0]), .ZN(n_3));
   INV_X1 i_31 (.A(B_in[2]), .ZN(n_4));
   AOI21_X1 i_32 (.A(n_5), .B1(B_in[4]), .B2(n_6), .ZN(p_0[4]));
   NOR2_X1 i_35 (.A1(B_in[4]), .A2(n_6), .ZN(n_5));
   OR4_X1 i_36 (.A1(B_in[3]), .A2(B_in[0]), .A3(n_7), .A4(B_in[1]), .ZN(n_6));
   INV_X1 i_37 (.A(n_4), .ZN(n_7));
   AOI21_X1 i_38 (.A(n_14), .B1(B_in[6]), .B2(n_12), .ZN(p_0[6]));
   INV_X1 i_39 (.A(n_13), .ZN(n_12));
   NOR2_X1 i_40 (.A1(B_in[5]), .A2(n_15), .ZN(n_13));
   NOR4_X1 i_41 (.A1(B_in[5]), .A2(B_in[4]), .A3(B_in[6]), .A4(n_6), .ZN(n_14));
   INV_X1 i_42 (.A(n_5), .ZN(n_15));
   INV_X1 i_44 (.A(B_in[4]), .ZN(n_16));
   INV_X1 i_45 (.A(B_in[5]), .ZN(n_17));
   INV_X1 i_46 (.A(B_in[6]), .ZN(n_18));
   INV_X1 i_47 (.A(n_24), .ZN(n_19));
   NOR4_X1 i_48 (.A1(B_in[10]), .A2(B_in[9]), .A3(B_in[8]), .A4(n_25), .ZN(n_24));
   INV_X1 i_49 (.A(n_26), .ZN(n_25));
   NOR2_X1 i_50 (.A1(n_6), .A2(n_27), .ZN(n_26));
   NAND4_X1 i_51 (.A1(n_17), .A2(n_16), .A3(n_28), .A4(n_18), .ZN(n_27));
   INV_X1 i_52 (.A(B_in[7]), .ZN(n_28));
   INV_X1 i_53 (.A(B_in[8]), .ZN(n_29));
   INV_X1 i_54 (.A(B_in[9]), .ZN(n_30));
   INV_X1 i_55 (.A(B_in[10]), .ZN(n_31));
   AOI21_X1 i_56 (.A(n_32), .B1(B_in[12]), .B2(n_33), .ZN(p_0[12]));
   NOR2_X1 i_57 (.A1(B_in[12]), .A2(n_33), .ZN(n_32));
   NAND3_X1 i_58 (.A1(n_37), .A2(n_36), .A3(n_34), .ZN(n_33));
   AND4_X1 i_59 (.A1(n_30), .A2(n_29), .A3(n_35), .A4(n_31), .ZN(n_34));
   INV_X1 i_60 (.A(B_in[11]), .ZN(n_35));
   INV_X1 i_61 (.A(n_27), .ZN(n_36));
   INV_X1 i_62 (.A(n_6), .ZN(n_37));
   AOI21_X1 i_63 (.A(n_40), .B1(B_in[14]), .B2(n_38), .ZN(p_0[14]));
   INV_X1 i_64 (.A(n_39), .ZN(n_38));
   NOR2_X1 i_65 (.A1(B_in[13]), .A2(n_41), .ZN(n_39));
   NOR4_X1 i_66 (.A1(B_in[13]), .A2(B_in[12]), .A3(B_in[14]), .A4(n_33), 
      .ZN(n_40));
   INV_X1 i_67 (.A(n_32), .ZN(n_41));
   INV_X1 i_68 (.A(B_in[12]), .ZN(n_42));
   INV_X1 i_69 (.A(B_in[13]), .ZN(n_43));
   INV_X1 i_70 (.A(B_in[14]), .ZN(n_44));
   INV_X1 i_71 (.A(n_45), .ZN(p_0[15]));
   OAI21_X1 i_72 (.A(n_51), .B1(n_53), .B2(n_40), .ZN(n_45));
   INV_X1 i_73 (.A(n_51), .ZN(n_46));
   NAND4_X1 i_74 (.A1(n_37), .A2(n_36), .A3(n_34), .A4(n_52), .ZN(n_51));
   AND4_X1 i_75 (.A1(n_43), .A2(n_42), .A3(n_53), .A4(n_44), .ZN(n_52));
   INV_X1 i_76 (.A(B_in[15]), .ZN(n_53));
   AOI22_X1 i_77 (.A1(n_46), .A2(n_57), .B1(B_in[19]), .B2(n_54), .ZN(p_0[19]));
   INV_X1 i_78 (.A(n_55), .ZN(n_54));
   NOR2_X1 i_79 (.A1(n_51), .A2(n_58), .ZN(n_55));
   NAND2_X1 i_80 (.A1(n_46), .A2(n_57), .ZN(n_56));
   NOR2_X1 i_81 (.A1(B_in[19]), .A2(n_58), .ZN(n_57));
   OR3_X1 i_82 (.A1(B_in[17]), .A2(B_in[16]), .A3(B_in[18]), .ZN(n_58));
   AOI21_X1 i_83 (.A(n_59), .B1(B_in[21]), .B2(n_60), .ZN(p_0[21]));
   NOR2_X1 i_84 (.A1(B_in[21]), .A2(n_60), .ZN(n_59));
   INV_X1 i_85 (.A(n_61), .ZN(n_60));
   NOR2_X1 i_86 (.A1(B_in[20]), .A2(n_56), .ZN(n_61));
   AOI21_X1 i_87 (.A(n_62), .B1(B_in[22]), .B2(n_65), .ZN(p_0[22]));
   INV_X1 i_88 (.A(n_63), .ZN(n_62));
   NAND4_X1 i_89 (.A1(n_66), .A2(n_52), .A3(n_57), .A4(n_64), .ZN(n_63));
   NOR3_X1 i_90 (.A1(B_in[22]), .A2(B_in[20]), .A3(B_in[21]), .ZN(n_64));
   INV_X1 i_91 (.A(n_59), .ZN(n_65));
   INV_X1 i_92 (.A(n_33), .ZN(n_66));
   INV_X1 i_93 (.A(n_67), .ZN(p_0[25]));
   OAI21_X1 i_94 (.A(n_68), .B1(n_72), .B2(n_69), .ZN(n_67));
   NAND2_X1 i_95 (.A1(n_72), .A2(n_69), .ZN(n_68));
   NOR2_X1 i_96 (.A1(B_in[24]), .A2(n_70), .ZN(n_69));
   NAND4_X1 i_97 (.A1(n_71), .A2(n_46), .A3(n_57), .A4(n_64), .ZN(n_70));
   INV_X1 i_98 (.A(B_in[23]), .ZN(n_71));
   INV_X1 i_99 (.A(B_in[25]), .ZN(n_72));
   AOI21_X1 i_100 (.A(n_73), .B1(B_in[26]), .B2(n_68), .ZN(p_0[26]));
   NOR2_X1 i_101 (.A1(n_70), .A2(n_74), .ZN(n_73));
   OR3_X1 i_102 (.A1(B_in[26]), .A2(B_in[24]), .A3(B_in[25]), .ZN(n_74));
   AOI21_X1 i_103 (.A(n_75), .B1(B_in[27]), .B2(n_77), .ZN(p_0[27]));
   NOR3_X1 i_104 (.A1(n_74), .A2(B_in[27]), .A3(n_70), .ZN(n_75));
   NOR2_X1 i_105 (.A1(n_74), .A2(B_in[27]), .ZN(n_76));
   INV_X1 i_106 (.A(n_73), .ZN(n_77));
   INV_X1 i_107 (.A(n_70), .ZN(n_78));
   NOR2_X1 i_108 (.A1(B_in[29]), .A2(B_in[28]), .ZN(n_79));
   INV_X1 i_109 (.A(B_in[30]), .ZN(n_80));
   NAND4_X1 i_110 (.A1(n_79), .A2(n_80), .A3(n_78), .A4(n_76), .ZN(n_81));
   INV_X1 i_111 (.A(n_81), .ZN(n_82));
   NAND4_X1 i_112 (.A1(n_79), .A2(n_62), .A3(n_76), .A4(n_71), .ZN(n_83));
   AOI21_X1 i_113 (.A(n_82), .B1(n_83), .B2(B_in[30]), .ZN(p_0[30]));
   XOR2_X1 i_114 (.A(n_81), .B(B_in[31]), .Z(p_0[31]));
endmodule

module datapath__0_67(p_0, p_1, p_2, p_3, p_4, p_5, p_6, p_7, p_8, p_9, p_10, 
      p_11, p_12, p_13, p_14, p_15, \aggregated_res[14] );
   input [63:0]p_0;
   input [63:0]p_1;
   input [63:0]p_2;
   input [63:0]p_3;
   input [63:0]p_4;
   input [63:0]p_5;
   input [63:0]p_6;
   input [63:0]p_7;
   input [63:0]p_8;
   input [63:0]p_9;
   input [63:0]p_10;
   input [63:0]p_11;
   input [63:0]p_12;
   input [63:0]p_13;
   input [63:0]p_14;
   input [63:0]p_15;
   output [63:0]\aggregated_res[14] ;

   OAI222_X1 i_0 (.A1(p_5[44]), .A2(n_1175), .B1(p_5[44]), .B2(n_1315), .C1(
      n_1315), .C2(n_1175), .ZN(n_16));
   INV_X1 i_1 (.A(n_912), .ZN(\aggregated_res[14] [2]));
   OAI21_X1 i_2 (.A(n_97), .B1(p_0[2]), .B2(p_15[2]), .ZN(n_912));
   XOR2_X1 i_3 (.A(n_97), .B(n_913), .Z(\aggregated_res[14] [3]));
   OAI21_X1 i_4 (.A(n_96), .B1(p_0[3]), .B2(p_15[3]), .ZN(n_913));
   XNOR2_X1 i_5 (.A(n_81), .B(n_914), .ZN(\aggregated_res[14] [4]));
   OAI21_X1 i_6 (.A(n_99), .B1(p_15[4]), .B2(n_38), .ZN(n_914));
   XOR2_X1 i_7 (.A(n_77), .B(n_915), .Z(\aggregated_res[14] [5]));
   XOR2_X1 i_8 (.A(n_49), .B(n_25), .Z(n_915));
   XOR2_X1 i_9 (.A(n_73), .B(n_922), .Z(\aggregated_res[14] [6]));
   XOR2_X1 i_10 (.A(n_69), .B(n_918), .Z(\aggregated_res[14] [7]));
   AOI21_X1 i_11 (.A(n_105), .B1(n_31), .B2(n_29), .ZN(n_918));
   OAI21_X1 i_12 (.A(n_71), .B1(n_23), .B2(n_27), .ZN(n_922));
   XOR2_X1 i_13 (.A(n_273), .B(n_926), .Z(\aggregated_res[14] [11]));
   AOI21_X1 i_14 (.A(n_271), .B1(n_145), .B2(n_185), .ZN(n_926));
   XOR2_X1 i_15 (.A(n_417), .B(n_932), .Z(\aggregated_res[14] [16]));
   NOR2_X1 i_16 (.A1(n_525), .A2(n_418), .ZN(n_932));
   XNOR2_X1 i_17 (.A(n_947), .B(n_941), .ZN(\aggregated_res[14] [21]));
   OAI21_X1 i_18 (.A(n_453), .B1(n_1137), .B2(n_943), .ZN(n_941));
   AOI21_X1 i_19 (.A(n_543), .B1(n_447), .B2(n_455), .ZN(n_947));
   XOR2_X1 i_20 (.A(n_953), .B(n_950), .Z(\aggregated_res[14] [23]));
   XOR2_X1 i_21 (.A(n_951), .B(n_948), .Z(\aggregated_res[14] [24]));
   NOR2_X1 i_22 (.A1(n_659), .A2(n_649), .ZN(n_948));
   XNOR2_X1 i_23 (.A(n_955), .B(n_949), .ZN(\aggregated_res[14] [25]));
   OAI21_X1 i_24 (.A(n_657), .B1(n_649), .B2(n_951), .ZN(n_949));
   NOR2_X1 i_25 (.A1(n_655), .A2(n_1121), .ZN(n_950));
   INV_X1 i_26 (.A(n_952), .ZN(n_951));
   OAI21_X1 i_27 (.A(n_653), .B1(n_1121), .B2(n_953), .ZN(n_952));
   AOI21_X1 i_28 (.A(n_636), .B1(n_511), .B2(n_507), .ZN(n_953));
   AOI21_X1 i_29 (.A(n_661), .B1(n_555), .B2(n_551), .ZN(n_955));
   XOR2_X1 i_30 (.A(n_961), .B(n_958), .Z(\aggregated_res[14] [27]));
   XOR2_X1 i_31 (.A(n_959), .B(n_956), .Z(\aggregated_res[14] [28]));
   NOR2_X1 i_32 (.A1(n_752), .A2(n_1131), .ZN(n_956));
   NOR2_X1 i_33 (.A1(n_1160), .A2(n_731), .ZN(n_958));
   XOR2_X1 i_34 (.A(n_983), .B(n_984), .Z(\aggregated_res[14] [34]));
   XOR2_X1 i_35 (.A(n_981), .B(n_944), .Z(\aggregated_res[14] [35]));
   OAI21_X1 i_36 (.A(n_1000), .B1(n_896), .B2(n_938), .ZN(n_984));
   XOR2_X1 i_37 (.A(n_1013), .B(n_992), .Z(\aggregated_res[14] [38]));
   XOR2_X1 i_38 (.A(n_991), .B(n_988), .Z(\aggregated_res[14] [39]));
   NOR2_X1 i_39 (.A1(n_1094), .A2(n_1097), .ZN(n_988));
   OAI21_X1 i_40 (.A(n_1072), .B1(n_1018), .B2(n_1078), .ZN(n_992));
   XOR2_X1 i_41 (.A(n_1007), .B(n_1218), .Z(\aggregated_res[14] [47]));
   XNOR2_X1 i_42 (.A(n_1003), .B(n_1002), .ZN(\aggregated_res[14] [48]));
   OAI22_X1 i_43 (.A1(n_1184), .A2(n_1208), .B1(n_1219), .B2(n_1007), .ZN(n_1002));
   NOR2_X1 i_44 (.A1(n_1216), .A2(n_1221), .ZN(n_1003));
   INV_X1 i_45 (.A(n_1217), .ZN(n_1007));
   XOR2_X1 i_46 (.A(n_1047), .B(n_1030), .Z(\aggregated_res[14] [54]));
   XOR2_X1 i_47 (.A(n_1029), .B(n_1026), .Z(\aggregated_res[14] [55]));
   NOR2_X1 i_48 (.A1(n_1393), .A2(n_1394), .ZN(n_1026));
   OAI21_X1 i_49 (.A(n_1250), .B1(n_1293), .B2(n_1384), .ZN(n_1030));
   AOI22_X1 i_50 (.A1(n_1039), .A2(n_1369), .B1(n_1040), .B2(n_1370), .ZN(
      \aggregated_res[14] [59]));
   INV_X1 i_51 (.A(n_651), .ZN(n_1121));
   AOI21_X1 i_52 (.A(n_1267), .B1(n_1207), .B2(n_1237), .ZN(n_1235));
   OAI211_X1 i_53 (.A(n_1309), .B(n_1241), .C1(n_1281), .C2(n_1292), .ZN(n_1238));
   INV_X1 i_54 (.A(p_14[61]), .ZN(n_1283));
   INV_X1 i_55 (.A(p_6[44]), .ZN(n_1315));
   INV_X1 i_56 (.A(n_451), .ZN(n_1137));
   XOR2_X1 i_57 (.A(n_519), .B(n_927), .Z(\aggregated_res[14] [18]));
   NAND2_X1 i_58 (.A1(n_1400), .A2(n_537), .ZN(n_927));
   XOR2_X1 i_59 (.A(n_931), .B(n_930), .Z(\aggregated_res[14] [19]));
   NAND2_X1 i_60 (.A1(n_533), .A2(n_539), .ZN(n_930));
   XNOR2_X1 i_61 (.A(n_449), .B(n_943), .ZN(\aggregated_res[14] [20]));
   AOI21_X1 i_62 (.A(n_535), .B1(n_539), .B2(n_931), .ZN(n_943));
   AOI21_X1 i_63 (.A(n_517), .B1(n_407), .B2(n_459), .ZN(n_931));
   XNOR2_X1 i_64 (.A(n_267), .B(n_994), .ZN(\aggregated_res[14] [12]));
   NAND2_X1 i_65 (.A1(n_275), .A2(n_263), .ZN(n_994));
   XOR2_X1 i_66 (.A(n_387), .B(n_363), .Z(\aggregated_res[14] [14]));
   INV_X1 i_67 (.A(n_1040), .ZN(n_1039));
   NAND2_X1 i_68 (.A1(n_1117), .A2(n_1347), .ZN(n_1040));
   OAI21_X1 i_69 (.A(n_1250), .B1(n_1047), .B2(n_1090), .ZN(n_1029));
   OAI21_X1 i_70 (.A(n_1072), .B1(n_1013), .B2(n_1365), .ZN(n_991));
   AOI21_X1 i_71 (.A(p_6[42]), .B1(p_5[42]), .B2(n_1044), .ZN(n_17));
   INV_X1 i_72 (.A(p_4[42]), .ZN(n_1044));
   INV_X1 i_674 (.A(p_5[42]), .ZN(n_19));
   INV_X1 i_685 (.A(p_1[36]), .ZN(n_21));
   XOR2_X1 i_73 (.A(n_1059), .B(n_1362), .Z(\aggregated_res[14] [40]));
   NAND2_X1 i_74 (.A1(n_1075), .A2(n_1367), .ZN(n_1059));
   NAND2_X1 i_75 (.A1(n_1169), .A2(n_1173), .ZN(n_1067));
   XNOR2_X1 i_76 (.A(n_1073), .B(n_1071), .ZN(\aggregated_res[14] [56]));
   NOR2_X1 i_77 (.A1(n_1391), .A2(n_1091), .ZN(n_1071));
   NAND2_X1 i_78 (.A1(n_1083), .A2(n_1392), .ZN(n_1073));
   NAND2_X1 i_79 (.A1(n_1076), .A2(n_1074), .ZN(\aggregated_res[14] [57]));
   OAI21_X1 i_80 (.A(n_1328), .B1(n_1081), .B2(n_1391), .ZN(n_1074));
   NAND2_X1 i_81 (.A1(n_1080), .A2(n_1327), .ZN(n_1076));
   NOR2_X1 i_82 (.A1(n_1081), .A2(n_1391), .ZN(n_1080));
   AOI21_X1 i_83 (.A(n_1091), .B1(n_1083), .B2(n_1392), .ZN(n_1081));
   OAI211_X1 i_84 (.A(n_1395), .B(n_1250), .C1(n_1047), .C2(n_1090), .ZN(n_1083));
   NAND2_X1 i_85 (.A1(n_1384), .A2(n_1293), .ZN(n_1250));
   NOR2_X1 i_86 (.A1(n_1384), .A2(n_1293), .ZN(n_1090));
   INV_X1 i_87 (.A(n_1396), .ZN(n_1091));
   NAND2_X1 i_88 (.A1(n_1098), .A2(n_1100), .ZN(\aggregated_res[14] [60]));
   NAND2_X1 i_89 (.A1(n_1099), .A2(n_1353), .ZN(n_1098));
   NAND2_X1 i_90 (.A1(n_1107), .A2(n_1101), .ZN(n_1099));
   NAND3_X1 i_91 (.A1(n_1107), .A2(n_1352), .A3(n_1101), .ZN(n_1100));
   OR2_X1 i_92 (.A1(n_1344), .A2(n_1350), .ZN(n_1101));
   NAND3_X1 i_93 (.A1(n_1117), .A2(n_1371), .A3(n_1347), .ZN(n_1107));
   NAND2_X1 i_94 (.A1(n_1111), .A2(n_1110), .ZN(\aggregated_res[14] [61]));
   NAND3_X1 i_95 (.A1(n_1114), .A2(n_1124), .A3(n_1118), .ZN(n_1110));
   NAND2_X1 i_96 (.A1(n_1113), .A2(n_1120), .ZN(n_1111));
   NAND2_X1 i_97 (.A1(n_1114), .A2(n_1118), .ZN(n_1113));
   NAND3_X1 i_98 (.A1(n_1117), .A2(n_1347), .A3(n_1368), .ZN(n_1114));
   NAND2_X1 i_99 (.A1(n_0), .A2(n_1348), .ZN(n_1117));
   OR2_X1 i_100 (.A1(n_1377), .A2(n_1355), .ZN(n_1118));
   INV_X1 i_101 (.A(n_1124), .ZN(n_1120));
   NAND2_X1 i_102 (.A1(n_1378), .A2(n_1379), .ZN(n_1124));
   NOR2_X1 i_103 (.A1(n_1125), .A2(n_1127), .ZN(\aggregated_res[14] [62]));
   INV_X1 i_104 (.A(n_1126), .ZN(n_1125));
   NAND3_X1 i_105 (.A1(n_1331), .A2(n_1374), .A3(n_1130), .ZN(n_1126));
   AOI21_X1 i_106 (.A(n_1130), .B1(n_1331), .B2(n_1374), .ZN(n_1127));
   XNOR2_X1 i_107 (.A(n_1283), .B(p_14[62]), .ZN(n_1130));
   NAND2_X1 i_108 (.A1(n_1281), .A2(n_1292), .ZN(n_1145));
   INV_X1 i_109 (.A(n_1269), .ZN(n_1241));
   INV_X1 i_110 (.A(n_1), .ZN(n_1331));
   NOR2_X1 i_111 (.A1(n_7), .A2(n_6), .ZN(n_1047));
   XOR2_X1 i_112 (.A(n_1342), .B(n_1339), .Z(\aggregated_res[14] [29]));
   OAI21_X1 i_113 (.A(n_739), .B1(n_959), .B2(n_1131), .ZN(n_1339));
   AOI21_X1 i_114 (.A(n_1160), .B1(n_1340), .B2(n_733), .ZN(n_959));
   INV_X1 i_115 (.A(n_961), .ZN(n_1340));
   NAND2_X1 i_116 (.A1(n_1341), .A2(n_614), .ZN(n_961));
   OAI21_X1 i_117 (.A(n_616), .B1(n_553), .B2(n_590), .ZN(n_1341));
   NOR2_X1 i_118 (.A1(n_665), .A2(n_592), .ZN(n_1160));
   INV_X1 i_119 (.A(n_727), .ZN(n_1131));
   NAND2_X1 i_120 (.A1(n_765), .A2(n_729), .ZN(n_1342));
   XNOR2_X1 i_121 (.A(n_1361), .B(n_1056), .ZN(\aggregated_res[14] [41]));
   AOI21_X1 i_122 (.A(n_1077), .B1(n_1362), .B2(n_1367), .ZN(n_1361));
   NAND2_X1 i_123 (.A1(n_1363), .A2(n_1095), .ZN(n_1362));
   OAI211_X1 i_124 (.A(n_1072), .B(n_1096), .C1(n_1013), .C2(n_1365), .ZN(n_1363));
   NAND2_X1 i_125 (.A1(n_1078), .A2(n_1018), .ZN(n_1072));
   NOR2_X1 i_126 (.A1(n_1078), .A2(n_1018), .ZN(n_1365));
   INV_X1 i_127 (.A(n_1136), .ZN(n_1013));
   NAND2_X1 i_128 (.A1(n_1033), .A2(n_1070), .ZN(n_1367));
   XNOR2_X1 i_129 (.A(n_1174), .B(n_1067), .ZN(\aggregated_res[14] [44]));
   INV_X1 i_130 (.A(n_1398), .ZN(\aggregated_res[14] [58]));
   XNOR2_X1 i_131 (.A(n_0), .B(n_1346), .ZN(n_1398));
   NAND2_X1 i_132 (.A1(n_4), .A2(n_1386), .ZN(n_0));
   OAI21_X1 i_133 (.A(n_9), .B1(n_1), .B2(n_1373), .ZN(\aggregated_res[14] [63]));
   AOI21_X1 i_134 (.A(n_2), .B1(n_4), .B2(n_1386), .ZN(n_1));
   NAND2_X1 i_135 (.A1(n_1348), .A2(n_3), .ZN(n_2));
   INV_X1 i_136 (.A(n_1376), .ZN(n_3));
   OAI211_X1 i_137 (.A(n_1389), .B(n_5), .C1(n_7), .C2(n_6), .ZN(n_4));
   OR2_X1 i_138 (.A1(n_1384), .A2(n_1293), .ZN(n_5));
   OAI221_X1 i_139 (.A(n_1145), .B1(n_1287), .B2(n_1306), .C1(n_1238), .C2(
      n_1235), .ZN(n_6));
   AND2_X1 i_140 (.A1(n_1245), .A2(n_8), .ZN(n_7));
   NOR2_X1 i_141 (.A1(n_1238), .A2(n_1274), .ZN(n_8));
   NAND2_X1 i_142 (.A1(n_1283), .A2(p_14[62]), .ZN(n_9));
   FA_X1 i_143 (.A(p_0[6]), .B(p_1[6]), .CI(p_2[6]), .CO(n_10), .S(n_23));
   FA_X1 i_144 (.A(p_0[5]), .B(p_1[5]), .CI(p_15[5]), .CO(n_11), .S(n_25));
   HA_X1 i_145 (.A(p_15[6]), .B(n_11), .CO(n_12), .S(n_27));
   FA_X1 i_146 (.A(p_15[7]), .B(n_10), .CI(n_12), .CO(n_13), .S(n_29));
   FA_X1 i_147 (.A(p_0[7]), .B(p_1[7]), .CI(p_2[7]), .CO(n_14), .S(n_31));
   HA_X1 i_148 (.A(p_0[4]), .B(p_1[4]), .CO(n_49), .S(n_38));
   FA_X1 i_149 (.A(p_3[8]), .B(p_15[8]), .CI(n_14), .CO(n_51), .S(n_15));
   HA_X1 i_150 (.A(n_13), .B(n_15), .CO(n_55), .S(n_53));
   FA_X1 i_151 (.A(p_0[8]), .B(p_1[8]), .CI(p_2[8]), .CO(n_58), .S(n_57));
   XNOR2_X1 i_152 (.A(n_65), .B(n_59), .ZN(\aggregated_res[14] [8]));
   OAI21_X1 i_153 (.A(n_63), .B1(n_53), .B2(n_57), .ZN(n_59));
   INV_X1 i_154 (.A(n_63), .ZN(n_61));
   NAND2_X1 i_155 (.A1(n_53), .A2(n_57), .ZN(n_63));
   AOI21_X1 i_156 (.A(n_105), .B1(n_103), .B2(n_67), .ZN(n_65));
   INV_X1 i_157 (.A(n_69), .ZN(n_67));
   AOI21_X1 i_158 (.A(n_101), .B1(n_73), .B2(n_71), .ZN(n_69));
   NAND2_X1 i_159 (.A1(n_23), .A2(n_27), .ZN(n_71));
   OAI22_X1 i_160 (.A1(n_25), .A2(n_49), .B1(n_77), .B2(n_75), .ZN(n_73));
   AND2_X1 i_161 (.A1(n_25), .A2(n_49), .ZN(n_75));
   NAND2_X1 i_162 (.A1(n_99), .A2(n_79), .ZN(n_77));
   OAI21_X1 i_163 (.A(n_81), .B1(n_38), .B2(p_15[4]), .ZN(n_79));
   AOI21_X1 i_164 (.A(n_83), .B1(n_97), .B2(n_96), .ZN(n_81));
   NOR2_X1 i_165 (.A1(p_0[3]), .A2(p_15[3]), .ZN(n_83));
   NAND2_X1 i_166 (.A1(p_0[3]), .A2(p_15[3]), .ZN(n_96));
   NAND2_X1 i_167 (.A1(p_0[2]), .A2(p_15[2]), .ZN(n_97));
   NAND2_X1 i_168 (.A1(n_38), .A2(p_15[4]), .ZN(n_99));
   NOR2_X1 i_169 (.A1(n_23), .A2(n_27), .ZN(n_101));
   NAND2_X1 i_170 (.A1(n_29), .A2(n_31), .ZN(n_103));
   NOR2_X1 i_171 (.A1(n_29), .A2(n_31), .ZN(n_105));
   FA_X1 i_172 (.A(p_3[9]), .B(p_15[9]), .CI(n_58), .CO(n_107), .S(n_20));
   FA_X1 i_173 (.A(p_0[9]), .B(p_1[9]), .CI(p_2[9]), .CO(n_109), .S(n_18));
   FA_X1 i_174 (.A(n_51), .B(n_20), .CI(n_18), .CO(n_110), .S(n_22));
   XNOR2_X1 i_175 (.A(n_122), .B(n_111), .ZN(\aggregated_res[14] [9]));
   OAI22_X1 i_176 (.A1(n_57), .A2(n_53), .B1(n_61), .B2(n_65), .ZN(n_111));
   AOI21_X1 i_177 (.A(n_126), .B1(n_55), .B2(n_22), .ZN(n_122));
   NAND2_X1 i_178 (.A1(n_55), .A2(n_22), .ZN(n_124));
   NOR2_X1 i_179 (.A1(n_55), .A2(n_22), .ZN(n_126));
   FA_X1 i_180 (.A(p_0[10]), .B(p_1[10]), .CI(p_2[10]), .CO(n_142), .S(n_24));
   HA_X1 i_181 (.A(n_24), .B(n_110), .CO(n_145), .S(n_30));
   FA_X1 i_182 (.A(p_3[10]), .B(p_4[10]), .CI(p_15[10]), .CO(n_147), .S(n_26));
   FA_X1 i_183 (.A(n_109), .B(n_107), .CI(n_26), .CO(n_149), .S(n_28));
   XOR2_X1 i_184 (.A(n_157), .B(n_151), .Z(\aggregated_res[14] [10]));
   OAI21_X1 i_185 (.A(n_153), .B1(n_30), .B2(n_28), .ZN(n_151));
   NAND2_X1 i_186 (.A1(n_30), .A2(n_28), .ZN(n_153));
   NOR2_X1 i_187 (.A1(n_30), .A2(n_28), .ZN(n_155));
   NAND2_X1 i_188 (.A1(n_181), .A2(n_159), .ZN(n_157));
   OAI211_X1 i_189 (.A(n_63), .B(n_124), .C1(n_178), .C2(n_161), .ZN(n_159));
   OAI21_X1 i_190 (.A(n_183), .B1(n_53), .B2(n_57), .ZN(n_161));
   INV_X1 i_191 (.A(n_179), .ZN(n_178));
   OAI211_X1 i_192 (.A(n_71), .B(n_103), .C1(n_73), .C2(n_101), .ZN(n_179));
   INV_X1 i_193 (.A(n_126), .ZN(n_181));
   INV_X1 i_194 (.A(n_105), .ZN(n_183));
   FA_X1 i_195 (.A(p_3[11]), .B(p_4[11]), .CI(p_15[11]), .CO(n_35), .S(n_34));
   FA_X1 i_196 (.A(n_147), .B(n_142), .CI(n_34), .CO(n_37), .S(n_36));
   FA_X1 i_197 (.A(p_0[11]), .B(p_1[11]), .CI(p_2[11]), .CO(n_33), .S(n_32));
   FA_X1 i_198 (.A(n_32), .B(n_149), .CI(n_36), .CO(n_39), .S(n_185));
   HA_X1 i_199 (.A(n_37), .B(n_39), .CO(n_187), .S(n_48));
   FA_X1 i_200 (.A(p_3[12]), .B(p_4[12]), .CI(p_5[12]), .CO(n_43), .S(n_42));
   FA_X1 i_201 (.A(p_0[12]), .B(p_1[12]), .CI(p_2[12]), .CO(n_41), .S(n_40));
   FA_X1 i_202 (.A(p_15[12]), .B(n_35), .CI(n_33), .CO(n_45), .S(n_44));
   FA_X1 i_203 (.A(n_42), .B(n_40), .CI(n_44), .CO(n_47), .S(n_46));
   FA_X1 i_204 (.A(p_15[13]), .B(n_43), .CI(n_41), .CO(n_189), .S(n_54));
   FA_X1 i_205 (.A(p_3[13]), .B(p_4[13]), .CI(p_5[13]), .CO(n_191), .S(n_52));
   FA_X1 i_206 (.A(p_0[13]), .B(p_1[13]), .CI(p_2[13]), .CO(n_193), .S(n_50));
   FA_X1 i_207 (.A(n_45), .B(n_52), .CI(n_50), .CO(n_195), .S(n_56));
   FA_X1 i_208 (.A(n_54), .B(n_47), .CI(n_56), .CO(n_198), .S(n_197));
   XOR2_X1 i_209 (.A(n_262), .B(n_199), .Z(\aggregated_res[14] [13]));
   OAI21_X1 i_210 (.A(n_241), .B1(n_187), .B2(n_197), .ZN(n_199));
   NAND2_X1 i_211 (.A1(n_187), .A2(n_197), .ZN(n_241));
   OAI21_X1 i_212 (.A(n_275), .B1(n_267), .B2(n_265), .ZN(n_262));
   INV_X1 i_213 (.A(n_265), .ZN(n_263));
   NOR2_X1 i_214 (.A1(n_279), .A2(n_277), .ZN(n_265));
   NOR2_X1 i_215 (.A1(n_271), .A2(n_269), .ZN(n_267));
   AOI21_X1 i_216 (.A(n_273), .B1(n_185), .B2(n_145), .ZN(n_269));
   NOR2_X1 i_217 (.A1(n_185), .A2(n_145), .ZN(n_271));
   AOI21_X1 i_218 (.A(n_155), .B1(n_157), .B2(n_153), .ZN(n_273));
   NAND2_X1 i_219 (.A1(n_279), .A2(n_277), .ZN(n_275));
   INV_X1 i_220 (.A(n_46), .ZN(n_277));
   INV_X1 i_221 (.A(n_48), .ZN(n_279));
   FA_X1 i_222 (.A(p_6[14]), .B(p_15[14]), .CI(n_191), .CO(n_281), .S(n_64));
   FA_X1 i_223 (.A(n_193), .B(n_189), .CI(n_64), .CO(n_283), .S(n_66));
   FA_X1 i_224 (.A(p_3[14]), .B(p_4[14]), .CI(p_5[14]), .CO(n_285), .S(n_62));
   FA_X1 i_225 (.A(p_0[14]), .B(p_1[14]), .CI(p_2[14]), .CO(n_286), .S(n_60));
   FA_X1 i_226 (.A(n_62), .B(n_60), .CI(n_195), .CO(n_287), .S(n_68));
   HA_X1 i_227 (.A(n_66), .B(n_68), .CO(n_310), .S(n_70));
   OAI21_X1 i_228 (.A(n_367), .B1(n_198), .B2(n_70), .ZN(n_363));
   NOR2_X1 i_229 (.A1(n_198), .A2(n_70), .ZN(n_365));
   NAND2_X1 i_230 (.A1(n_198), .A2(n_70), .ZN(n_367));
   FA_X1 i_231 (.A(p_6[15]), .B(p_15[15]), .CI(n_285), .CO(n_369), .S(n_76));
   FA_X1 i_232 (.A(n_286), .B(n_281), .CI(n_76), .CO(n_371), .S(n_78));
   FA_X1 i_233 (.A(p_3[15]), .B(p_4[15]), .CI(p_5[15]), .CO(n_373), .S(n_74));
   FA_X1 i_234 (.A(p_0[15]), .B(p_1[15]), .CI(p_2[15]), .CO(n_375), .S(n_72));
   FA_X1 i_235 (.A(n_74), .B(n_72), .CI(n_283), .CO(n_377), .S(n_80));
   FA_X1 i_236 (.A(n_78), .B(n_287), .CI(n_80), .CO(n_379), .S(n_82));
   XNOR2_X1 i_237 (.A(n_383), .B(n_381), .ZN(\aggregated_res[14] [15]));
   AOI21_X1 i_238 (.A(n_391), .B1(n_310), .B2(n_82), .ZN(n_381));
   INV_X1 i_239 (.A(n_385), .ZN(n_383));
   OAI21_X1 i_240 (.A(n_367), .B1(n_365), .B2(n_387), .ZN(n_385));
   OAI21_X1 i_241 (.A(n_389), .B1(n_187), .B2(n_197), .ZN(n_387));
   NAND2_X1 i_242 (.A1(n_262), .A2(n_241), .ZN(n_389));
   NAND2_X1 i_243 (.A1(n_310), .A2(n_82), .ZN(n_390));
   NOR2_X1 i_244 (.A1(n_310), .A2(n_82), .ZN(n_391));
   FA_X1 i_245 (.A(p_6[17]), .B(p_7[17]), .CI(p_15[17]), .CO(n_393), .S(n_102));
   FA_X1 i_246 (.A(p_3[17]), .B(p_4[17]), .CI(p_5[17]), .CO(n_395), .S(n_100));
   FA_X1 i_247 (.A(p_0[17]), .B(p_1[17]), .CI(p_2[17]), .CO(n_397), .S(n_98));
   FA_X1 i_248 (.A(n_102), .B(n_100), .CI(n_98), .CO(n_399), .S(n_106));
   FA_X1 i_249 (.A(n_373), .B(n_375), .CI(n_369), .CO(n_91), .S(n_90));
   FA_X1 i_250 (.A(n_90), .B(n_371), .CI(n_377), .CO(n_95), .S(n_94));
   FA_X1 i_251 (.A(p_6[16]), .B(p_7[16]), .CI(p_15[16]), .CO(n_89), .S(n_88));
   FA_X1 i_252 (.A(p_3[16]), .B(p_4[16]), .CI(p_5[16]), .CO(n_87), .S(n_86));
   FA_X1 i_253 (.A(p_0[16]), .B(p_1[16]), .CI(p_2[16]), .CO(n_85), .S(n_84));
   FA_X1 i_254 (.A(n_89), .B(n_87), .CI(n_85), .CO(n_401), .S(n_104));
   FA_X1 i_255 (.A(n_88), .B(n_86), .CI(n_84), .CO(n_93), .S(n_92));
   FA_X1 i_256 (.A(n_91), .B(n_104), .CI(n_93), .CO(n_403), .S(n_108));
   FA_X1 i_257 (.A(n_106), .B(n_95), .CI(n_108), .CO(n_407), .S(n_405));
   HA_X1 i_258 (.A(n_92), .B(n_94), .CO(n_411), .S(n_409));
   XOR2_X1 i_259 (.A(n_415), .B(n_413), .Z(\aggregated_res[14] [17]));
   OAI22_X1 i_260 (.A1(n_409), .A2(n_379), .B1(n_418), .B2(n_417), .ZN(n_413));
   OAI21_X1 i_261 (.A(n_421), .B1(n_405), .B2(n_411), .ZN(n_415));
   AOI21_X1 i_262 (.A(n_391), .B1(n_423), .B2(n_390), .ZN(n_417));
   INV_X1 i_263 (.A(n_419), .ZN(n_418));
   NAND2_X1 i_264 (.A1(n_409), .A2(n_379), .ZN(n_419));
   NAND2_X1 i_265 (.A1(n_405), .A2(n_411), .ZN(n_421));
   INV_X1 i_266 (.A(n_385), .ZN(n_423));
   FA_X1 i_267 (.A(p_3[19]), .B(p_4[19]), .CI(p_5[19]), .CO(n_131), .S(n_130));
   FA_X1 i_268 (.A(p_0[19]), .B(p_1[19]), .CI(p_2[19]), .CO(n_129), .S(n_128));
   FA_X1 i_269 (.A(p_6[18]), .B(p_7[18]), .CI(p_8[18]), .CO(n_117), .S(n_116));
   FA_X1 i_270 (.A(p_3[18]), .B(p_4[18]), .CI(p_5[18]), .CO(n_115), .S(n_114));
   FA_X1 i_271 (.A(p_15[19]), .B(n_117), .CI(n_115), .CO(n_135), .S(n_134));
   FA_X1 i_272 (.A(n_130), .B(n_128), .CI(n_134), .CO(n_139), .S(n_138));
   FA_X1 i_273 (.A(n_397), .B(n_401), .CI(n_116), .CO(n_121), .S(n_120));
   FA_X1 i_274 (.A(n_399), .B(n_120), .CI(n_403), .CO(n_125), .S(n_425));
   FA_X1 i_275 (.A(p_0[18]), .B(p_1[18]), .CI(p_2[18]), .CO(n_113), .S(n_112));
   FA_X1 i_276 (.A(p_15[18]), .B(n_393), .CI(n_395), .CO(n_119), .S(n_118));
   FA_X1 i_277 (.A(p_6[19]), .B(p_7[19]), .CI(p_8[19]), .CO(n_133), .S(n_132));
   FA_X1 i_278 (.A(n_113), .B(n_119), .CI(n_132), .CO(n_137), .S(n_136));
   FA_X1 i_279 (.A(n_114), .B(n_112), .CI(n_118), .CO(n_123), .S(n_427));
   FA_X1 i_280 (.A(n_121), .B(n_136), .CI(n_123), .CO(n_141), .S(n_140));
   FA_X1 i_281 (.A(n_138), .B(n_125), .CI(n_140), .CO(n_143), .S(n_429));
   FA_X1 i_282 (.A(p_0[20]), .B(p_1[20]), .CI(p_2[20]), .CO(n_431), .S(n_144));
   FA_X1 i_283 (.A(n_131), .B(n_129), .CI(n_135), .CO(n_433), .S(n_152));
   FA_X1 i_284 (.A(n_144), .B(n_152), .CI(n_137), .CO(n_435), .S(n_156));
   FA_X1 i_285 (.A(p_9[20]), .B(p_15[20]), .CI(n_133), .CO(n_437), .S(n_150));
   FA_X1 i_286 (.A(p_6[20]), .B(p_7[20]), .CI(p_8[20]), .CO(n_439), .S(n_148));
   FA_X1 i_287 (.A(p_3[20]), .B(p_4[20]), .CI(p_5[20]), .CO(n_441), .S(n_146));
   FA_X1 i_288 (.A(n_150), .B(n_148), .CI(n_146), .CO(n_443), .S(n_154));
   FA_X1 i_289 (.A(n_139), .B(n_154), .CI(n_141), .CO(n_445), .S(n_158));
   HA_X1 i_290 (.A(n_156), .B(n_158), .CO(n_447), .S(n_160));
   NAND2_X1 i_291 (.A1(n_453), .A2(n_451), .ZN(n_449));
   NAND2_X1 i_292 (.A1(n_143), .A2(n_160), .ZN(n_451));
   OR2_X1 i_293 (.A1(n_143), .A2(n_160), .ZN(n_453));
   FA_X1 i_294 (.A(p_0[21]), .B(p_1[21]), .CI(p_2[21]), .CO(n_163), .S(n_162));
   FA_X1 i_295 (.A(n_441), .B(n_431), .CI(n_437), .CO(n_171), .S(n_170));
   FA_X1 i_296 (.A(n_162), .B(n_433), .CI(n_170), .CO(n_175), .S(n_174));
   FA_X1 i_297 (.A(p_9[21]), .B(p_15[21]), .CI(n_439), .CO(n_169), .S(n_168));
   FA_X1 i_298 (.A(p_6[21]), .B(p_7[21]), .CI(p_8[21]), .CO(n_167), .S(n_166));
   FA_X1 i_299 (.A(p_3[21]), .B(p_4[21]), .CI(p_5[21]), .CO(n_165), .S(n_164));
   FA_X1 i_300 (.A(n_168), .B(n_166), .CI(n_164), .CO(n_173), .S(n_172));
   FA_X1 i_301 (.A(n_443), .B(n_435), .CI(n_172), .CO(n_177), .S(n_176));
   FA_X1 i_302 (.A(n_174), .B(n_445), .CI(n_176), .CO(n_457), .S(n_455));
   HA_X1 i_303 (.A(n_427), .B(n_425), .CO(n_127), .S(n_459));
   FA_X1 i_304 (.A(p_3[22]), .B(p_4[22]), .CI(p_5[22]), .CO(n_461), .S(n_182));
   FA_X1 i_305 (.A(p_0[22]), .B(p_1[22]), .CI(p_2[22]), .CO(n_463), .S(n_180));
   FA_X1 i_306 (.A(n_182), .B(n_180), .CI(n_171), .CO(n_465), .S(n_192));
   FA_X1 i_307 (.A(p_9[22]), .B(p_10[22]), .CI(p_15[22]), .CO(n_467), .S(n_186));
   FA_X1 i_308 (.A(p_6[22]), .B(p_7[22]), .CI(p_8[22]), .CO(n_469), .S(n_184));
   FA_X1 i_309 (.A(n_169), .B(n_186), .CI(n_184), .CO(n_471), .S(n_190));
   FA_X1 i_310 (.A(n_167), .B(n_165), .CI(n_163), .CO(n_472), .S(n_188));
   FA_X1 i_311 (.A(n_188), .B(n_173), .CI(n_175), .CO(n_473), .S(n_194));
   FA_X1 i_312 (.A(n_192), .B(n_190), .CI(n_194), .CO(n_498), .S(n_196));
   HA_X1 i_313 (.A(n_177), .B(n_196), .CO(n_503), .S(n_501));
   XNOR2_X1 i_314 (.A(n_509), .B(n_505), .ZN(\aggregated_res[14] [22]));
   OAI21_X1 i_315 (.A(n_511), .B1(n_457), .B2(n_501), .ZN(n_505));
   INV_X1 i_316 (.A(n_509), .ZN(n_507));
   OAI211_X1 i_317 (.A(n_527), .B(n_513), .C1(n_531), .C2(n_515), .ZN(n_509));
   NAND2_X1 i_318 (.A1(n_457), .A2(n_501), .ZN(n_511));
   AOI22_X1 i_319 (.A1(n_455), .A2(n_447), .B1(n_545), .B2(n_541), .ZN(n_513));
   INV_X1 i_320 (.A(n_517), .ZN(n_515));
   AOI21_X1 i_321 (.A(n_519), .B1(n_549), .B2(n_547), .ZN(n_517));
   OAI22_X1 i_322 (.A1(n_411), .A2(n_405), .B1(n_523), .B2(n_521), .ZN(n_519));
   NAND2_X1 i_323 (.A1(n_421), .A2(n_419), .ZN(n_521));
   AOI211_X1 i_324 (.A(n_525), .B(n_391), .C1(n_390), .C2(n_383), .ZN(n_523));
   NOR2_X1 i_325 (.A1(n_409), .A2(n_379), .ZN(n_525));
   INV_X1 i_326 (.A(n_529), .ZN(n_527));
   AOI21_X1 i_327 (.A(n_531), .B1(n_539), .B2(n_537), .ZN(n_529));
   NAND3_X1 i_328 (.A1(n_453), .A2(n_533), .A3(n_541), .ZN(n_531));
   INV_X1 i_329 (.A(n_535), .ZN(n_533));
   NOR2_X1 i_330 (.A1(n_429), .A2(n_127), .ZN(n_535));
   NAND2_X1 i_331 (.A1(n_459), .A2(n_407), .ZN(n_537));
   NAND2_X1 i_332 (.A1(n_429), .A2(n_127), .ZN(n_539));
   INV_X1 i_333 (.A(n_543), .ZN(n_541));
   NOR2_X1 i_334 (.A1(n_455), .A2(n_447), .ZN(n_543));
   INV_X1 i_335 (.A(n_451), .ZN(n_545));
   INV_X1 i_336 (.A(n_407), .ZN(n_547));
   INV_X1 i_337 (.A(n_459), .ZN(n_549));
   FA_X1 i_338 (.A(p_15[25]), .B(n_227), .CI(n_225), .CO(n_251), .S(n_250));
   FA_X1 i_339 (.A(n_226), .B(n_224), .CI(n_222), .CO(n_233), .S(n_232));
   FA_X1 i_340 (.A(n_220), .B(n_230), .CI(n_228), .CO(n_235), .S(n_234));
   FA_X1 i_341 (.A(n_250), .B(n_233), .CI(n_235), .CO(n_259), .S(n_258));
   FA_X1 i_342 (.A(n_213), .B(n_211), .CI(n_215), .CO(n_237), .S(n_236));
   FA_X1 i_343 (.A(n_232), .B(n_236), .CI(n_234), .CO(n_239), .S(n_238));
   FA_X1 i_344 (.A(n_248), .B(n_246), .CI(n_244), .CO(n_255), .S(n_254));
   FA_X1 i_345 (.A(n_242), .B(n_231), .CI(n_252), .CO(n_257), .S(n_256));
   FA_X1 i_346 (.A(n_254), .B(n_256), .CI(n_237), .CO(n_261), .S(n_260));
   FA_X1 i_347 (.A(n_258), .B(n_239), .CI(n_260), .CO(n_553), .S(n_551));
   FA_X1 i_348 (.A(n_463), .B(n_472), .CI(n_206), .CO(n_211), .S(n_210));
   FA_X1 i_349 (.A(n_204), .B(n_202), .CI(n_200), .CO(n_213), .S(n_212));
   FA_X1 i_350 (.A(n_210), .B(n_212), .CI(n_473), .CO(n_217), .S(n_216));
   HA_X1 i_351 (.A(n_217), .B(n_238), .CO(n_555), .S(n_240));
   FA_X1 i_352 (.A(n_467), .B(n_469), .CI(n_461), .CO(n_209), .S(n_208));
   FA_X1 i_353 (.A(n_208), .B(n_471), .CI(n_465), .CO(n_215), .S(n_214));
   FA_X1 i_354 (.A(n_214), .B(n_498), .CI(n_216), .CO(n_219), .S(n_218));
   FA_X1 i_355 (.A(p_0[25]), .B(p_1[25]), .CI(p_2[25]), .CO(n_243), .S(n_242));
   FA_X1 i_356 (.A(p_3[23]), .B(p_4[23]), .CI(p_5[23]), .CO(n_203), .S(n_202));
   FA_X1 i_357 (.A(p_0[23]), .B(p_1[23]), .CI(p_2[23]), .CO(n_201), .S(n_200));
   FA_X1 i_358 (.A(n_203), .B(n_201), .CI(n_209), .CO(n_231), .S(n_230));
   FA_X1 i_359 (.A(p_3[24]), .B(p_4[24]), .CI(p_5[24]), .CO(n_223), .S(n_222));
   FA_X1 i_360 (.A(p_0[24]), .B(p_1[24]), .CI(p_2[24]), .CO(n_221), .S(n_220));
   FA_X1 i_361 (.A(p_9[23]), .B(p_10[23]), .CI(p_15[23]), .CO(n_207), .S(n_206));
   FA_X1 i_362 (.A(p_6[23]), .B(p_7[23]), .CI(p_8[23]), .CO(n_205), .S(n_204));
   FA_X1 i_363 (.A(p_15[24]), .B(n_207), .CI(n_205), .CO(n_229), .S(n_228));
   FA_X1 i_364 (.A(n_223), .B(n_221), .CI(n_229), .CO(n_253), .S(n_252));
   FA_X1 i_365 (.A(p_6[26]), .B(p_7[26]), .CI(p_8[26]), .CO(n_557), .S(n_268));
   FA_X1 i_366 (.A(p_3[26]), .B(p_4[26]), .CI(p_5[26]), .CO(n_559), .S(n_266));
   FA_X1 i_367 (.A(p_0[26]), .B(p_1[26]), .CI(p_2[26]), .CO(n_561), .S(n_264));
   FA_X1 i_368 (.A(n_268), .B(n_266), .CI(n_264), .CO(n_563), .S(n_278));
   FA_X1 i_369 (.A(p_9[24]), .B(p_10[24]), .CI(p_11[24]), .CO(n_227), .S(n_226));
   FA_X1 i_370 (.A(p_6[24]), .B(p_7[24]), .CI(p_8[24]), .CO(n_225), .S(n_224));
   FA_X1 i_371 (.A(p_9[25]), .B(p_10[25]), .CI(p_11[25]), .CO(n_249), .S(n_248));
   FA_X1 i_372 (.A(p_12[26]), .B(p_15[26]), .CI(n_249), .CO(n_565), .S(n_272));
   FA_X1 i_373 (.A(p_9[26]), .B(p_10[26]), .CI(p_11[26]), .CO(n_567), .S(n_270));
   FA_X1 i_374 (.A(n_251), .B(n_272), .CI(n_270), .CO(n_569), .S(n_276));
   FA_X1 i_375 (.A(n_257), .B(n_278), .CI(n_276), .CO(n_571), .S(n_282));
   FA_X1 i_376 (.A(p_6[25]), .B(p_7[25]), .CI(p_8[25]), .CO(n_247), .S(n_246));
   FA_X1 i_377 (.A(p_3[25]), .B(p_4[25]), .CI(p_5[25]), .CO(n_245), .S(n_244));
   FA_X1 i_378 (.A(n_247), .B(n_245), .CI(n_243), .CO(n_572), .S(n_274));
   FA_X1 i_379 (.A(n_253), .B(n_274), .CI(n_255), .CO(n_573), .S(n_280));
   FA_X1 i_380 (.A(n_259), .B(n_280), .CI(n_261), .CO(n_588), .S(n_284));
   HA_X1 i_381 (.A(n_282), .B(n_284), .CO(n_592), .S(n_590));
   XNOR2_X1 i_382 (.A(n_616), .B(n_594), .ZN(\aggregated_res[14] [26]));
   OAI21_X1 i_383 (.A(n_614), .B1(n_553), .B2(n_590), .ZN(n_594));
   NAND2_X1 i_384 (.A1(n_553), .A2(n_590), .ZN(n_614));
   OAI21_X1 i_385 (.A(n_639), .B1(n_507), .B2(n_617), .ZN(n_616));
   OR2_X1 i_386 (.A1(n_645), .A2(n_636), .ZN(n_617));
   NOR2_X1 i_387 (.A1(n_501), .A2(n_457), .ZN(n_636));
   INV_X1 i_388 (.A(n_641), .ZN(n_639));
   OAI22_X1 i_389 (.A1(n_647), .A2(n_645), .B1(n_661), .B2(n_643), .ZN(n_641));
   AOI21_X1 i_390 (.A(n_649), .B1(n_551), .B2(n_555), .ZN(n_643));
   OR3_X1 i_391 (.A1(n_661), .A2(n_655), .A3(n_659), .ZN(n_645));
   AND2_X1 i_392 (.A1(n_511), .A2(n_651), .ZN(n_647));
   AND2_X1 i_393 (.A1(n_240), .A2(n_219), .ZN(n_649));
   NAND2_X1 i_394 (.A1(n_503), .A2(n_218), .ZN(n_651));
   INV_X1 i_395 (.A(n_655), .ZN(n_653));
   NOR2_X1 i_396 (.A1(n_503), .A2(n_218), .ZN(n_655));
   INV_X1 i_397 (.A(n_659), .ZN(n_657));
   NOR2_X1 i_398 (.A1(n_240), .A2(n_219), .ZN(n_659));
   NOR2_X1 i_399 (.A1(n_551), .A2(n_555), .ZN(n_661));
   FA_X1 i_400 (.A(n_314), .B(n_312), .CI(n_322), .CO(n_329), .S(n_328));
   FA_X1 i_401 (.A(n_340), .B(n_338), .CI(n_325), .CO(n_355), .S(n_354));
   FA_X1 i_402 (.A(n_346), .B(n_344), .CI(n_342), .CO(n_353), .S(n_352));
   FA_X1 i_403 (.A(n_329), .B(n_354), .CI(n_352), .CO(n_359), .S(n_358));
   FA_X1 i_404 (.A(n_569), .B(n_300), .CI(n_573), .CO(n_307), .S(n_306));
   FA_X1 i_405 (.A(n_303), .B(n_301), .CI(n_324), .CO(n_331), .S(n_330));
   FA_X1 i_406 (.A(n_302), .B(n_304), .CI(n_571), .CO(n_309), .S(n_308));
   FA_X1 i_407 (.A(n_307), .B(n_330), .CI(n_309), .CO(n_335), .S(n_334));
   FA_X1 i_408 (.A(n_350), .B(n_348), .CI(n_327), .CO(n_357), .S(n_356));
   FA_X1 i_409 (.A(n_305), .B(n_328), .CI(n_326), .CO(n_333), .S(n_332));
   FA_X1 i_410 (.A(n_331), .B(n_356), .CI(n_333), .CO(n_361), .S(n_360));
   FA_X1 i_411 (.A(n_358), .B(n_335), .CI(n_360), .CO(n_663), .S(n_362));
   FA_X1 i_412 (.A(n_288), .B(n_298), .CI(n_563), .CO(n_305), .S(n_304));
   FA_X1 i_413 (.A(n_320), .B(n_318), .CI(n_316), .CO(n_327), .S(n_326));
   HA_X1 i_414 (.A(n_332), .B(n_334), .CO(n_337), .S(n_336));
   FA_X1 i_415 (.A(n_572), .B(n_565), .CI(n_296), .CO(n_301), .S(n_300));
   FA_X1 i_416 (.A(n_294), .B(n_292), .CI(n_290), .CO(n_303), .S(n_302));
   FA_X1 i_417 (.A(n_306), .B(n_588), .CI(n_308), .CO(n_311), .S(n_665));
   FA_X1 i_418 (.A(p_6[30]), .B(p_7[30]), .CI(p_8[30]), .CO(n_667), .S(n_368));
   FA_X1 i_419 (.A(p_3[30]), .B(p_4[30]), .CI(p_5[30]), .CO(n_669), .S(n_366));
   FA_X1 i_420 (.A(p_0[30]), .B(p_1[30]), .CI(p_2[30]), .CO(n_671), .S(n_364));
   FA_X1 i_421 (.A(n_368), .B(n_366), .CI(n_364), .CO(n_673), .S(n_380));
   FA_X1 i_422 (.A(p_12[28]), .B(p_13[28]), .CI(p_15[28]), .CO(n_321), .S(n_320));
   FA_X1 i_423 (.A(p_9[28]), .B(p_10[28]), .CI(p_11[28]), .CO(n_319), .S(n_318));
   FA_X1 i_424 (.A(p_6[28]), .B(p_7[28]), .CI(p_8[28]), .CO(n_317), .S(n_316));
   FA_X1 i_425 (.A(n_321), .B(n_319), .CI(n_317), .CO(n_349), .S(n_348));
   FA_X1 i_426 (.A(p_12[30]), .B(p_13[30]), .CI(p_14[30]), .CO(n_675), .S(n_372));
   FA_X1 i_427 (.A(p_9[30]), .B(p_10[30]), .CI(p_11[30]), .CO(n_677), .S(n_370));
   FA_X1 i_428 (.A(n_349), .B(n_372), .CI(n_370), .CO(n_679), .S(n_378));
   FA_X1 i_429 (.A(p_3[28]), .B(p_4[28]), .CI(p_5[28]), .CO(n_315), .S(n_314));
   FA_X1 i_430 (.A(p_0[28]), .B(p_1[28]), .CI(p_2[28]), .CO(n_313), .S(n_312));
   FA_X1 i_431 (.A(p_9[27]), .B(p_10[27]), .CI(p_11[27]), .CO(n_295), .S(n_294));
   FA_X1 i_432 (.A(p_6[27]), .B(p_7[27]), .CI(p_8[27]), .CO(n_293), .S(n_292));
   FA_X1 i_433 (.A(p_3[27]), .B(p_4[27]), .CI(p_5[27]), .CO(n_291), .S(n_290));
   FA_X1 i_434 (.A(n_295), .B(n_293), .CI(n_291), .CO(n_323), .S(n_322));
   FA_X1 i_435 (.A(n_315), .B(n_313), .CI(n_323), .CO(n_351), .S(n_350));
   FA_X1 i_436 (.A(p_6[29]), .B(p_7[29]), .CI(p_8[29]), .CO(n_343), .S(n_342));
   FA_X1 i_437 (.A(p_3[29]), .B(p_4[29]), .CI(p_5[29]), .CO(n_341), .S(n_340));
   FA_X1 i_438 (.A(p_0[29]), .B(p_1[29]), .CI(p_2[29]), .CO(n_339), .S(n_338));
   FA_X1 i_439 (.A(n_343), .B(n_341), .CI(n_339), .CO(n_681), .S(n_376));
   FA_X1 i_440 (.A(p_12[29]), .B(p_13[29]), .CI(p_15[29]), .CO(n_347), .S(n_346));
   FA_X1 i_441 (.A(p_9[29]), .B(p_10[29]), .CI(p_11[29]), .CO(n_345), .S(n_344));
   FA_X1 i_442 (.A(p_15[30]), .B(n_347), .CI(n_345), .CO(n_683), .S(n_374));
   FA_X1 i_443 (.A(n_351), .B(n_376), .CI(n_374), .CO(n_685), .S(n_382));
   FA_X1 i_444 (.A(n_380), .B(n_378), .CI(n_382), .CO(n_687), .S(n_386));
   FA_X1 i_445 (.A(p_0[27]), .B(p_1[27]), .CI(p_2[27]), .CO(n_289), .S(n_288));
   FA_X1 i_446 (.A(n_557), .B(n_559), .CI(n_561), .CO(n_299), .S(n_298));
   FA_X1 i_447 (.A(p_12[27]), .B(p_15[27]), .CI(n_567), .CO(n_297), .S(n_296));
   FA_X1 i_448 (.A(n_289), .B(n_299), .CI(n_297), .CO(n_325), .S(n_324));
   FA_X1 i_449 (.A(n_353), .B(n_355), .CI(n_357), .CO(n_689), .S(n_384));
   FA_X1 i_450 (.A(n_359), .B(n_384), .CI(n_361), .CO(n_691), .S(n_388));
   HA_X1 i_451 (.A(n_386), .B(n_388), .CO(n_711), .S(n_693));
   XNOR2_X1 i_452 (.A(n_717), .B(n_712), .ZN(\aggregated_res[14] [30]));
   OAI21_X1 i_453 (.A(n_715), .B1(n_663), .B2(n_693), .ZN(n_712));
   NAND2_X1 i_454 (.A1(n_663), .A2(n_693), .ZN(n_715));
   OAI21_X1 i_455 (.A(n_721), .B1(n_738), .B2(n_719), .ZN(n_717));
   NAND2_X1 i_456 (.A1(n_616), .A2(n_735), .ZN(n_719));
   INV_X1 i_457 (.A(n_723), .ZN(n_721));
   OAI211_X1 i_458 (.A(n_729), .B(n_725), .C1(n_767), .C2(n_727), .ZN(n_723));
   OAI21_X1 i_459 (.A(n_737), .B1(n_769), .B2(n_731), .ZN(n_725));
   NAND2_X1 i_460 (.A1(n_336), .A2(n_311), .ZN(n_727));
   NAND2_X1 i_461 (.A1(n_362), .A2(n_337), .ZN(n_729));
   INV_X1 i_462 (.A(n_733), .ZN(n_731));
   NAND2_X1 i_463 (.A1(n_665), .A2(n_592), .ZN(n_733));
   OR2_X1 i_464 (.A1(n_590), .A2(n_553), .ZN(n_735));
   INV_X1 i_465 (.A(n_738), .ZN(n_737));
   OAI211_X1 i_466 (.A(n_739), .B(n_765), .C1(n_665), .C2(n_592), .ZN(n_738));
   INV_X1 i_467 (.A(n_752), .ZN(n_739));
   NOR2_X1 i_468 (.A1(n_336), .A2(n_311), .ZN(n_752));
   INV_X1 i_469 (.A(n_767), .ZN(n_765));
   NOR2_X1 i_470 (.A1(n_362), .A2(n_337), .ZN(n_767));
   INV_X1 i_471 (.A(n_614), .ZN(n_769));
   FA_X1 i_472 (.A(p_9[31]), .B(p_10[31]), .CI(p_11[31]), .CO(n_771), .S(n_398));
   FA_X1 i_473 (.A(p_6[31]), .B(p_7[31]), .CI(p_8[31]), .CO(n_773), .S(n_396));
   FA_X1 i_474 (.A(p_3[31]), .B(p_4[31]), .CI(p_5[31]), .CO(n_775), .S(n_394));
   FA_X1 i_475 (.A(n_398), .B(n_396), .CI(n_394), .CO(n_776), .S(n_408));
   FA_X1 i_476 (.A(n_685), .B(n_408), .CI(n_689), .CO(n_777), .S(n_414));
   FA_X1 i_477 (.A(p_12[31]), .B(p_13[31]), .CI(p_14[31]), .CO(n_779), .S(n_400));
   FA_X1 i_478 (.A(n_681), .B(n_683), .CI(n_400), .CO(n_781), .S(n_406));
   FA_X1 i_479 (.A(n_673), .B(n_679), .CI(n_406), .CO(n_783), .S(n_412));
   FA_X1 i_480 (.A(p_0[31]), .B(p_1[31]), .CI(p_2[31]), .CO(n_785), .S(n_392));
   FA_X1 i_481 (.A(n_667), .B(n_669), .CI(n_671), .CO(n_786), .S(n_404));
   FA_X1 i_482 (.A(p_15[31]), .B(n_675), .CI(n_677), .CO(n_787), .S(n_402));
   FA_X1 i_483 (.A(n_392), .B(n_404), .CI(n_402), .CO(n_789), .S(n_410));
   FA_X1 i_484 (.A(n_412), .B(n_410), .CI(n_687), .CO(n_791), .S(n_416));
   FA_X1 i_485 (.A(n_414), .B(n_691), .CI(n_416), .CO(n_795), .S(n_793));
   OAI21_X1 i_486 (.A(n_717), .B1(n_663), .B2(n_693), .ZN(n_797));
   NAND2_X1 i_487 (.A1(n_797), .A2(n_715), .ZN(n_799));
   NAND2_X1 i_488 (.A1(n_793), .A2(n_711), .ZN(n_801));
   INV_X1 i_489 (.A(n_801), .ZN(n_803));
   OAI21_X1 i_490 (.A(n_801), .B1(n_793), .B2(n_711), .ZN(n_805));
   XNOR2_X1 i_491 (.A(n_799), .B(n_805), .ZN(\aggregated_res[14] [31]));
   FA_X1 i_492 (.A(n_785), .B(n_786), .CI(n_787), .CO(n_807), .S(n_430));
   FA_X1 i_493 (.A(p_5[32]), .B(p_6[32]), .CI(p_7[32]), .CO(n_809), .S(n_422));
   FA_X1 i_494 (.A(p_2[32]), .B(p_3[32]), .CI(p_4[32]), .CO(n_811), .S(n_420));
   FA_X1 i_495 (.A(n_422), .B(n_420), .CI(n_910), .CO(n_812), .S(n_434));
   FA_X1 i_496 (.A(n_430), .B(n_789), .CI(n_434), .CO(n_813), .S(n_438));
   FA_X1 i_497 (.A(p_11[32]), .B(p_12[32]), .CI(p_13[32]), .CO(n_814), .S(n_426));
   FA_X1 i_498 (.A(p_8[32]), .B(p_9[32]), .CI(p_10[32]), .CO(n_818), .S(n_424));
   FA_X1 i_499 (.A(n_907), .B(n_426), .CI(n_424), .CO(n_822), .S(n_432));
   FA_X1 i_500 (.A(n_771), .B(n_773), .CI(n_775), .CO(n_828), .S(n_428));
   FA_X1 i_501 (.A(n_428), .B(n_776), .CI(n_781), .CO(n_829), .S(n_436));
   FA_X1 i_502 (.A(n_432), .B(n_783), .CI(n_436), .CO(n_831), .S(n_440));
   FA_X1 i_503 (.A(n_777), .B(n_438), .CI(n_440), .CO(n_832), .S(n_442));
   HA_X1 i_504 (.A(n_791), .B(n_442), .CO(n_833), .S(n_444));
   XNOR2_X1 i_505 (.A(p_15[32]), .B(n_835), .ZN(n_907));
   XOR2_X1 i_506 (.A(n_779), .B(p_14[32]), .Z(n_835));
   OAI21_X1 i_507 (.A(n_846), .B1(n_856), .B2(n_854), .ZN(n_910));
   XOR2_X1 i_508 (.A(n_839), .B(n_836), .Z(\aggregated_res[14] [32]));
   NAND2_X1 i_509 (.A1(n_844), .A2(n_841), .ZN(n_836));
   OAI22_X1 i_510 (.A1(n_793), .A2(n_711), .B1(n_799), .B2(n_803), .ZN(n_839));
   NAND2_X1 i_511 (.A1(n_795), .A2(n_444), .ZN(n_841));
   OR2_X1 i_512 (.A1(n_795), .A2(n_444), .ZN(n_844));
   NAND2_X1 i_513 (.A1(n_856), .A2(n_854), .ZN(n_846));
   INV_X1 i_514 (.A(p_15[32]), .ZN(n_851));
   INV_X1 i_515 (.A(p_1[32]), .ZN(n_854));
   INV_X1 i_516 (.A(p_0[32]), .ZN(n_856));
   FA_X1 i_517 (.A(p_11[33]), .B(p_12[33]), .CI(p_13[33]), .CO(n_859), .S(n_452));
   FA_X1 i_518 (.A(n_828), .B(n_905), .CI(n_452), .CO(n_861), .S(n_458));
   FA_X1 i_519 (.A(p_8[33]), .B(p_9[33]), .CI(p_10[33]), .CO(n_864), .S(n_450));
   FA_X1 i_520 (.A(p_5[33]), .B(p_6[33]), .CI(p_7[33]), .CO(n_866), .S(n_448));
   FA_X1 i_521 (.A(p_2[33]), .B(p_3[33]), .CI(p_4[33]), .CO(n_871), .S(n_446));
   FA_X1 i_522 (.A(n_450), .B(n_448), .CI(n_446), .CO(n_874), .S(n_460));
   FA_X1 i_523 (.A(n_458), .B(n_829), .CI(n_460), .CO(n_876), .S(n_466));
   FA_X1 i_524 (.A(n_809), .B(n_811), .CI(n_846), .CO(n_877), .S(n_456));
   FA_X1 i_525 (.A(n_903), .B(n_807), .CI(n_456), .CO(n_879), .S(n_462));
   FA_X1 i_526 (.A(p_14[33]), .B(n_814), .CI(n_818), .CO(n_881), .S(n_454));
   FA_X1 i_527 (.A(n_454), .B(n_812), .CI(n_822), .CO(n_884), .S(n_464));
   FA_X1 i_528 (.A(n_462), .B(n_464), .CI(n_813), .CO(n_886), .S(n_468));
   FA_X1 i_529 (.A(n_466), .B(n_831), .CI(n_468), .CO(n_891), .S(n_470));
   HA_X1 i_530 (.A(n_832), .B(n_470), .CO(n_896), .S(n_894));
   OAI21_X1 i_531 (.A(n_909), .B1(n_917), .B2(n_916), .ZN(n_903));
   NAND2_X1 i_532 (.A1(n_901), .A2(n_899), .ZN(n_905));
   OAI21_X1 i_533 (.A(p_14[32]), .B1(n_851), .B2(n_779), .ZN(n_899));
   NAND2_X1 i_534 (.A1(n_851), .A2(n_779), .ZN(n_901));
   XNOR2_X1 i_535 (.A(n_906), .B(n_904), .ZN(\aggregated_res[14] [33]));
   AOI21_X1 i_536 (.A(n_911), .B1(n_839), .B2(n_841), .ZN(n_904));
   OAI21_X1 i_537 (.A(n_908), .B1(n_894), .B2(n_833), .ZN(n_906));
   NAND2_X1 i_538 (.A1(n_894), .A2(n_833), .ZN(n_908));
   NAND2_X1 i_539 (.A1(n_917), .A2(n_916), .ZN(n_909));
   INV_X1 i_540 (.A(n_844), .ZN(n_911));
   INV_X1 i_541 (.A(p_1[33]), .ZN(n_916));
   INV_X1 i_542 (.A(p_0[33]), .ZN(n_917));
   FA_X1 i_543 (.A(n_861), .B(n_884), .CI(n_879), .CO(n_493), .S(n_492));
   FA_X1 i_544 (.A(n_876), .B(n_492), .CI(n_886), .CO(n_497), .S(n_496));
   FA_X1 i_545 (.A(p_12[34]), .B(p_13[34]), .CI(p_14[34]), .CO(n_481), .S(n_480));
   FA_X1 i_546 (.A(p_9[34]), .B(p_10[34]), .CI(p_11[34]), .CO(n_479), .S(n_478));
   FA_X1 i_547 (.A(n_881), .B(n_480), .CI(n_478), .CO(n_487), .S(n_486));
   FA_X1 i_548 (.A(n_871), .B(n_909), .CI(n_877), .CO(n_485), .S(n_484));
   FA_X1 i_549 (.A(n_859), .B(n_864), .CI(n_866), .CO(n_483), .S(n_482));
   FA_X1 i_550 (.A(n_484), .B(n_482), .CI(n_874), .CO(n_491), .S(n_490));
   FA_X1 i_551 (.A(p_3[35]), .B(p_4[35]), .CI(p_5[35]), .CO(n_919), .S(n_500));
   FA_X1 i_552 (.A(n_500), .B(n_898), .CI(n_485), .CO(n_920), .S(n_514));
   FA_X1 i_553 (.A(n_487), .B(n_491), .CI(n_514), .CO(n_921), .S(n_518));
   FA_X1 i_554 (.A(p_6[34]), .B(p_7[34]), .CI(p_8[34]), .CO(n_477), .S(n_476));
   FA_X1 i_555 (.A(p_3[34]), .B(p_4[34]), .CI(p_5[34]), .CO(n_475), .S(n_474));
   FA_X1 i_556 (.A(n_476), .B(n_474), .CI(n_900), .CO(n_489), .S(n_488));
   FA_X1 i_557 (.A(n_488), .B(n_486), .CI(n_490), .CO(n_495), .S(n_494));
   FA_X1 i_558 (.A(p_12[35]), .B(p_13[35]), .CI(p_14[35]), .CO(n_923), .S(n_506));
   FA_X1 i_559 (.A(p_9[35]), .B(p_10[35]), .CI(p_11[35]), .CO(n_924), .S(n_504));
   FA_X1 i_560 (.A(p_6[35]), .B(p_7[35]), .CI(p_8[35]), .CO(n_925), .S(n_502));
   FA_X1 i_561 (.A(n_506), .B(n_504), .CI(n_502), .CO(n_928), .S(n_512));
   FA_X1 i_562 (.A(n_475), .B(n_902), .CI(n_483), .CO(n_929), .S(n_510));
   FA_X1 i_563 (.A(n_481), .B(n_479), .CI(n_477), .CO(n_933), .S(n_508));
   FA_X1 i_564 (.A(n_510), .B(n_508), .CI(n_489), .CO(n_934), .S(n_516));
   FA_X1 i_565 (.A(n_512), .B(n_493), .CI(n_516), .CO(n_935), .S(n_520));
   FA_X1 i_566 (.A(n_518), .B(n_495), .CI(n_520), .CO(n_936), .S(n_522));
   HA_X1 i_567 (.A(n_497), .B(n_522), .CO(n_937), .S(n_524));
   FA_X1 i_568 (.A(n_494), .B(n_496), .CI(n_891), .CO(n_499), .S(n_938));
   AOI21_X1 i_569 (.A(n_939), .B1(n_962), .B2(p_0[34]), .ZN(n_902));
   NOR2_X1 i_570 (.A1(p_2[34]), .A2(n_942), .ZN(n_939));
   XOR2_X1 i_571 (.A(p_2[34]), .B(n_940), .Z(n_900));
   AOI21_X1 i_572 (.A(n_942), .B1(n_962), .B2(p_0[34]), .ZN(n_940));
   NOR2_X1 i_573 (.A1(n_962), .A2(p_0[34]), .ZN(n_942));
   OAI21_X1 i_574 (.A(n_957), .B1(n_963), .B2(n_960), .ZN(n_898));
   NOR2_X1 i_575 (.A1(n_954), .A2(n_945), .ZN(n_944));
   INV_X1 i_576 (.A(n_946), .ZN(n_945));
   NAND2_X1 i_577 (.A1(n_524), .A2(n_499), .ZN(n_946));
   NOR2_X1 i_578 (.A1(n_524), .A2(n_499), .ZN(n_954));
   NAND2_X1 i_579 (.A1(n_963), .A2(n_960), .ZN(n_957));
   INV_X1 i_580 (.A(p_2[35]), .ZN(n_960));
   INV_X1 i_581 (.A(p_1[34]), .ZN(n_962));
   INV_X1 i_582 (.A(p_1[35]), .ZN(n_963));
   FA_X1 i_583 (.A(p_10[36]), .B(p_11[36]), .CI(p_12[36]), .CO(n_964), .S(n_530));
   FA_X1 i_584 (.A(p_7[36]), .B(p_8[36]), .CI(p_9[36]), .CO(n_965), .S(n_528));
   FA_X1 i_585 (.A(p_4[36]), .B(p_5[36]), .CI(p_6[36]), .CO(n_966), .S(n_526));
   FA_X1 i_586 (.A(n_530), .B(n_528), .CI(n_526), .CO(n_967), .S(n_538));
   FA_X1 i_587 (.A(n_924), .B(n_925), .CI(n_919), .CO(n_968), .S(n_534));
   FA_X1 i_588 (.A(n_895), .B(n_929), .CI(n_534), .CO(n_969), .S(n_540));
   FA_X1 i_589 (.A(n_934), .B(n_538), .CI(n_540), .CO(n_970), .S(n_544));
   FA_X1 i_590 (.A(p_13[36]), .B(p_14[36]), .CI(n_923), .CO(n_971), .S(n_532));
   FA_X1 i_591 (.A(n_957), .B(n_933), .CI(n_532), .CO(n_972), .S(n_536));
   FA_X1 i_592 (.A(n_928), .B(n_920), .CI(n_536), .CO(n_973), .S(n_542));
   FA_X1 i_593 (.A(n_921), .B(n_542), .CI(n_935), .CO(n_974), .S(n_546));
   FA_X1 i_594 (.A(n_544), .B(n_546), .CI(n_936), .CO(n_975), .S(n_548));
   XNOR2_X1 i_595 (.A(p_1[36]), .B(n_976), .ZN(n_895));
   XOR2_X1 i_596 (.A(p_3[36]), .B(p_2[36]), .Z(n_976));
   XOR2_X1 i_597 (.A(n_980), .B(n_977), .Z(\aggregated_res[14] [36]));
   OAI21_X1 i_598 (.A(n_978), .B1(n_937), .B2(n_548), .ZN(n_977));
   NAND2_X1 i_599 (.A1(n_937), .A2(n_548), .ZN(n_978));
   NOR2_X1 i_600 (.A1(n_937), .A2(n_548), .ZN(n_979));
   OAI21_X1 i_601 (.A(n_1001), .B1(n_945), .B2(n_981), .ZN(n_980));
   OAI21_X1 i_602 (.A(n_1000), .B1(n_983), .B2(n_982), .ZN(n_981));
   NOR2_X1 i_603 (.A1(n_938), .A2(n_896), .ZN(n_982));
   INV_X1 i_604 (.A(n_985), .ZN(n_983));
   OAI211_X1 i_605 (.A(n_908), .B(n_986), .C1(n_997), .C2(n_990), .ZN(n_985));
   OAI21_X1 i_606 (.A(n_987), .B1(n_894), .B2(n_833), .ZN(n_986));
   OAI21_X1 i_607 (.A(n_841), .B1(n_999), .B2(n_989), .ZN(n_987));
   AOI21_X1 i_608 (.A(n_803), .B1(n_693), .B2(n_663), .ZN(n_989));
   NOR2_X1 i_609 (.A1(n_723), .A2(n_993), .ZN(n_990));
   AND3_X1 i_610 (.A1(n_737), .A2(n_735), .A3(n_995), .ZN(n_993));
   OAI21_X1 i_611 (.A(n_639), .B1(n_617), .B2(n_996), .ZN(n_995));
   AND3_X1 i_612 (.A1(n_527), .A2(n_513), .A3(n_1397), .ZN(n_996));
   OAI221_X1 i_613 (.A(n_998), .B1(n_894), .B2(n_833), .C1(n_693), .C2(n_663), 
      .ZN(n_997));
   INV_X1 i_614 (.A(n_999), .ZN(n_998));
   OAI21_X1 i_615 (.A(n_844), .B1(n_711), .B2(n_793), .ZN(n_999));
   NAND2_X1 i_616 (.A1(n_938), .A2(n_896), .ZN(n_1000));
   INV_X1 i_617 (.A(n_954), .ZN(n_1001));
   FA_X1 i_618 (.A(p_13[37]), .B(p_14[37]), .CI(n_964), .CO(n_1004), .S(n_556));
   FA_X1 i_619 (.A(n_968), .B(n_971), .CI(n_556), .CO(n_1005), .S(n_560));
   FA_X1 i_620 (.A(n_972), .B(n_560), .CI(n_969), .CO(n_1006), .S(n_566));
   FA_X1 i_621 (.A(p_10[37]), .B(p_11[37]), .CI(p_12[37]), .CO(n_1008), .S(n_554));
   FA_X1 i_622 (.A(p_7[37]), .B(p_8[37]), .CI(p_9[37]), .CO(n_1009), .S(n_552));
   FA_X1 i_623 (.A(p_4[37]), .B(p_5[37]), .CI(p_6[37]), .CO(n_1010), .S(n_550));
   FA_X1 i_624 (.A(n_554), .B(n_552), .CI(n_550), .CO(n_1011), .S(n_562));
   FA_X1 i_625 (.A(n_965), .B(n_966), .CI(n_897), .CO(n_1012), .S(n_558));
   FA_X1 i_626 (.A(n_893), .B(n_558), .CI(n_967), .CO(n_1014), .S(n_564));
   FA_X1 i_627 (.A(n_562), .B(n_973), .CI(n_564), .CO(n_1015), .S(n_568));
   FA_X1 i_628 (.A(n_970), .B(n_566), .CI(n_568), .CO(n_1016), .S(n_570));
   HA_X1 i_629 (.A(n_974), .B(n_570), .CO(n_1018), .S(n_1017));
   AOI21_X1 i_630 (.A(n_1019), .B1(n_1025), .B2(p_1[36]), .ZN(n_897));
   AOI21_X1 i_631 (.A(p_3[36]), .B1(p_2[36]), .B2(n_21), .ZN(n_1019));
   OAI21_X1 i_632 (.A(n_1023), .B1(n_1027), .B2(n_1024), .ZN(n_893));
   XOR2_X1 i_633 (.A(n_1021), .B(n_1020), .Z(\aggregated_res[14] [37]));
   AOI21_X1 i_634 (.A(n_1022), .B1(n_1017), .B2(n_975), .ZN(n_1020));
   AOI21_X1 i_635 (.A(n_979), .B1(n_980), .B2(n_978), .ZN(n_1021));
   NOR2_X1 i_636 (.A1(n_1017), .A2(n_975), .ZN(n_1022));
   NAND2_X1 i_637 (.A1(n_1027), .A2(n_1024), .ZN(n_1023));
   INV_X1 i_638 (.A(p_3[37]), .ZN(n_1024));
   INV_X1 i_639 (.A(p_2[36]), .ZN(n_1025));
   INV_X1 i_640 (.A(p_2[37]), .ZN(n_1027));
   FA_X1 i_641 (.A(p_11[38]), .B(p_12[38]), .CI(p_13[38]), .CO(n_579), .S(n_578));
   FA_X1 i_642 (.A(p_8[38]), .B(p_9[38]), .CI(p_10[38]), .CO(n_577), .S(n_576));
   FA_X1 i_643 (.A(p_14[39]), .B(n_579), .CI(n_577), .CO(n_603), .S(n_602));
   FA_X1 i_644 (.A(p_12[40]), .B(p_13[40]), .CI(p_14[40]), .CO(n_623), .S(n_622));
   FA_X1 i_645 (.A(n_889), .B(n_603), .CI(n_622), .CO(n_627), .S(n_626));
   FA_X1 i_646 (.A(n_1010), .B(n_1023), .CI(n_1012), .CO(n_583), .S(n_582));
   FA_X1 i_647 (.A(p_5[38]), .B(p_6[38]), .CI(p_7[38]), .CO(n_575), .S(n_574));
   FA_X1 i_648 (.A(p_14[38]), .B(n_1008), .CI(n_1009), .CO(n_581), .S(n_580));
   FA_X1 i_649 (.A(n_575), .B(n_892), .CI(n_581), .CO(n_605), .S(n_604));
   FA_X1 i_650 (.A(n_888), .B(n_583), .CI(n_604), .CO(n_609), .S(n_608));
   FA_X1 i_651 (.A(p_9[40]), .B(p_10[40]), .CI(p_11[40]), .CO(n_621), .S(n_620));
   FA_X1 i_652 (.A(p_6[40]), .B(p_7[40]), .CI(p_8[40]), .CO(n_619), .S(n_618));
   FA_X1 i_653 (.A(n_620), .B(n_618), .CI(n_885), .CO(n_629), .S(n_628));
   FA_X1 i_654 (.A(n_626), .B(n_609), .CI(n_628), .CO(n_633), .S(n_632));
   FA_X1 i_655 (.A(n_1004), .B(n_578), .CI(n_576), .CO(n_585), .S(n_584));
   FA_X1 i_656 (.A(n_580), .B(n_1011), .CI(n_1005), .CO(n_589), .S(n_1028));
   FA_X1 i_657 (.A(n_602), .B(n_585), .CI(n_589), .CO(n_611), .S(n_610));
   FA_X1 i_658 (.A(p_11[39]), .B(p_12[39]), .CI(p_13[39]), .CO(n_601), .S(n_600));
   FA_X1 i_659 (.A(p_8[39]), .B(p_9[39]), .CI(p_10[39]), .CO(n_599), .S(n_598));
   FA_X1 i_660 (.A(p_5[39]), .B(p_6[39]), .CI(p_7[39]), .CO(n_597), .S(n_596));
   FA_X1 i_661 (.A(n_601), .B(n_599), .CI(n_597), .CO(n_625), .S(n_624));
   FA_X1 i_662 (.A(n_600), .B(n_598), .CI(n_596), .CO(n_607), .S(n_606));
   FA_X1 i_663 (.A(n_605), .B(n_624), .CI(n_607), .CO(n_631), .S(n_630));
   FA_X1 i_664 (.A(n_574), .B(n_890), .CI(n_582), .CO(n_587), .S(n_586));
   FA_X1 i_665 (.A(n_587), .B(n_606), .CI(n_608), .CO(n_613), .S(n_612));
   FA_X1 i_666 (.A(n_611), .B(n_630), .CI(n_613), .CO(n_635), .S(n_634));
   FA_X1 i_667 (.A(n_1014), .B(n_586), .CI(n_584), .CO(n_591), .S(n_1031));
   FA_X1 i_668 (.A(n_610), .B(n_591), .CI(n_612), .CO(n_615), .S(n_1032));
   FA_X1 i_669 (.A(n_632), .B(n_634), .CI(n_615), .CO(n_637), .S(n_1033));
   FA_X1 i_670 (.A(n_623), .B(n_621), .CI(n_619), .CO(n_1034), .S(n_644));
   FA_X1 i_671 (.A(n_644), .B(n_629), .CI(n_627), .CO(n_1035), .S(n_650));
   FA_X1 i_672 (.A(p_12[41]), .B(p_13[41]), .CI(p_14[41]), .CO(n_1036), .S(n_642));
   FA_X1 i_673 (.A(n_887), .B(n_625), .CI(n_642), .CO(n_1037), .S(n_646));
   FA_X1 i_675 (.A(p_9[41]), .B(p_10[41]), .CI(p_11[41]), .CO(n_1038), .S(n_640));
   FA_X1 i_676 (.A(p_6[41]), .B(p_7[41]), .CI(p_8[41]), .CO(n_1041), .S(n_638));
   FA_X1 i_677 (.A(n_640), .B(n_638), .CI(n_883), .CO(n_1042), .S(n_648));
   FA_X1 i_678 (.A(n_646), .B(n_631), .CI(n_648), .CO(n_1043), .S(n_652));
   FA_X1 i_679 (.A(n_650), .B(n_633), .CI(n_652), .CO(n_1045), .S(n_654));
   HA_X1 i_680 (.A(n_635), .B(n_654), .CO(n_1046), .S(n_656));
   OAI21_X1 i_681 (.A(n_1060), .B1(n_1064), .B2(n_1062), .ZN(n_883));
   NAND2_X1 i_682 (.A1(n_1052), .A2(n_1048), .ZN(n_887));
   NAND2_X1 i_683 (.A1(p_4[40]), .A2(n_1051), .ZN(n_1048));
   XNOR2_X1 i_684 (.A(p_4[38]), .B(n_1049), .ZN(n_890));
   OAI21_X1 i_686 (.A(n_1055), .B1(p_3[38]), .B2(n_1061), .ZN(n_1049));
   XNOR2_X1 i_687 (.A(p_4[40]), .B(n_1050), .ZN(n_885));
   NAND2_X1 i_688 (.A1(n_1052), .A2(n_1051), .ZN(n_1050));
   OR2_X1 i_689 (.A1(n_1066), .A2(p_5[40]), .ZN(n_1051));
   NAND2_X1 i_690 (.A1(n_1066), .A2(p_5[40]), .ZN(n_1052));
   INV_X1 i_691 (.A(n_1053), .ZN(n_892));
   OAI22_X1 i_692 (.A1(p_3[38]), .A2(n_1061), .B1(p_4[38]), .B2(n_1054), 
      .ZN(n_1053));
   INV_X1 i_693 (.A(n_1055), .ZN(n_1054));
   NAND2_X1 i_694 (.A1(p_3[38]), .A2(n_1061), .ZN(n_1055));
   OAI21_X1 i_695 (.A(n_889), .B1(n_1065), .B2(n_1063), .ZN(n_888));
   NAND2_X1 i_696 (.A1(n_1065), .A2(n_1063), .ZN(n_889));
   NAND2_X1 i_697 (.A1(n_1058), .A2(n_1057), .ZN(n_1056));
   NAND2_X1 i_698 (.A1(n_637), .A2(n_656), .ZN(n_1057));
   OR2_X1 i_699 (.A1(n_637), .A2(n_656), .ZN(n_1058));
   NAND2_X1 i_700 (.A1(n_1064), .A2(n_1062), .ZN(n_1060));
   INV_X1 i_701 (.A(p_2[38]), .ZN(n_1061));
   INV_X1 i_702 (.A(p_5[41]), .ZN(n_1062));
   INV_X1 i_703 (.A(p_4[39]), .ZN(n_1063));
   INV_X1 i_704 (.A(p_4[41]), .ZN(n_1064));
   INV_X1 i_705 (.A(p_3[39]), .ZN(n_1065));
   INV_X1 i_706 (.A(p_3[40]), .ZN(n_1066));
   FA_X1 i_707 (.A(n_1006), .B(n_1028), .CI(n_1015), .CO(n_593), .S(n_1068));
   HA_X1 i_708 (.A(n_593), .B(n_1032), .CO(n_1070), .S(n_1069));
   INV_X1 i_709 (.A(n_1077), .ZN(n_1075));
   NOR2_X1 i_710 (.A1(n_1070), .A2(n_1033), .ZN(n_1077));
   FA_X1 i_711 (.A(n_1031), .B(n_1068), .CI(n_1016), .CO(n_595), .S(n_1078));
   FA_X1 i_712 (.A(p_7[42]), .B(p_8[42]), .CI(p_9[42]), .CO(n_1079), .S(n_658));
   FA_X1 i_713 (.A(n_1038), .B(n_1041), .CI(n_1060), .CO(n_1082), .S(n_664));
   FA_X1 i_714 (.A(n_658), .B(n_880), .CI(n_664), .CO(n_1084), .S(n_668));
   FA_X1 i_715 (.A(p_13[42]), .B(p_14[42]), .CI(n_1036), .CO(n_1085), .S(n_662));
   FA_X1 i_716 (.A(p_10[42]), .B(p_11[42]), .CI(p_12[42]), .CO(n_1086), .S(n_660));
   FA_X1 i_717 (.A(n_1034), .B(n_662), .CI(n_660), .CO(n_1087), .S(n_666));
   FA_X1 i_718 (.A(n_1042), .B(n_1037), .CI(n_1035), .CO(n_1088), .S(n_670));
   FA_X1 i_719 (.A(n_668), .B(n_666), .CI(n_670), .CO(n_1089), .S(n_672));
   FA_X1 i_720 (.A(n_1043), .B(n_672), .CI(n_1045), .CO(n_1092), .S(n_674));
   XNOR2_X1 i_721 (.A(p_6[42]), .B(p_5[42]), .ZN(n_1093));
   XOR2_X1 i_722 (.A(n_1093), .B(p_4[42]), .Z(n_880));
   NOR2_X1 i_723 (.A1(n_1069), .A2(n_595), .ZN(n_1094));
   INV_X1 i_724 (.A(n_1094), .ZN(n_1095));
   NAND2_X1 i_725 (.A1(n_1069), .A2(n_595), .ZN(n_1096));
   INV_X1 i_726 (.A(n_1096), .ZN(n_1097));
   NAND3_X1 i_727 (.A1(n_1070), .A2(n_1033), .A3(n_1058), .ZN(n_1102));
   AOI21_X1 i_728 (.A(n_1097), .B1(n_1078), .B2(n_1018), .ZN(n_1103));
   NAND3_X1 i_729 (.A1(n_1095), .A2(n_1075), .A3(n_1058), .ZN(n_1104));
   OAI211_X1 i_730 (.A(n_1057), .B(n_1102), .C1(n_1103), .C2(n_1104), .ZN(n_1105));
   INV_X1 i_731 (.A(n_1105), .ZN(n_1106));
   NAND2_X1 i_732 (.A1(n_1017), .A2(n_975), .ZN(n_1108));
   AND2_X1 i_733 (.A1(n_946), .A2(n_1000), .ZN(n_1109));
   INV_X1 i_734 (.A(n_1001), .ZN(n_1112));
   OR3_X1 i_735 (.A1(n_1112), .A2(n_979), .A3(n_1022), .ZN(n_1115));
   OAI221_X1 i_736 (.A(n_1108), .B1(n_978), .B2(n_1022), .C1(n_1109), .C2(n_1115), 
      .ZN(n_1116));
   NOR4_X1 i_737 (.A1(n_1112), .A2(n_979), .A3(n_1022), .A4(n_982), .ZN(n_1119));
   INV_X1 i_738 (.A(n_1104), .ZN(n_1122));
   AOI21_X1 i_739 (.A(n_1116), .B1(n_985), .B2(n_1119), .ZN(n_1123));
   OAI21_X1 i_740 (.A(n_1122), .B1(n_1078), .B2(n_1018), .ZN(n_1128));
   OAI21_X1 i_741 (.A(n_1106), .B1(n_1123), .B2(n_1128), .ZN(n_1129));
   NOR2_X1 i_742 (.A1(n_1046), .A2(n_674), .ZN(n_1132));
   INV_X1 i_743 (.A(n_1132), .ZN(n_1133));
   NAND2_X1 i_744 (.A1(n_1046), .A2(n_674), .ZN(n_1134));
   NAND2_X1 i_745 (.A1(n_1133), .A2(n_1134), .ZN(n_1135));
   XNOR2_X1 i_746 (.A(n_1129), .B(n_1135), .ZN(\aggregated_res[14] [42]));
   INV_X1 i_747 (.A(n_1123), .ZN(n_1136));
   FA_X1 i_748 (.A(p_13[43]), .B(p_14[43]), .CI(n_1086), .CO(n_1138), .S(n_680));
   FA_X1 i_749 (.A(p_10[43]), .B(p_11[43]), .CI(p_12[43]), .CO(n_1139), .S(n_678));
   FA_X1 i_750 (.A(n_1085), .B(n_680), .CI(n_678), .CO(n_1140), .S(n_684));
   FA_X1 i_751 (.A(p_7[43]), .B(p_8[43]), .CI(p_9[43]), .CO(n_1141), .S(n_676));
   FA_X1 i_752 (.A(n_1079), .B(n_882), .CI(n_1082), .CO(n_1142), .S(n_682));
   FA_X1 i_753 (.A(n_676), .B(n_878), .CI(n_682), .CO(n_1143), .S(n_686));
   FA_X1 i_754 (.A(n_1087), .B(n_1084), .CI(n_686), .CO(n_1144), .S(n_688));
   FA_X1 i_755 (.A(n_684), .B(n_1088), .CI(n_688), .CO(n_1146), .S(n_690));
   HA_X1 i_756 (.A(n_1089), .B(n_690), .CO(n_1147), .S(n_692));
   AOI21_X1 i_757 (.A(n_17), .B1(p_4[42]), .B2(n_19), .ZN(n_882));
   OAI21_X1 i_758 (.A(n_1152), .B1(n_1155), .B2(n_1154), .ZN(n_878));
   XOR2_X1 i_759 (.A(n_1153), .B(n_1148), .Z(\aggregated_res[14] [43]));
   NAND2_X1 i_760 (.A1(n_1150), .A2(n_1149), .ZN(n_1148));
   NAND2_X1 i_761 (.A1(n_1092), .A2(n_692), .ZN(n_1149));
   INV_X1 i_762 (.A(n_1151), .ZN(n_1150));
   NOR2_X1 i_763 (.A1(n_1092), .A2(n_692), .ZN(n_1151));
   NAND2_X1 i_764 (.A1(n_1155), .A2(n_1154), .ZN(n_1152));
   AOI21_X1 i_765 (.A(n_1156), .B1(n_1129), .B2(n_1133), .ZN(n_1153));
   INV_X1 i_766 (.A(p_6[43]), .ZN(n_1154));
   INV_X1 i_767 (.A(p_5[43]), .ZN(n_1155));
   INV_X1 i_768 (.A(n_1134), .ZN(n_1156));
   FA_X1 i_769 (.A(p_8[44]), .B(p_9[44]), .CI(p_10[44]), .CO(n_695), .S(n_694));
   FA_X1 i_770 (.A(n_694), .B(n_875), .CI(n_1142), .CO(n_703), .S(n_702));
   FA_X1 i_771 (.A(p_14[44]), .B(n_1139), .CI(n_1141), .CO(n_699), .S(n_698));
   FA_X1 i_772 (.A(p_11[44]), .B(p_12[44]), .CI(p_13[44]), .CO(n_697), .S(n_696));
   FA_X1 i_773 (.A(n_1152), .B(n_1138), .CI(n_696), .CO(n_701), .S(n_700));
   FA_X1 i_774 (.A(n_698), .B(n_1140), .CI(n_700), .CO(n_705), .S(n_704));
   FA_X1 i_775 (.A(n_1143), .B(n_702), .CI(n_704), .CO(n_707), .S(n_706));
   FA_X1 i_776 (.A(n_1144), .B(n_706), .CI(n_1146), .CO(n_709), .S(n_708));
   FA_X1 i_777 (.A(p_8[45]), .B(p_9[45]), .CI(p_10[45]), .CO(n_1157), .S(n_710));
   FA_X1 i_778 (.A(p_14[45]), .B(n_697), .CI(n_695), .CO(n_1158), .S(n_714));
   FA_X1 i_779 (.A(n_710), .B(n_873), .CI(n_714), .CO(n_1159), .S(n_718));
   FA_X1 i_780 (.A(n_16), .B(n_699), .CI(n_1176), .CO(n_1161), .S(n_716));
   FA_X1 i_781 (.A(n_701), .B(n_703), .CI(n_716), .CO(n_1162), .S(n_720));
   FA_X1 i_782 (.A(n_718), .B(n_705), .CI(n_720), .CO(n_1163), .S(n_722));
   HA_X1 i_783 (.A(n_707), .B(n_722), .CO(n_1164), .S(n_724));
   OAI21_X1 i_784 (.A(n_1188), .B1(n_1197), .B2(n_1196), .ZN(n_873));
   XNOR2_X1 i_785 (.A(p_7[44]), .B(n_1165), .ZN(n_875));
   XOR2_X1 i_786 (.A(p_5[44]), .B(p_6[44]), .Z(n_1165));
   XNOR2_X1 i_787 (.A(n_1168), .B(n_1166), .ZN(\aggregated_res[14] [45]));
   NAND2_X1 i_788 (.A1(n_1173), .A2(n_1167), .ZN(n_1166));
   NAND2_X1 i_789 (.A1(n_1174), .A2(n_1169), .ZN(n_1167));
   NAND2_X1 i_790 (.A1(n_1171), .A2(n_1170), .ZN(n_1168));
   OR2_X1 i_791 (.A1(n_1147), .A2(n_708), .ZN(n_1169));
   NAND2_X1 i_792 (.A1(n_709), .A2(n_724), .ZN(n_1170));
   INV_X1 i_793 (.A(n_1172), .ZN(n_1171));
   NOR2_X1 i_794 (.A1(n_709), .A2(n_724), .ZN(n_1172));
   NAND2_X1 i_795 (.A1(n_1147), .A2(n_708), .ZN(n_1173));
   OAI21_X1 i_796 (.A(n_1149), .B1(n_1153), .B2(n_1151), .ZN(n_1174));
   INV_X1 i_797 (.A(p_7[44]), .ZN(n_1175));
   FA_X1 i_798 (.A(p_11[45]), .B(p_12[45]), .CI(p_13[45]), .CO(n_713), .S(n_1176));
   FA_X1 i_799 (.A(n_713), .B(n_1157), .CI(n_1188), .CO(n_1177), .S(n_730));
   FA_X1 i_800 (.A(n_870), .B(n_730), .CI(n_1161), .CO(n_1178), .S(n_734));
   FA_X1 i_801 (.A(p_12[46]), .B(p_13[46]), .CI(p_14[46]), .CO(n_1179), .S(n_728));
   FA_X1 i_802 (.A(p_9[46]), .B(p_10[46]), .CI(p_11[46]), .CO(n_1180), .S(n_726));
   FA_X1 i_803 (.A(n_1158), .B(n_728), .CI(n_726), .CO(n_1181), .S(n_732));
   FA_X1 i_804 (.A(n_1159), .B(n_732), .CI(n_1162), .CO(n_1182), .S(n_736));
   FA_X1 i_805 (.A(n_734), .B(n_1163), .CI(n_736), .CO(n_1184), .S(n_1183));
   XNOR2_X1 i_806 (.A(p_8[46]), .B(n_1185), .ZN(n_870));
   XOR2_X1 i_807 (.A(p_6[46]), .B(p_7[46]), .Z(n_1185));
   XNOR2_X1 i_808 (.A(n_1189), .B(n_1186), .ZN(\aggregated_res[14] [46]));
   OAI21_X1 i_809 (.A(n_1187), .B1(n_1183), .B2(n_1164), .ZN(n_1186));
   NAND2_X1 i_810 (.A1(n_1183), .A2(n_1164), .ZN(n_1187));
   NAND2_X1 i_811 (.A1(n_1197), .A2(n_1196), .ZN(n_1188));
   OAI21_X1 i_812 (.A(n_1192), .B1(n_1199), .B2(n_1190), .ZN(n_1189));
   OR2_X1 i_813 (.A1(n_1132), .A2(n_1195), .ZN(n_1190));
   INV_X1 i_814 (.A(n_1192), .ZN(n_1191));
   NOR2_X1 i_815 (.A1(n_1194), .A2(n_1193), .ZN(n_1192));
   OAI21_X1 i_816 (.A(n_1170), .B1(n_1172), .B2(n_1173), .ZN(n_1193));
   AOI21_X1 i_817 (.A(n_1195), .B1(n_1149), .B2(n_1134), .ZN(n_1194));
   NAND3_X1 i_818 (.A1(n_1169), .A2(n_1150), .A3(n_1171), .ZN(n_1195));
   INV_X1 i_819 (.A(p_7[45]), .ZN(n_1196));
   INV_X1 i_820 (.A(p_6[45]), .ZN(n_1197));
   INV_X1 i_821 (.A(p_8[46]), .ZN(n_1198));
   INV_X1 i_822 (.A(n_1129), .ZN(n_1199));
   FA_X1 i_823 (.A(p_12[47]), .B(p_13[47]), .CI(p_14[47]), .CO(n_743), .S(n_742));
   FA_X1 i_824 (.A(p_13[48]), .B(p_14[48]), .CI(n_743), .CO(n_757), .S(n_756));
   FA_X1 i_825 (.A(p_10[48]), .B(p_11[48]), .CI(p_12[48]), .CO(n_755), .S(n_754));
   FA_X1 i_826 (.A(n_756), .B(n_754), .CI(n_865), .CO(n_761), .S(n_760));
   FA_X1 i_827 (.A(p_9[47]), .B(p_10[47]), .CI(p_11[47]), .CO(n_741), .S(n_740));
   FA_X1 i_828 (.A(n_1179), .B(n_1180), .CI(n_872), .CO(n_745), .S(n_744));
   FA_X1 i_829 (.A(n_741), .B(n_869), .CI(n_745), .CO(n_759), .S(n_758));
   FA_X1 i_830 (.A(n_1177), .B(n_742), .CI(n_740), .CO(n_747), .S(n_746));
   FA_X1 i_831 (.A(n_868), .B(n_744), .CI(n_1181), .CO(n_749), .S(n_748));
   FA_X1 i_832 (.A(n_758), .B(n_747), .CI(n_749), .CO(n_763), .S(n_762));
   FA_X1 i_833 (.A(n_1178), .B(n_746), .CI(n_748), .CO(n_751), .S(n_750));
   FA_X1 i_834 (.A(n_760), .B(n_762), .CI(n_751), .CO(n_1200), .S(n_764));
   FA_X1 i_835 (.A(p_13[49]), .B(p_14[49]), .CI(n_755), .CO(n_1201), .S(n_768));
   FA_X1 i_836 (.A(n_867), .B(n_757), .CI(n_768), .CO(n_1202), .S(n_770));
   FA_X1 i_837 (.A(p_10[49]), .B(p_11[49]), .CI(p_12[49]), .CO(n_1203), .S(n_766));
   FA_X1 i_838 (.A(n_766), .B(n_863), .CI(n_759), .CO(n_1204), .S(n_772));
   FA_X1 i_839 (.A(n_761), .B(n_770), .CI(n_772), .CO(n_1205), .S(n_774));
   HA_X1 i_840 (.A(n_763), .B(n_774), .CO(n_1207), .S(n_1206));
   HA_X1 i_841 (.A(n_1182), .B(n_750), .CO(n_753), .S(n_1208));
   OAI21_X1 i_842 (.A(n_1224), .B1(n_1231), .B2(n_1227), .ZN(n_863));
   NAND2_X1 i_843 (.A1(n_1212), .A2(n_1209), .ZN(n_867));
   NAND2_X1 i_844 (.A1(p_9[48]), .A2(n_1211), .ZN(n_1209));
   OAI21_X1 i_845 (.A(n_869), .B1(n_1229), .B2(n_1226), .ZN(n_868));
   OAI222_X1 i_846 (.A1(p_6[46]), .A2(n_1198), .B1(n_1228), .B2(p_6[46]), 
      .C1(n_1228), .C2(n_1198), .ZN(n_872));
   NAND2_X1 i_847 (.A1(n_1229), .A2(n_1226), .ZN(n_869));
   XNOR2_X1 i_848 (.A(p_9[48]), .B(n_1210), .ZN(n_865));
   NAND2_X1 i_849 (.A1(n_1212), .A2(n_1211), .ZN(n_1210));
   OR2_X1 i_850 (.A1(n_1230), .A2(p_8[48]), .ZN(n_1211));
   NAND2_X1 i_851 (.A1(n_1230), .A2(p_8[48]), .ZN(n_1212));
   XOR2_X1 i_852 (.A(n_1215), .B(n_1213), .Z(\aggregated_res[14] [49]));
   OR2_X1 i_853 (.A1(n_1221), .A2(n_1214), .ZN(n_1213));
   AOI211_X1 i_854 (.A(n_1220), .B(n_1216), .C1(n_1218), .C2(n_1217), .ZN(n_1214));
   AOI21_X1 i_855 (.A(n_1223), .B1(n_1200), .B2(n_1206), .ZN(n_1215));
   NOR2_X1 i_856 (.A1(n_764), .A2(n_753), .ZN(n_1216));
   OAI22_X1 i_857 (.A1(n_1225), .A2(n_1189), .B1(n_1164), .B2(n_1183), .ZN(
      n_1217));
   NOR2_X1 i_858 (.A1(n_1220), .A2(n_1219), .ZN(n_1218));
   AND2_X1 i_859 (.A1(n_1208), .A2(n_1184), .ZN(n_1219));
   NOR2_X1 i_860 (.A1(n_1208), .A2(n_1184), .ZN(n_1220));
   INV_X1 i_861 (.A(n_1222), .ZN(n_1221));
   NAND2_X1 i_862 (.A1(n_764), .A2(n_753), .ZN(n_1222));
   NOR2_X1 i_863 (.A1(n_1200), .A2(n_1206), .ZN(n_1223));
   NAND2_X1 i_864 (.A1(n_1231), .A2(n_1227), .ZN(n_1224));
   INV_X1 i_865 (.A(n_1187), .ZN(n_1225));
   INV_X1 i_866 (.A(p_8[47]), .ZN(n_1226));
   INV_X1 i_867 (.A(p_8[49]), .ZN(n_1227));
   INV_X1 i_868 (.A(p_7[46]), .ZN(n_1228));
   INV_X1 i_869 (.A(p_7[47]), .ZN(n_1229));
   INV_X1 i_870 (.A(p_7[48]), .ZN(n_1230));
   INV_X1 i_871 (.A(p_9[49]), .ZN(n_1231));
   FA_X1 i_872 (.A(p_11[50]), .B(p_12[50]), .CI(p_13[50]), .CO(n_1232), .S(n_778));
   FA_X1 i_873 (.A(n_1201), .B(n_778), .CI(n_860), .CO(n_1233), .S(n_782));
   FA_X1 i_874 (.A(p_14[50]), .B(n_1203), .CI(n_1224), .CO(n_1234), .S(n_780));
   FA_X1 i_875 (.A(n_780), .B(n_1202), .CI(n_1204), .CO(n_1236), .S(n_784));
   FA_X1 i_876 (.A(n_782), .B(n_784), .CI(n_1205), .CO(n_1239), .S(n_1237));
   XNOR2_X1 i_877 (.A(p_10[50]), .B(n_1240), .ZN(n_860));
   XOR2_X1 i_878 (.A(p_8[50]), .B(p_9[50]), .Z(n_1240));
   XNOR2_X1 i_879 (.A(n_1245), .B(n_1242), .ZN(\aggregated_res[14] [50]));
   OAI21_X1 i_880 (.A(n_1243), .B1(n_1237), .B2(n_1207), .ZN(n_1242));
   NAND2_X1 i_881 (.A1(n_1237), .A2(n_1207), .ZN(n_1243));
   INV_X1 i_882 (.A(n_1245), .ZN(n_1244));
   NAND4_X1 i_883 (.A1(n_1248), .A2(n_1246), .A3(n_1252), .A4(n_1253), .ZN(
      n_1245));
   OAI21_X1 i_884 (.A(n_1256), .B1(n_1191), .B2(n_1247), .ZN(n_1246));
   NOR2_X1 i_885 (.A1(n_1190), .A2(n_1106), .ZN(n_1247));
   AOI21_X1 i_886 (.A(n_1249), .B1(n_1206), .B2(n_1200), .ZN(n_1248));
   OAI21_X1 i_887 (.A(n_1251), .B1(n_1223), .B2(n_1222), .ZN(n_1249));
   OAI21_X1 i_888 (.A(n_1258), .B1(n_1225), .B2(n_1219), .ZN(n_1251));
   NAND2_X1 i_889 (.A1(n_1116), .A2(n_1254), .ZN(n_1252));
   NAND3_X1 i_890 (.A1(n_1119), .A2(n_985), .A3(n_1254), .ZN(n_1253));
   NOR4_X1 i_891 (.A1(n_1257), .A2(n_1255), .A3(n_1260), .A4(n_1190), .ZN(n_1254));
   NOR2_X1 i_892 (.A1(n_1018), .A2(n_1078), .ZN(n_1255));
   INV_X1 i_893 (.A(n_1257), .ZN(n_1256));
   OAI21_X1 i_894 (.A(n_1258), .B1(n_1164), .B2(n_1183), .ZN(n_1257));
   NOR3_X1 i_895 (.A1(n_1223), .A2(n_1220), .A3(n_1216), .ZN(n_1258));
   INV_X1 i_896 (.A(p_10[50]), .ZN(n_1259));
   INV_X1 i_897 (.A(n_1122), .ZN(n_1260));
   FA_X1 i_898 (.A(p_11[51]), .B(p_12[51]), .CI(p_13[51]), .CO(n_1261), .S(n_788));
   FA_X1 i_899 (.A(n_1234), .B(n_788), .CI(n_858), .CO(n_1262), .S(n_792));
   FA_X1 i_900 (.A(p_14[51]), .B(n_1232), .CI(n_862), .CO(n_1263), .S(n_790));
   FA_X1 i_901 (.A(n_790), .B(n_1233), .CI(n_1236), .CO(n_1264), .S(n_794));
   HA_X1 i_902 (.A(n_792), .B(n_794), .CO(n_1265), .S(n_796));
   OAI222_X1 i_903 (.A1(p_8[50]), .A2(n_1259), .B1(n_1276), .B2(p_8[50]), 
      .C1(n_1276), .C2(n_1259), .ZN(n_862));
   OAI21_X1 i_904 (.A(n_1270), .B1(n_1277), .B2(n_1275), .ZN(n_858));
   XNOR2_X1 i_905 (.A(n_1271), .B(n_1266), .ZN(\aggregated_res[14] [51]));
   NOR2_X1 i_906 (.A1(n_1269), .A2(n_1267), .ZN(n_1266));
   INV_X1 i_907 (.A(n_1268), .ZN(n_1267));
   NAND2_X1 i_908 (.A1(n_1239), .A2(n_796), .ZN(n_1268));
   NOR2_X1 i_909 (.A1(n_1239), .A2(n_796), .ZN(n_1269));
   NAND2_X1 i_910 (.A1(n_1277), .A2(n_1275), .ZN(n_1270));
   INV_X1 i_911 (.A(n_1272), .ZN(n_1271));
   AOI21_X1 i_912 (.A(n_1274), .B1(n_1244), .B2(n_1243), .ZN(n_1272));
   INV_X1 i_913 (.A(n_1274), .ZN(n_1273));
   NOR2_X1 i_914 (.A1(n_1237), .A2(n_1207), .ZN(n_1274));
   INV_X1 i_915 (.A(p_10[51]), .ZN(n_1275));
   INV_X1 i_916 (.A(p_9[50]), .ZN(n_1276));
   INV_X1 i_917 (.A(p_9[51]), .ZN(n_1277));
   FA_X1 i_918 (.A(p_12[52]), .B(p_13[52]), .CI(p_14[52]), .CO(n_1278), .S(n_798));
   FA_X1 i_919 (.A(n_1261), .B(n_1270), .CI(n_1263), .CO(n_1279), .S(n_800));
   FA_X1 i_920 (.A(n_798), .B(n_855), .CI(n_800), .CO(n_1280), .S(n_802));
   FA_X1 i_921 (.A(n_1262), .B(n_802), .CI(n_1264), .CO(n_1281), .S(n_804));
   XNOR2_X1 i_922 (.A(p_11[52]), .B(n_1282), .ZN(n_855));
   XOR2_X1 i_923 (.A(p_9[52]), .B(p_10[52]), .Z(n_1282));
   XNOR2_X1 i_924 (.A(n_1285), .B(n_1284), .ZN(\aggregated_res[14] [52]));
   AOI21_X1 i_925 (.A(n_1269), .B1(n_1271), .B2(n_1268), .ZN(n_1284));
   OAI21_X1 i_926 (.A(n_1287), .B1(n_1265), .B2(n_804), .ZN(n_1285));
   NOR2_X1 i_927 (.A1(n_1265), .A2(n_804), .ZN(n_1286));
   NAND2_X1 i_928 (.A1(n_1265), .A2(n_804), .ZN(n_1287));
   INV_X1 i_929 (.A(p_11[52]), .ZN(n_1288));
   FA_X1 i_930 (.A(p_12[53]), .B(p_13[53]), .CI(p_14[53]), .CO(n_1289), .S(n_806));
   FA_X1 i_931 (.A(n_1278), .B(n_857), .CI(n_806), .CO(n_1290), .S(n_808));
   FA_X1 i_932 (.A(n_853), .B(n_1279), .CI(n_808), .CO(n_1291), .S(n_810));
   HA_X1 i_933 (.A(n_1280), .B(n_810), .CO(n_1293), .S(n_1292));
   OAI222_X1 i_934 (.A1(p_9[52]), .A2(n_1288), .B1(n_1311), .B2(p_9[52]), 
      .C1(n_1311), .C2(n_1288), .ZN(n_857));
   OAI21_X1 i_935 (.A(n_1307), .B1(n_1312), .B2(n_1310), .ZN(n_853));
   AOI211_X1 i_936 (.A(n_1294), .B(n_1299), .C1(n_1304), .C2(n_1302), .ZN(
      \aggregated_res[14] [53]));
   OAI33_X1 i_937 (.A1(n_1301), .A2(n_1297), .A3(n_1305), .B1(n_1286), .B2(
      n_1304), .B3(n_1295), .ZN(n_1294));
   INV_X1 i_938 (.A(n_1296), .ZN(n_1295));
   OAI21_X1 i_939 (.A(n_1287), .B1(n_1269), .B2(n_1298), .ZN(n_1296));
   NAND3_X1 i_940 (.A1(n_1248), .A2(n_1287), .A3(n_1298), .ZN(n_1297));
   AND2_X1 i_941 (.A1(n_1268), .A2(n_1243), .ZN(n_1298));
   NOR3_X1 i_942 (.A1(n_1286), .A2(n_1269), .A3(n_1300), .ZN(n_1299));
   OAI211_X1 i_943 (.A(n_1305), .B(n_1273), .C1(n_1313), .C2(n_1301), .ZN(n_1300));
   NAND3_X1 i_944 (.A1(n_1246), .A2(n_1253), .A3(n_1252), .ZN(n_1301));
   OAI21_X1 i_945 (.A(n_1309), .B1(n_1308), .B2(n_1303), .ZN(n_1302));
   AOI21_X1 i_946 (.A(n_1269), .B1(n_1268), .B2(n_1274), .ZN(n_1303));
   INV_X1 i_947 (.A(n_1305), .ZN(n_1304));
   AOI21_X1 i_948 (.A(n_1306), .B1(n_1292), .B2(n_1281), .ZN(n_1305));
   NOR2_X1 i_949 (.A1(n_1292), .A2(n_1281), .ZN(n_1306));
   NAND2_X1 i_950 (.A1(n_1312), .A2(n_1310), .ZN(n_1307));
   INV_X1 i_951 (.A(n_1287), .ZN(n_1308));
   INV_X1 i_952 (.A(n_1286), .ZN(n_1309));
   INV_X1 i_953 (.A(p_11[53]), .ZN(n_1310));
   INV_X1 i_954 (.A(p_10[52]), .ZN(n_1311));
   INV_X1 i_955 (.A(p_10[53]), .ZN(n_1312));
   INV_X1 i_956 (.A(n_1248), .ZN(n_1313));
   FA_X1 i_957 (.A(p_13[55]), .B(p_14[55]), .CI(n_852), .CO(n_821), .S(n_820));
   FA_X1 i_958 (.A(p_14[56]), .B(n_849), .CI(n_821), .CO(n_827), .S(n_826));
   FA_X1 i_959 (.A(p_13[54]), .B(p_14[54]), .CI(n_1289), .CO(n_815), .S(n_1314));
   FA_X1 i_960 (.A(n_815), .B(n_820), .CI(n_848), .CO(n_823), .S(n_1316));
   FA_X1 i_961 (.A(n_845), .B(n_826), .CI(n_823), .CO(n_1318), .S(n_1317));
   FA_X1 i_962 (.A(p_14[57]), .B(n_847), .CI(n_843), .CO(n_1319), .S(n_830));
   HA_X1 i_963 (.A(n_827), .B(n_830), .CO(n_1321), .S(n_1320));
   OAI21_X1 i_964 (.A(n_1332), .B1(n_1343), .B2(n_1336), .ZN(n_843));
   NAND2_X1 i_965 (.A1(n_1326), .A2(n_1322), .ZN(n_847));
   NAND2_X1 i_966 (.A1(p_13[56]), .A2(n_1325), .ZN(n_1322));
   OAI21_X1 i_967 (.A(n_849), .B1(n_1337), .B2(n_1335), .ZN(n_848));
   OAI21_X1 i_968 (.A(n_1323), .B1(n_1334), .B2(p_10[54]), .ZN(n_852));
   OAI21_X1 i_969 (.A(p_11[54]), .B1(p_12[54]), .B2(n_1333), .ZN(n_1323));
   NAND2_X1 i_970 (.A1(n_1337), .A2(n_1335), .ZN(n_849));
   XNOR2_X1 i_971 (.A(p_13[56]), .B(n_1324), .ZN(n_845));
   NAND2_X1 i_972 (.A1(n_1326), .A2(n_1325), .ZN(n_1324));
   OR2_X1 i_973 (.A1(n_1338), .A2(p_12[56]), .ZN(n_1325));
   NAND2_X1 i_974 (.A1(n_1338), .A2(p_12[56]), .ZN(n_1326));
   INV_X1 i_975 (.A(n_1328), .ZN(n_1327));
   AOI21_X1 i_976 (.A(n_1330), .B1(n_1318), .B2(n_1320), .ZN(n_1328));
   NAND2_X1 i_977 (.A1(n_1318), .A2(n_1320), .ZN(n_1329));
   NOR2_X1 i_978 (.A1(n_1318), .A2(n_1320), .ZN(n_1330));
   NAND2_X1 i_979 (.A1(n_1343), .A2(n_1336), .ZN(n_1332));
   INV_X1 i_980 (.A(p_10[54]), .ZN(n_1333));
   INV_X1 i_981 (.A(p_12[54]), .ZN(n_1334));
   INV_X1 i_982 (.A(p_12[55]), .ZN(n_1335));
   INV_X1 i_983 (.A(p_12[57]), .ZN(n_1336));
   INV_X1 i_984 (.A(p_11[55]), .ZN(n_1337));
   INV_X1 i_985 (.A(p_11[56]), .ZN(n_1338));
   INV_X1 i_986 (.A(p_13[57]), .ZN(n_1343));
   FA_X1 i_987 (.A(n_1332), .B(n_840), .CI(n_1319), .CO(n_1344), .S(n_834));
   XNOR2_X1 i_988 (.A(p_14[58]), .B(n_1345), .ZN(n_840));
   XOR2_X1 i_989 (.A(p_12[58]), .B(p_13[58]), .Z(n_1345));
   AND2_X1 i_990 (.A1(n_1348), .A2(n_1347), .ZN(n_1346));
   NAND2_X1 i_991 (.A1(n_1321), .A2(n_834), .ZN(n_1347));
   OR2_X1 i_992 (.A1(n_1321), .A2(n_834), .ZN(n_1348));
   INV_X1 i_993 (.A(p_14[58]), .ZN(n_1349));
   HA_X1 i_994 (.A(n_842), .B(n_838), .CO(n_837), .S(n_1350));
   INV_X1 i_995 (.A(n_1351), .ZN(n_838));
   AOI21_X1 i_996 (.A(n_1360), .B1(p_13[59]), .B2(p_14[59]), .ZN(n_1351));
   OAI222_X1 i_997 (.A1(p_12[58]), .A2(n_1349), .B1(n_1364), .B2(p_12[58]), 
      .C1(n_1364), .C2(n_1349), .ZN(n_842));
   INV_X1 i_998 (.A(n_1353), .ZN(n_1352));
   NOR2_X1 i_999 (.A1(n_1355), .A2(n_1354), .ZN(n_1353));
   NOR2_X1 i_1000 (.A1(n_837), .A2(n_1356), .ZN(n_1354));
   AND2_X1 i_1001 (.A1(n_837), .A2(n_1356), .ZN(n_1355));
   XOR2_X1 i_1002 (.A(n_1360), .B(n_1357), .Z(n_1356));
   OAI21_X1 i_1003 (.A(n_1358), .B1(n_1366), .B2(p_14[60]), .ZN(n_1357));
   NAND2_X1 i_1004 (.A1(n_1366), .A2(p_14[60]), .ZN(n_1358));
   INV_X1 i_1005 (.A(n_1360), .ZN(n_1359));
   NOR2_X1 i_1006 (.A1(p_13[59]), .A2(p_14[59]), .ZN(n_1360));
   INV_X1 i_1007 (.A(p_13[58]), .ZN(n_1364));
   INV_X1 i_1008 (.A(p_13[60]), .ZN(n_1366));
   NOR2_X1 i_1009 (.A1(n_1355), .A2(n_1369), .ZN(n_1368));
   INV_X1 i_1010 (.A(n_1370), .ZN(n_1369));
   AOI21_X1 i_1011 (.A(n_1372), .B1(n_1344), .B2(n_1350), .ZN(n_1370));
   NAND2_X1 i_1012 (.A1(n_1344), .A2(n_1350), .ZN(n_1371));
   NOR2_X1 i_1013 (.A1(n_1344), .A2(n_1350), .ZN(n_1372));
   OAI21_X1 i_1014 (.A(n_1374), .B1(p_14[62]), .B2(n_1382), .ZN(n_1373));
   AOI211_X1 i_1015 (.A(n_1375), .B(n_1380), .C1(n_1355), .C2(n_1378), .ZN(
      n_1374));
   AOI21_X1 i_1016 (.A(n_1376), .B1(n_1347), .B2(n_1371), .ZN(n_1375));
   NAND2_X1 i_1017 (.A1(n_1378), .A2(n_1377), .ZN(n_1376));
   NOR2_X1 i_1018 (.A1(n_1372), .A2(n_1354), .ZN(n_1377));
   NAND2_X1 i_1019 (.A1(p_14[61]), .A2(n_1381), .ZN(n_1378));
   INV_X1 i_1020 (.A(n_1380), .ZN(n_1379));
   NOR2_X1 i_1021 (.A1(p_14[61]), .A2(n_1381), .ZN(n_1380));
   OAI22_X1 i_1022 (.A1(p_14[60]), .A2(n_1366), .B1(n_1383), .B2(n_1359), 
      .ZN(n_1381));
   INV_X1 i_1023 (.A(p_14[61]), .ZN(n_1382));
   INV_X1 i_1024 (.A(n_1358), .ZN(n_1383));
   FA_X1 i_1025 (.A(n_1307), .B(n_1314), .CI(n_850), .CO(n_817), .S(n_816));
   HA_X1 i_1026 (.A(n_817), .B(n_1316), .CO(n_825), .S(n_824));
   FA_X1 i_1027 (.A(n_1290), .B(n_1291), .CI(n_816), .CO(n_819), .S(n_1384));
   XOR2_X1 i_1028 (.A(n_1334), .B(n_1385), .Z(n_850));
   XOR2_X1 i_1029 (.A(p_10[54]), .B(p_11[54]), .Z(n_1385));
   INV_X1 i_1030 (.A(n_1387), .ZN(n_1386));
   OAI221_X1 i_1031 (.A(n_1329), .B1(n_1330), .B2(n_1396), .C1(n_1390), .C2(
      n_1388), .ZN(n_1387));
   AOI21_X1 i_1032 (.A(n_1394), .B1(n_1384), .B2(n_1293), .ZN(n_1388));
   INV_X1 i_1033 (.A(n_1390), .ZN(n_1389));
   OAI221_X1 i_1034 (.A(n_1392), .B1(n_1317), .B2(n_825), .C1(n_1318), .C2(
      n_1320), .ZN(n_1390));
   NOR2_X1 i_1035 (.A1(n_1317), .A2(n_825), .ZN(n_1391));
   INV_X1 i_1036 (.A(n_1393), .ZN(n_1392));
   NOR2_X1 i_1037 (.A1(n_824), .A2(n_819), .ZN(n_1393));
   INV_X1 i_1038 (.A(n_1395), .ZN(n_1394));
   NAND2_X1 i_1039 (.A1(n_824), .A2(n_819), .ZN(n_1395));
   NAND2_X1 i_1040 (.A1(n_1317), .A2(n_825), .ZN(n_1396));
   NAND4_X1 i_1041 (.A1(n_541), .A2(n_453), .A3(n_1399), .A4(n_533), .ZN(n_1397));
   AOI21_X1 i_1042 (.A(n_519), .B1(n_549), .B2(n_547), .ZN(n_1399));
   NAND2_X1 i_1043 (.A1(n_549), .A2(n_547), .ZN(n_1400));
endmodule

module datapath__0_68(\aggregated_res[14] , p_0);
   input [63:0]\aggregated_res[14] ;
   output [63:0]p_0;

   AOI21_X1 i_0 (.A(n_13), .B1(\aggregated_res[14] [1]), .B2(
      \aggregated_res[14] [0]), .ZN(p_0[1]));
   AOI21_X1 i_1 (.A(n_10), .B1(\aggregated_res[14] [2]), .B2(n_11), .ZN(p_0[2]));
   AOI21_X1 i_2 (.A(n_8), .B1(\aggregated_res[14] [3]), .B2(n_9), .ZN(p_0[3]));
   AOI21_X1 i_3 (.A(n_5), .B1(\aggregated_res[14] [4]), .B2(n_7), .ZN(p_0[4]));
   AOI21_X1 i_4 (.A(n_3), .B1(\aggregated_res[14] [5]), .B2(n_4), .ZN(p_0[5]));
   AOI21_X1 i_5 (.A(n_6), .B1(\aggregated_res[14] [6]), .B2(n_2), .ZN(p_0[6]));
   INV_X1 i_6 (.A(n_3), .ZN(n_2));
   NOR2_X1 i_7 (.A1(\aggregated_res[14] [5]), .A2(n_4), .ZN(n_3));
   INV_X1 i_8 (.A(n_5), .ZN(n_4));
   NOR2_X1 i_9 (.A1(\aggregated_res[14] [4]), .A2(n_7), .ZN(n_5));
   AOI21_X1 i_10 (.A(n_32), .B1(\aggregated_res[14] [8]), .B2(n_39), .ZN(p_0[8]));
   AOI21_X1 i_11 (.A(n_15), .B1(\aggregated_res[14] [9]), .B2(n_17), .ZN(p_0[9]));
   AOI21_X1 i_23 (.A(n_47), .B1(\aggregated_res[14] [12]), .B2(n_41), .ZN(
      p_0[12]));
   AOI21_X1 i_24 (.A(n_45), .B1(\aggregated_res[14] [13]), .B2(n_46), .ZN(
      p_0[13]));
   AOI21_X1 i_12 (.A(n_53), .B1(\aggregated_res[14] [15]), .B2(n_12), .ZN(
      p_0[15]));
   INV_X1 i_13 (.A(n_43), .ZN(n_12));
   AOI21_X1 i_14 (.A(n_66), .B1(\aggregated_res[14] [18]), .B2(n_58), .ZN(
      p_0[18]));
   AOI21_X1 i_36 (.A(n_63), .B1(\aggregated_res[14] [19]), .B2(n_65), .ZN(
      p_0[19]));
   AOI21_X1 i_39 (.A(n_72), .B1(\aggregated_res[14] [22]), .B2(n_68), .ZN(
      p_0[22]));
   AOI21_X1 i_15 (.A(n_93), .B1(\aggregated_res[14] [26]), .B2(n_77), .ZN(
      p_0[26]));
   AOI21_X1 i_45 (.A(n_87), .B1(\aggregated_res[14] [28]), .B2(n_81), .ZN(
      p_0[28]));
   AOI21_X1 i_16 (.A(n_89), .B1(\aggregated_res[14] [30]), .B2(n_86), .ZN(
      p_0[30]));
   AOI21_X1 i_49 (.A(n_23), .B1(\aggregated_res[14] [32]), .B2(n_92), .ZN(
      p_0[32]));
   AOI21_X1 i_50 (.A(n_21), .B1(\aggregated_res[14] [33]), .B2(n_22), .ZN(
      p_0[33]));
   AOI21_X1 i_51 (.A(n_19), .B1(\aggregated_res[14] [34]), .B2(n_20), .ZN(
      p_0[34]));
   AOI21_X1 i_17 (.A(n_31), .B1(\aggregated_res[14] [35]), .B2(n_18), .ZN(
      p_0[35]));
   INV_X1 i_18 (.A(n_19), .ZN(n_18));
   NOR2_X1 i_19 (.A1(\aggregated_res[14] [34]), .A2(n_20), .ZN(n_19));
   INV_X1 i_20 (.A(n_21), .ZN(n_20));
   NOR2_X1 i_21 (.A1(\aggregated_res[14] [33]), .A2(n_22), .ZN(n_21));
   INV_X1 i_22 (.A(n_23), .ZN(n_22));
   NOR2_X1 i_25 (.A1(\aggregated_res[14] [32]), .A2(n_92), .ZN(n_23));
   AOI21_X1 i_26 (.A(n_29), .B1(\aggregated_res[14] [36]), .B2(n_30), .ZN(
      p_0[36]));
   AOI21_X1 i_27 (.A(n_27), .B1(\aggregated_res[14] [37]), .B2(n_28), .ZN(
      p_0[37]));
   AOI21_X1 i_28 (.A(n_25), .B1(\aggregated_res[14] [38]), .B2(n_26), .ZN(
      p_0[38]));
   AOI21_X1 i_29 (.A(n_78), .B1(\aggregated_res[14] [39]), .B2(n_24), .ZN(
      p_0[39]));
   INV_X1 i_30 (.A(n_25), .ZN(n_24));
   NOR2_X1 i_31 (.A1(\aggregated_res[14] [38]), .A2(n_26), .ZN(n_25));
   INV_X1 i_32 (.A(n_27), .ZN(n_26));
   NOR2_X1 i_33 (.A1(\aggregated_res[14] [37]), .A2(n_28), .ZN(n_27));
   INV_X1 i_34 (.A(n_29), .ZN(n_28));
   NOR2_X1 i_35 (.A1(\aggregated_res[14] [36]), .A2(n_30), .ZN(n_29));
   INV_X1 i_37 (.A(n_31), .ZN(n_30));
   NOR2_X1 i_38 (.A1(n_92), .A2(n_80), .ZN(n_31));
   AOI21_X1 i_40 (.A(n_37), .B1(\aggregated_res[14] [40]), .B2(n_98), .ZN(
      p_0[40]));
   AOI21_X1 i_41 (.A(n_35), .B1(\aggregated_res[14] [41]), .B2(n_36), .ZN(
      p_0[41]));
   AOI21_X1 i_42 (.A(n_97), .B1(\aggregated_res[14] [42]), .B2(n_34), .ZN(
      p_0[42]));
   INV_X1 i_43 (.A(n_35), .ZN(n_34));
   NOR2_X1 i_44 (.A1(\aggregated_res[14] [41]), .A2(n_36), .ZN(n_35));
   INV_X1 i_46 (.A(n_37), .ZN(n_36));
   NOR2_X1 i_47 (.A1(\aggregated_res[14] [40]), .A2(n_98), .ZN(n_37));
   AOI21_X1 i_82 (.A(n_112), .B1(\aggregated_res[14] [45]), .B2(n_107), .ZN(
      p_0[45]));
   AOI21_X1 i_48 (.A(n_140), .B1(\aggregated_res[14] [52]), .B2(n_130), .ZN(
      p_0[52]));
   INV_X1 i_52 (.A(n_98), .ZN(n_78));
   INV_X1 i_53 (.A(n_128), .ZN(p_0[49]));
   INV_X1 i_54 (.A(n_167), .ZN(p_0[59]));
   INV_X1 i_55 (.A(n_83), .ZN(n_93));
   AOI21_X1 i_56 (.A(n_152), .B1(n_151), .B2(\aggregated_res[14] [62]), .ZN(
      p_0[62]));
   NAND4_X1 i_57 (.A1(n_115), .A2(n_180), .A3(n_146), .A4(n_177), .ZN(n_151));
   OAI21_X1 i_58 (.A(n_178), .B1(\aggregated_res[14] [63]), .B2(n_152), .ZN(
      p_0[63]));
   NOR2_X1 i_59 (.A1(n_176), .A2(n_153), .ZN(n_152));
   NAND2_X1 i_60 (.A1(n_181), .A2(n_180), .ZN(n_153));
   AOI21_X1 i_61 (.A(n_172), .B1(n_169), .B2(\aggregated_res[14] [60]), .ZN(
      p_0[60]));
   INV_X1 i_62 (.A(n_101), .ZN(n_80));
   AOI21_X1 i_63 (.A(n_0), .B1(\aggregated_res[14] [7]), .B2(n_1), .ZN(p_0[7]));
   NOR2_X1 i_64 (.A1(\aggregated_res[14] [7]), .A2(n_1), .ZN(n_0));
   INV_X1 i_65 (.A(n_6), .ZN(n_1));
   NOR4_X1 i_66 (.A1(\aggregated_res[14] [6]), .A2(\aggregated_res[14] [5]), 
      .A3(\aggregated_res[14] [4]), .A4(n_7), .ZN(n_6));
   INV_X1 i_67 (.A(n_8), .ZN(n_7));
   NOR2_X1 i_68 (.A1(\aggregated_res[14] [3]), .A2(n_9), .ZN(n_8));
   INV_X1 i_69 (.A(n_10), .ZN(n_9));
   NOR2_X1 i_70 (.A1(\aggregated_res[14] [2]), .A2(n_11), .ZN(n_10));
   INV_X1 i_71 (.A(n_13), .ZN(n_11));
   NOR2_X1 i_72 (.A1(\aggregated_res[14] [1]), .A2(\aggregated_res[14] [0]), 
      .ZN(n_13));
   AOI21_X1 i_73 (.A(n_14), .B1(\aggregated_res[14] [10]), .B2(n_16), .ZN(
      p_0[10]));
   NOR2_X1 i_74 (.A1(\aggregated_res[14] [10]), .A2(n_16), .ZN(n_14));
   INV_X1 i_75 (.A(n_16), .ZN(n_15));
   NAND2_X1 i_76 (.A1(n_0), .A2(n_33), .ZN(n_16));
   INV_X1 i_77 (.A(n_32), .ZN(n_17));
   NOR2_X1 i_78 (.A1(n_39), .A2(\aggregated_res[14] [8]), .ZN(n_32));
   NOR2_X1 i_79 (.A1(\aggregated_res[14] [9]), .A2(\aggregated_res[14] [8]), 
      .ZN(n_33));
   INV_X1 i_80 (.A(\aggregated_res[14] [10]), .ZN(n_38));
   INV_X1 i_81 (.A(n_0), .ZN(n_39));
   INV_X1 i_83 (.A(n_40), .ZN(p_0[11]));
   OAI21_X1 i_84 (.A(n_41), .B1(n_42), .B2(n_14), .ZN(n_40));
   NAND4_X1 i_85 (.A1(n_0), .A2(n_38), .A3(n_33), .A4(n_42), .ZN(n_41));
   INV_X1 i_86 (.A(\aggregated_res[14] [11]), .ZN(n_42));
   AOI21_X1 i_87 (.A(n_43), .B1(\aggregated_res[14] [14]), .B2(n_44), .ZN(
      p_0[14]));
   NOR2_X1 i_88 (.A1(\aggregated_res[14] [14]), .A2(n_44), .ZN(n_43));
   INV_X1 i_89 (.A(n_45), .ZN(n_44));
   NOR2_X1 i_90 (.A1(\aggregated_res[14] [13]), .A2(n_46), .ZN(n_45));
   INV_X1 i_91 (.A(n_47), .ZN(n_46));
   NOR2_X1 i_92 (.A1(\aggregated_res[14] [12]), .A2(n_41), .ZN(n_47));
   INV_X1 i_93 (.A(\aggregated_res[14] [12]), .ZN(n_48));
   INV_X1 i_94 (.A(\aggregated_res[14] [13]), .ZN(n_49));
   INV_X1 i_95 (.A(\aggregated_res[14] [14]), .ZN(n_50));
   AOI21_X1 i_96 (.A(n_51), .B1(\aggregated_res[14] [16]), .B2(n_52), .ZN(
      p_0[16]));
   NOR2_X1 i_97 (.A1(\aggregated_res[14] [16]), .A2(n_52), .ZN(n_51));
   INV_X1 i_98 (.A(n_53), .ZN(n_52));
   NOR2_X1 i_99 (.A1(n_41), .A2(n_54), .ZN(n_53));
   NAND4_X1 i_100 (.A1(n_55), .A2(n_50), .A3(n_49), .A4(n_48), .ZN(n_54));
   INV_X1 i_101 (.A(\aggregated_res[14] [15]), .ZN(n_55));
   INV_X1 i_102 (.A(\aggregated_res[14] [16]), .ZN(n_56));
   INV_X1 i_103 (.A(n_57), .ZN(p_0[17]));
   OAI21_X1 i_104 (.A(n_58), .B1(n_60), .B2(n_51), .ZN(n_57));
   NAND3_X1 i_105 (.A1(n_60), .A2(n_59), .A3(n_56), .ZN(n_58));
   NOR2_X1 i_106 (.A1(n_54), .A2(n_41), .ZN(n_59));
   INV_X1 i_107 (.A(\aggregated_res[14] [17]), .ZN(n_60));
   INV_X1 i_108 (.A(n_61), .ZN(p_0[20]));
   OAI21_X1 i_109 (.A(n_62), .B1(n_67), .B2(n_63), .ZN(n_61));
   NAND2_X1 i_110 (.A1(n_67), .A2(n_63), .ZN(n_62));
   NOR2_X1 i_111 (.A1(\aggregated_res[14] [19]), .A2(n_65), .ZN(n_63));
   NOR2_X1 i_112 (.A1(\aggregated_res[14] [20]), .A2(\aggregated_res[14] [19]), 
      .ZN(n_64));
   INV_X1 i_113 (.A(n_66), .ZN(n_65));
   NOR2_X1 i_114 (.A1(n_58), .A2(\aggregated_res[14] [18]), .ZN(n_66));
   INV_X1 i_115 (.A(\aggregated_res[14] [20]), .ZN(n_67));
   AOI22_X1 i_116 (.A1(n_64), .A2(n_69), .B1(\aggregated_res[14] [21]), .B2(n_62), 
      .ZN(p_0[21]));
   NAND2_X1 i_117 (.A1(n_64), .A2(n_69), .ZN(n_68));
   NOR3_X1 i_118 (.A1(n_58), .A2(\aggregated_res[14] [21]), .A3(
      \aggregated_res[14] [18]), .ZN(n_69));
   INV_X1 i_119 (.A(n_70), .ZN(p_0[23]));
   OAI21_X1 i_120 (.A(n_71), .B1(n_73), .B2(n_72), .ZN(n_70));
   NAND2_X1 i_121 (.A1(n_73), .A2(n_72), .ZN(n_71));
   NOR2_X1 i_122 (.A1(n_68), .A2(\aggregated_res[14] [22]), .ZN(n_72));
   INV_X1 i_123 (.A(\aggregated_res[14] [23]), .ZN(n_73));
   AOI21_X1 i_124 (.A(n_74), .B1(\aggregated_res[14] [24]), .B2(n_71), .ZN(
      p_0[24]));
   NOR4_X1 i_125 (.A1(n_68), .A2(\aggregated_res[14] [24]), .A3(n_75), .A4(
      \aggregated_res[14] [22]), .ZN(n_74));
   INV_X1 i_126 (.A(n_73), .ZN(n_75));
   INV_X1 i_127 (.A(n_76), .ZN(p_0[25]));
   OAI21_X1 i_128 (.A(n_77), .B1(n_79), .B2(n_74), .ZN(n_76));
   NAND2_X1 i_129 (.A1(n_79), .A2(n_74), .ZN(n_77));
   INV_X1 i_130 (.A(\aggregated_res[14] [25]), .ZN(n_79));
   AOI21_X1 i_131 (.A(n_82), .B1(\aggregated_res[14] [27]), .B2(n_83), .ZN(
      p_0[27]));
   INV_X1 i_132 (.A(n_82), .ZN(n_81));
   NOR2_X1 i_133 (.A1(\aggregated_res[14] [27]), .A2(n_83), .ZN(n_82));
   NAND3_X1 i_134 (.A1(n_74), .A2(n_79), .A3(n_84), .ZN(n_83));
   INV_X1 i_135 (.A(\aggregated_res[14] [26]), .ZN(n_84));
   INV_X1 i_136 (.A(n_85), .ZN(p_0[29]));
   OAI21_X1 i_137 (.A(n_86), .B1(n_88), .B2(n_87), .ZN(n_85));
   NAND2_X1 i_138 (.A1(n_88), .A2(n_87), .ZN(n_86));
   NOR2_X1 i_139 (.A1(n_81), .A2(\aggregated_res[14] [28]), .ZN(n_87));
   INV_X1 i_140 (.A(\aggregated_res[14] [29]), .ZN(n_88));
   INV_X1 i_141 (.A(n_90), .ZN(n_89));
   NAND3_X1 i_142 (.A1(n_82), .A2(n_88), .A3(n_91), .ZN(n_90));
   NOR2_X1 i_143 (.A1(\aggregated_res[14] [30]), .A2(\aggregated_res[14] [28]), 
      .ZN(n_91));
   AOI21_X1 i_144 (.A(n_94), .B1(n_90), .B2(\aggregated_res[14] [31]), .ZN(
      p_0[31]));
   INV_X1 i_145 (.A(n_94), .ZN(n_92));
   NOR2_X1 i_146 (.A1(n_90), .A2(\aggregated_res[14] [31]), .ZN(n_94));
   INV_X1 i_147 (.A(n_95), .ZN(p_0[43]));
   OAI21_X1 i_148 (.A(n_96), .B1(n_105), .B2(n_97), .ZN(n_95));
   NAND2_X1 i_149 (.A1(n_105), .A2(n_97), .ZN(n_96));
   NOR2_X1 i_150 (.A1(n_102), .A2(n_98), .ZN(n_97));
   NAND4_X1 i_151 (.A1(n_104), .A2(n_100), .A3(n_101), .A4(n_94), .ZN(n_98));
   AND4_X1 i_152 (.A1(n_104), .A2(n_100), .A3(n_101), .A4(n_105), .ZN(n_99));
   NOR3_X1 i_153 (.A1(\aggregated_res[14] [39]), .A2(\aggregated_res[14] [38]), 
      .A3(\aggregated_res[14] [37]), .ZN(n_100));
   NOR4_X1 i_154 (.A1(\aggregated_res[14] [35]), .A2(\aggregated_res[14] [33]), 
      .A3(\aggregated_res[14] [34]), .A4(\aggregated_res[14] [32]), .ZN(n_101));
   INV_X1 i_155 (.A(n_103), .ZN(n_102));
   NOR3_X1 i_156 (.A1(\aggregated_res[14] [42]), .A2(\aggregated_res[14] [40]), 
      .A3(\aggregated_res[14] [41]), .ZN(n_103));
   INV_X1 i_157 (.A(\aggregated_res[14] [36]), .ZN(n_104));
   INV_X1 i_158 (.A(\aggregated_res[14] [43]), .ZN(n_105));
   AOI21_X1 i_159 (.A(n_106), .B1(\aggregated_res[14] [44]), .B2(n_96), .ZN(
      p_0[44]));
   INV_X1 i_160 (.A(n_107), .ZN(n_106));
   NAND3_X1 i_161 (.A1(n_99), .A2(n_108), .A3(n_94), .ZN(n_107));
   AND2_X1 i_162 (.A1(n_109), .A2(n_103), .ZN(n_108));
   INV_X1 i_163 (.A(\aggregated_res[14] [44]), .ZN(n_109));
   INV_X1 i_164 (.A(n_110), .ZN(p_0[46]));
   OAI21_X1 i_165 (.A(n_111), .B1(n_113), .B2(n_112), .ZN(n_110));
   NAND2_X1 i_166 (.A1(n_113), .A2(n_112), .ZN(n_111));
   NOR2_X1 i_167 (.A1(\aggregated_res[14] [45]), .A2(n_107), .ZN(n_112));
   INV_X1 i_168 (.A(\aggregated_res[14] [46]), .ZN(n_113));
   AOI21_X1 i_169 (.A(n_115), .B1(\aggregated_res[14] [47]), .B2(n_111), 
      .ZN(p_0[47]));
   INV_X1 i_170 (.A(n_115), .ZN(n_114));
   NOR2_X1 i_171 (.A1(n_107), .A2(n_116), .ZN(n_115));
   NAND2_X1 i_172 (.A1(n_119), .A2(n_118), .ZN(n_116));
   INV_X1 i_173 (.A(n_118), .ZN(n_117));
   NOR2_X1 i_174 (.A1(\aggregated_res[14] [47]), .A2(\aggregated_res[14] [46]), 
      .ZN(n_118));
   INV_X1 i_175 (.A(\aggregated_res[14] [45]), .ZN(n_119));
   AOI22_X1 i_176 (.A1(n_121), .A2(n_115), .B1(\aggregated_res[14] [48]), 
      .B2(n_114), .ZN(p_0[48]));
   NAND2_X1 i_177 (.A1(n_121), .A2(n_115), .ZN(n_120));
   INV_X1 i_178 (.A(\aggregated_res[14] [48]), .ZN(n_121));
   OR4_X1 i_179 (.A1(\aggregated_res[14] [45]), .A2(\aggregated_res[14] [43]), 
      .A3(\aggregated_res[14] [39]), .A4(\aggregated_res[14] [38]), .ZN(n_122));
   NAND2_X1 i_180 (.A1(n_94), .A2(n_101), .ZN(n_123));
   NOR4_X1 i_181 (.A1(n_122), .A2(\aggregated_res[14] [37]), .A3(
      \aggregated_res[14] [36]), .A4(n_123), .ZN(n_124));
   NAND4_X1 i_182 (.A1(n_124), .A2(n_109), .A3(n_118), .A4(n_103), .ZN(n_125));
   OR3_X1 i_183 (.A1(n_125), .A2(\aggregated_res[14] [48]), .A3(
      \aggregated_res[14] [49]), .ZN(n_126));
   NAND2_X1 i_184 (.A1(n_120), .A2(\aggregated_res[14] [49]), .ZN(n_127));
   NAND2_X1 i_185 (.A1(n_126), .A2(n_127), .ZN(n_128));
   XOR2_X1 i_186 (.A(n_126), .B(\aggregated_res[14] [50]), .Z(p_0[50]));
   AND2_X1 i_187 (.A1(n_130), .A2(n_129), .ZN(p_0[51]));
   OAI21_X1 i_188 (.A(\aggregated_res[14] [51]), .B1(\aggregated_res[14] [50]), 
      .B2(n_126), .ZN(n_129));
   NAND2_X1 i_189 (.A1(n_115), .A2(n_131), .ZN(n_130));
   INV_X1 i_190 (.A(n_132), .ZN(n_131));
   NAND2_X1 i_191 (.A1(n_134), .A2(n_133), .ZN(n_132));
   NOR3_X1 i_192 (.A1(\aggregated_res[14] [51]), .A2(\aggregated_res[14] [48]), 
      .A3(\aggregated_res[14] [50]), .ZN(n_133));
   INV_X1 i_193 (.A(\aggregated_res[14] [49]), .ZN(n_134));
   NAND4_X1 i_194 (.A1(n_119), .A2(n_108), .A3(n_94), .A4(n_99), .ZN(n_135));
   INV_X1 i_195 (.A(n_131), .ZN(n_136));
   OR4_X1 i_196 (.A1(n_135), .A2(n_136), .A3(\aggregated_res[14] [52]), .A4(
      n_117), .ZN(n_137));
   XOR2_X1 i_197 (.A(n_137), .B(\aggregated_res[14] [53]), .Z(p_0[53]));
   NOR2_X1 i_198 (.A1(n_139), .A2(n_138), .ZN(p_0[54]));
   AOI21_X1 i_199 (.A(n_143), .B1(n_142), .B2(n_140), .ZN(n_138));
   NOR4_X1 i_200 (.A1(n_130), .A2(\aggregated_res[14] [52]), .A3(
      \aggregated_res[14] [53]), .A4(\aggregated_res[14] [54]), .ZN(n_139));
   INV_X1 i_201 (.A(n_137), .ZN(n_140));
   INV_X1 i_202 (.A(\aggregated_res[14] [52]), .ZN(n_141));
   INV_X1 i_203 (.A(\aggregated_res[14] [53]), .ZN(n_142));
   INV_X1 i_204 (.A(\aggregated_res[14] [54]), .ZN(n_143));
   INV_X1 i_205 (.A(n_144), .ZN(p_0[55]));
   OAI21_X1 i_206 (.A(n_145), .B1(n_149), .B2(n_139), .ZN(n_144));
   NAND3_X1 i_207 (.A1(n_150), .A2(n_106), .A3(n_146), .ZN(n_145));
   AND3_X1 i_208 (.A1(n_134), .A2(n_133), .A3(n_147), .ZN(n_146));
   INV_X1 i_209 (.A(n_148), .ZN(n_147));
   NAND4_X1 i_210 (.A1(n_149), .A2(n_142), .A3(n_143), .A4(n_141), .ZN(n_148));
   INV_X1 i_211 (.A(\aggregated_res[14] [55]), .ZN(n_149));
   INV_X1 i_212 (.A(n_116), .ZN(n_150));
   OAI22_X1 i_213 (.A1(n_155), .A2(\aggregated_res[14] [56]), .B1(n_145), 
      .B2(n_154), .ZN(p_0[56]));
   INV_X1 i_214 (.A(\aggregated_res[14] [56]), .ZN(n_154));
   INV_X1 i_215 (.A(n_145), .ZN(n_155));
   INV_X1 i_216 (.A(n_156), .ZN(p_0[57]));
   AOI21_X1 i_217 (.A(n_157), .B1(\aggregated_res[14] [57]), .B2(n_158), 
      .ZN(n_156));
   AOI21_X1 i_218 (.A(\aggregated_res[14] [57]), .B1(n_155), .B2(n_154), 
      .ZN(n_157));
   NOR2_X1 i_219 (.A1(\aggregated_res[14] [56]), .A2(n_145), .ZN(n_158));
   AOI22_X1 i_220 (.A1(n_164), .A2(n_162), .B1(\aggregated_res[14] [58]), 
      .B2(n_159), .ZN(p_0[58]));
   OR3_X1 i_221 (.A1(n_165), .A2(n_163), .A3(n_148), .ZN(n_159));
   NAND2_X1 i_222 (.A1(n_164), .A2(n_162), .ZN(n_160));
   INV_X1 i_223 (.A(n_162), .ZN(n_161));
   NOR2_X1 i_224 (.A1(\aggregated_res[14] [58]), .A2(n_163), .ZN(n_162));
   OR2_X1 i_225 (.A1(\aggregated_res[14] [57]), .A2(\aggregated_res[14] [56]), 
      .ZN(n_163));
   NOR2_X1 i_226 (.A1(n_166), .A2(n_165), .ZN(n_164));
   OR2_X1 i_227 (.A1(n_132), .A2(n_125), .ZN(n_165));
   INV_X1 i_228 (.A(n_147), .ZN(n_166));
   NAND2_X1 i_229 (.A1(n_169), .A2(n_168), .ZN(n_167));
   NAND2_X1 i_230 (.A1(n_160), .A2(\aggregated_res[14] [59]), .ZN(n_168));
   NAND2_X1 i_231 (.A1(n_155), .A2(n_171), .ZN(n_169));
   INV_X1 i_232 (.A(n_171), .ZN(n_170));
   NOR2_X1 i_233 (.A1(\aggregated_res[14] [59]), .A2(n_161), .ZN(n_171));
   INV_X1 i_234 (.A(n_173), .ZN(n_172));
   NAND3_X1 i_235 (.A1(n_164), .A2(n_162), .A3(n_174), .ZN(n_173));
   NOR2_X1 i_236 (.A1(\aggregated_res[14] [60]), .A2(\aggregated_res[14] [59]), 
      .ZN(n_174));
   AOI21_X1 i_237 (.A(n_175), .B1(\aggregated_res[14] [61]), .B2(n_173), 
      .ZN(p_0[61]));
   NOR2_X1 i_238 (.A1(\aggregated_res[14] [61]), .A2(n_176), .ZN(n_175));
   NAND4_X1 i_239 (.A1(n_106), .A2(n_150), .A3(n_146), .A4(n_177), .ZN(n_176));
   NOR2_X1 i_240 (.A1(n_170), .A2(\aggregated_res[14] [60]), .ZN(n_177));
   NAND4_X1 i_241 (.A1(n_180), .A2(n_155), .A3(n_177), .A4(n_179), .ZN(n_178));
   AND2_X1 i_242 (.A1(\aggregated_res[14] [63]), .A2(n_181), .ZN(n_179));
   INV_X1 i_243 (.A(\aggregated_res[14] [61]), .ZN(n_180));
   INV_X1 i_244 (.A(\aggregated_res[14] [62]), .ZN(n_181));
endmodule

module boothAlgoR4(Res, OVF, A, B, clk, reset, enable);
   output [63:0]Res;
   output OVF;
   input [31:0]A;
   input [31:0]B;
   input clk;
   input reset;
   input enable;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire [31:0]A_imm_2s_complement;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire [63:0]\aggregated_res[14] ;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire A_in;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire B_in;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_1_74;
   wire n_0_1_75;
   wire n_0_1_76;
   wire n_0_1_77;
   wire n_0_1_79;
   wire n_0_1_80;
   wire n_0_1_81;
   wire n_0_1_82;
   wire n_0_317;
   wire n_0_318;
   wire n_0_1_90;
   wire n_0_1_91;
   wire n_0_319;
   wire n_0_1_92;
   wire n_0_320;
   wire n_0_1_93;
   wire n_0_321;
   wire n_0_1_94;
   wire n_0_322;
   wire n_0_1_95;
   wire n_0_323;
   wire n_0_1_96;
   wire n_0_324;
   wire n_0_1_97;
   wire n_0_325;
   wire n_0_1_98;
   wire n_0_326;
   wire n_0_1_99;
   wire n_0_327;
   wire n_0_1_100;
   wire n_0_328;
   wire n_0_1_101;
   wire n_0_329;
   wire n_0_1_102;
   wire n_0_330;
   wire n_0_1_103;
   wire n_0_331;
   wire n_0_1_104;
   wire n_0_332;
   wire n_0_1_105;
   wire n_0_333;
   wire n_0_1_106;
   wire n_0_334;
   wire n_0_1_107;
   wire n_0_335;
   wire n_0_1_108;
   wire n_0_336;
   wire n_0_1_109;
   wire n_0_337;
   wire n_0_1_110;
   wire n_0_338;
   wire n_0_1_111;
   wire n_0_339;
   wire n_0_1_112;
   wire n_0_340;
   wire n_0_1_113;
   wire n_0_341;
   wire n_0_1_114;
   wire n_0_342;
   wire n_0_1_115;
   wire n_0_343;
   wire n_0_1_116;
   wire n_0_344;
   wire n_0_1_117;
   wire n_0_345;
   wire n_0_1_118;
   wire n_0_346;
   wire n_0_1_119;
   wire n_0_347;
   wire n_0_1_120;
   wire n_0_348;
   wire n_0_1_121;
   wire n_0_349;
   wire n_0_1_122;
   wire n_0_1_123;
   wire n_0_1_124;
   wire n_0_1_125;
   wire n_0_1_126;
   wire n_0_1_127;
   wire n_0_1_128;
   wire n_0_1_129;
   wire n_0_1_130;
   wire n_0_1_131;
   wire n_0_1_132;
   wire n_0_1_133;
   wire n_0_350;
   wire n_0_351;
   wire n_0_1_134;
   wire n_0_1_135;
   wire n_0_352;
   wire n_0_1_136;
   wire n_0_353;
   wire n_0_1_137;
   wire n_0_354;
   wire n_0_1_138;
   wire n_0_355;
   wire n_0_1_139;
   wire n_0_356;
   wire n_0_1_140;
   wire n_0_357;
   wire n_0_1_141;
   wire n_0_358;
   wire n_0_1_142;
   wire n_0_359;
   wire n_0_1_143;
   wire n_0_360;
   wire n_0_1_144;
   wire n_0_361;
   wire n_0_1_145;
   wire n_0_362;
   wire n_0_1_146;
   wire n_0_363;
   wire n_0_1_147;
   wire n_0_364;
   wire n_0_1_148;
   wire n_0_365;
   wire n_0_1_149;
   wire n_0_366;
   wire n_0_1_150;
   wire n_0_367;
   wire n_0_1_151;
   wire n_0_368;
   wire n_0_1_152;
   wire n_0_369;
   wire n_0_1_153;
   wire n_0_370;
   wire n_0_1_154;
   wire n_0_371;
   wire n_0_1_155;
   wire n_0_372;
   wire n_0_1_156;
   wire n_0_373;
   wire n_0_1_157;
   wire n_0_374;
   wire n_0_1_158;
   wire n_0_375;
   wire n_0_1_159;
   wire n_0_376;
   wire n_0_1_160;
   wire n_0_377;
   wire n_0_1_161;
   wire n_0_378;
   wire n_0_1_162;
   wire n_0_379;
   wire n_0_1_163;
   wire n_0_380;
   wire n_0_1_164;
   wire n_0_381;
   wire n_0_1_165;
   wire n_0_1_166;
   wire n_0_1_167;
   wire n_0_1_168;
   wire n_0_1_169;
   wire n_0_1_170;
   wire n_0_382;
   wire n_0_1_171;
   wire n_0_1_172;
   wire n_0_1_173;
   wire n_0_1_174;
   wire n_0_1_175;
   wire n_0_1_176;
   wire n_0_1_177;
   wire n_0_1_178;
   wire n_0_1_179;
   wire n_0_383;
   wire n_0_384;
   wire n_0_1_180;
   wire n_0_1_181;
   wire n_0_385;
   wire n_0_1_182;
   wire n_0_386;
   wire n_0_1_183;
   wire n_0_387;
   wire n_0_1_184;
   wire n_0_388;
   wire n_0_1_185;
   wire n_0_389;
   wire n_0_1_186;
   wire n_0_390;
   wire n_0_1_187;
   wire n_0_391;
   wire n_0_1_188;
   wire n_0_392;
   wire n_0_1_189;
   wire n_0_393;
   wire n_0_1_190;
   wire n_0_394;
   wire n_0_1_191;
   wire n_0_395;
   wire n_0_1_192;
   wire n_0_396;
   wire n_0_1_193;
   wire n_0_397;
   wire n_0_1_194;
   wire n_0_398;
   wire n_0_1_195;
   wire n_0_399;
   wire n_0_1_196;
   wire n_0_400;
   wire n_0_1_197;
   wire n_0_401;
   wire n_0_1_198;
   wire n_0_402;
   wire n_0_1_199;
   wire n_0_403;
   wire n_0_1_200;
   wire n_0_404;
   wire n_0_1_201;
   wire n_0_405;
   wire n_0_1_202;
   wire n_0_406;
   wire n_0_1_203;
   wire n_0_407;
   wire n_0_1_204;
   wire n_0_408;
   wire n_0_1_205;
   wire n_0_409;
   wire n_0_1_206;
   wire n_0_410;
   wire n_0_1_207;
   wire n_0_411;
   wire n_0_1_208;
   wire n_0_412;
   wire n_0_1_209;
   wire n_0_413;
   wire n_0_1_210;
   wire n_0_414;
   wire n_0_1_211;
   wire n_0_1_212;
   wire n_0_1_213;
   wire n_0_1_214;
   wire n_0_1_215;
   wire n_0_1_216;
   wire n_0_415;
   wire n_0_1_217;
   wire n_0_1_218;
   wire n_0_1_219;
   wire n_0_1_220;
   wire n_0_1_221;
   wire n_0_1_222;
   wire n_0_416;
   wire n_0_417;
   wire n_0_1_223;
   wire n_0_1_224;
   wire n_0_418;
   wire n_0_1_225;
   wire n_0_419;
   wire n_0_1_226;
   wire n_0_420;
   wire n_0_1_227;
   wire n_0_421;
   wire n_0_1_228;
   wire n_0_422;
   wire n_0_1_229;
   wire n_0_423;
   wire n_0_1_230;
   wire n_0_424;
   wire n_0_1_231;
   wire n_0_425;
   wire n_0_1_232;
   wire n_0_426;
   wire n_0_1_233;
   wire n_0_427;
   wire n_0_1_234;
   wire n_0_428;
   wire n_0_1_235;
   wire n_0_429;
   wire n_0_1_236;
   wire n_0_430;
   wire n_0_1_237;
   wire n_0_431;
   wire n_0_1_238;
   wire n_0_432;
   wire n_0_1_239;
   wire n_0_433;
   wire n_0_1_240;
   wire n_0_434;
   wire n_0_1_241;
   wire n_0_435;
   wire n_0_1_242;
   wire n_0_436;
   wire n_0_1_243;
   wire n_0_437;
   wire n_0_1_244;
   wire n_0_438;
   wire n_0_1_245;
   wire n_0_439;
   wire n_0_1_246;
   wire n_0_440;
   wire n_0_1_247;
   wire n_0_441;
   wire n_0_1_248;
   wire n_0_442;
   wire n_0_1_249;
   wire n_0_443;
   wire n_0_1_250;
   wire n_0_444;
   wire n_0_1_251;
   wire n_0_445;
   wire n_0_1_252;
   wire n_0_446;
   wire n_0_1_253;
   wire n_0_447;
   wire n_0_1_254;
   wire n_0_1_255;
   wire n_0_1_256;
   wire n_0_1_257;
   wire n_0_1_258;
   wire n_0_1_259;
   wire n_0_448;
   wire n_0_1_260;
   wire n_0_1_261;
   wire n_0_1_262;
   wire n_0_1_263;
   wire n_0_1_264;
   wire n_0_1_265;
   wire n_0_449;
   wire n_0_450;
   wire n_0_1_266;
   wire n_0_1_267;
   wire n_0_451;
   wire n_0_1_268;
   wire n_0_452;
   wire n_0_1_269;
   wire n_0_453;
   wire n_0_1_270;
   wire n_0_454;
   wire n_0_1_271;
   wire n_0_455;
   wire n_0_1_272;
   wire n_0_456;
   wire n_0_1_273;
   wire n_0_457;
   wire n_0_1_274;
   wire n_0_458;
   wire n_0_1_275;
   wire n_0_459;
   wire n_0_1_276;
   wire n_0_460;
   wire n_0_1_277;
   wire n_0_461;
   wire n_0_1_278;
   wire n_0_462;
   wire n_0_1_279;
   wire n_0_463;
   wire n_0_1_280;
   wire n_0_464;
   wire n_0_1_281;
   wire n_0_465;
   wire n_0_1_282;
   wire n_0_466;
   wire n_0_1_283;
   wire n_0_467;
   wire n_0_1_284;
   wire n_0_468;
   wire n_0_1_285;
   wire n_0_469;
   wire n_0_1_286;
   wire n_0_470;
   wire n_0_1_287;
   wire n_0_471;
   wire n_0_1_288;
   wire n_0_472;
   wire n_0_1_289;
   wire n_0_473;
   wire n_0_1_290;
   wire n_0_474;
   wire n_0_1_291;
   wire n_0_475;
   wire n_0_1_292;
   wire n_0_476;
   wire n_0_1_293;
   wire n_0_477;
   wire n_0_1_294;
   wire n_0_478;
   wire n_0_1_295;
   wire n_0_479;
   wire n_0_1_296;
   wire n_0_480;
   wire n_0_1_297;
   wire n_0_1_298;
   wire n_0_1_299;
   wire n_0_1_300;
   wire n_0_1_301;
   wire n_0_1_302;
   wire n_0_481;
   wire n_0_1_303;
   wire n_0_1_304;
   wire n_0_1_305;
   wire n_0_1_306;
   wire n_0_1_307;
   wire n_0_1_308;
   wire n_0_482;
   wire n_0_483;
   wire n_0_1_309;
   wire n_0_1_310;
   wire n_0_484;
   wire n_0_1_311;
   wire n_0_485;
   wire n_0_1_312;
   wire n_0_486;
   wire n_0_1_313;
   wire n_0_487;
   wire n_0_1_314;
   wire n_0_488;
   wire n_0_1_315;
   wire n_0_489;
   wire n_0_1_316;
   wire n_0_490;
   wire n_0_1_317;
   wire n_0_491;
   wire n_0_1_318;
   wire n_0_492;
   wire n_0_1_319;
   wire n_0_493;
   wire n_0_1_320;
   wire n_0_494;
   wire n_0_1_321;
   wire n_0_495;
   wire n_0_1_322;
   wire n_0_496;
   wire n_0_1_323;
   wire n_0_497;
   wire n_0_1_324;
   wire n_0_498;
   wire n_0_1_325;
   wire n_0_499;
   wire n_0_1_326;
   wire n_0_500;
   wire n_0_1_327;
   wire n_0_501;
   wire n_0_1_328;
   wire n_0_502;
   wire n_0_1_329;
   wire n_0_503;
   wire n_0_1_330;
   wire n_0_504;
   wire n_0_1_331;
   wire n_0_505;
   wire n_0_1_332;
   wire n_0_506;
   wire n_0_1_333;
   wire n_0_507;
   wire n_0_1_334;
   wire n_0_508;
   wire n_0_1_335;
   wire n_0_509;
   wire n_0_1_336;
   wire n_0_510;
   wire n_0_1_337;
   wire n_0_511;
   wire n_0_1_338;
   wire n_0_512;
   wire n_0_1_339;
   wire n_0_513;
   wire n_0_1_340;
   wire n_0_1_341;
   wire n_0_1_342;
   wire n_0_1_343;
   wire n_0_1_344;
   wire n_0_1_345;
   wire n_0_514;
   wire n_0_1_346;
   wire n_0_1_347;
   wire n_0_1_348;
   wire n_0_1_349;
   wire n_0_1_350;
   wire n_0_1_351;
   wire n_0_515;
   wire n_0_516;
   wire n_0_1_352;
   wire n_0_1_353;
   wire n_0_517;
   wire n_0_1_354;
   wire n_0_518;
   wire n_0_1_355;
   wire n_0_519;
   wire n_0_1_356;
   wire n_0_520;
   wire n_0_1_357;
   wire n_0_521;
   wire n_0_1_358;
   wire n_0_522;
   wire n_0_1_359;
   wire n_0_523;
   wire n_0_1_360;
   wire n_0_524;
   wire n_0_1_361;
   wire n_0_525;
   wire n_0_1_362;
   wire n_0_526;
   wire n_0_1_363;
   wire n_0_527;
   wire n_0_1_364;
   wire n_0_528;
   wire n_0_1_365;
   wire n_0_529;
   wire n_0_1_366;
   wire n_0_530;
   wire n_0_1_367;
   wire n_0_531;
   wire n_0_1_368;
   wire n_0_532;
   wire n_0_1_369;
   wire n_0_533;
   wire n_0_1_370;
   wire n_0_534;
   wire n_0_1_371;
   wire n_0_535;
   wire n_0_1_372;
   wire n_0_536;
   wire n_0_1_373;
   wire n_0_537;
   wire n_0_1_374;
   wire n_0_538;
   wire n_0_1_375;
   wire n_0_539;
   wire n_0_1_376;
   wire n_0_540;
   wire n_0_1_377;
   wire n_0_541;
   wire n_0_1_378;
   wire n_0_542;
   wire n_0_1_379;
   wire n_0_543;
   wire n_0_1_380;
   wire n_0_544;
   wire n_0_1_381;
   wire n_0_545;
   wire n_0_1_382;
   wire n_0_546;
   wire n_0_1_383;
   wire n_0_1_384;
   wire n_0_1_385;
   wire n_0_1_386;
   wire n_0_1_387;
   wire n_0_1_388;
   wire n_0_547;
   wire n_0_1_389;
   wire n_0_1_390;
   wire n_0_1_391;
   wire n_0_1_392;
   wire n_0_1_393;
   wire n_0_1_394;
   wire n_0_548;
   wire n_0_549;
   wire n_0_1_395;
   wire n_0_1_396;
   wire n_0_550;
   wire n_0_1_397;
   wire n_0_551;
   wire n_0_1_398;
   wire n_0_552;
   wire n_0_1_399;
   wire n_0_553;
   wire n_0_1_400;
   wire n_0_554;
   wire n_0_1_401;
   wire n_0_555;
   wire n_0_1_402;
   wire n_0_556;
   wire n_0_1_403;
   wire n_0_557;
   wire n_0_1_404;
   wire n_0_558;
   wire n_0_1_405;
   wire n_0_559;
   wire n_0_1_406;
   wire n_0_560;
   wire n_0_1_407;
   wire n_0_561;
   wire n_0_1_408;
   wire n_0_562;
   wire n_0_1_409;
   wire n_0_563;
   wire n_0_1_410;
   wire n_0_564;
   wire n_0_1_411;
   wire n_0_565;
   wire n_0_1_412;
   wire n_0_566;
   wire n_0_1_413;
   wire n_0_567;
   wire n_0_1_414;
   wire n_0_568;
   wire n_0_1_415;
   wire n_0_569;
   wire n_0_1_416;
   wire n_0_570;
   wire n_0_1_417;
   wire n_0_571;
   wire n_0_1_418;
   wire n_0_572;
   wire n_0_1_419;
   wire n_0_573;
   wire n_0_1_420;
   wire n_0_574;
   wire n_0_1_421;
   wire n_0_575;
   wire n_0_1_422;
   wire n_0_576;
   wire n_0_1_423;
   wire n_0_577;
   wire n_0_1_424;
   wire n_0_578;
   wire n_0_1_425;
   wire n_0_579;
   wire n_0_1_426;
   wire n_0_1_427;
   wire n_0_1_428;
   wire n_0_1_429;
   wire n_0_1_430;
   wire n_0_1_431;
   wire n_0_580;
   wire n_0_1_432;
   wire n_0_1_433;
   wire n_0_1_434;
   wire n_0_1_435;
   wire n_0_1_436;
   wire n_0_1_437;
   wire n_0_581;
   wire n_0_582;
   wire n_0_1_438;
   wire n_0_1_439;
   wire n_0_583;
   wire n_0_1_440;
   wire n_0_584;
   wire n_0_1_441;
   wire n_0_585;
   wire n_0_1_442;
   wire n_0_586;
   wire n_0_1_443;
   wire n_0_587;
   wire n_0_1_444;
   wire n_0_588;
   wire n_0_1_445;
   wire n_0_589;
   wire n_0_1_446;
   wire n_0_590;
   wire n_0_1_447;
   wire n_0_591;
   wire n_0_1_448;
   wire n_0_592;
   wire n_0_1_449;
   wire n_0_593;
   wire n_0_1_450;
   wire n_0_594;
   wire n_0_1_451;
   wire n_0_595;
   wire n_0_1_452;
   wire n_0_596;
   wire n_0_1_453;
   wire n_0_597;
   wire n_0_1_454;
   wire n_0_598;
   wire n_0_1_455;
   wire n_0_599;
   wire n_0_1_456;
   wire n_0_600;
   wire n_0_1_457;
   wire n_0_601;
   wire n_0_1_458;
   wire n_0_602;
   wire n_0_1_459;
   wire n_0_603;
   wire n_0_1_460;
   wire n_0_604;
   wire n_0_1_461;
   wire n_0_605;
   wire n_0_1_462;
   wire n_0_606;
   wire n_0_1_463;
   wire n_0_607;
   wire n_0_1_464;
   wire n_0_608;
   wire n_0_1_465;
   wire n_0_609;
   wire n_0_1_466;
   wire n_0_610;
   wire n_0_1_467;
   wire n_0_611;
   wire n_0_1_468;
   wire n_0_612;
   wire n_0_1_469;
   wire n_0_1_470;
   wire n_0_1_471;
   wire n_0_1_472;
   wire n_0_1_473;
   wire n_0_1_474;
   wire n_0_613;
   wire n_0_1_475;
   wire n_0_1_476;
   wire n_0_1_477;
   wire n_0_1_478;
   wire n_0_1_479;
   wire n_0_1_480;
   wire n_0_614;
   wire n_0_615;
   wire n_0_1_481;
   wire n_0_1_482;
   wire n_0_616;
   wire n_0_1_483;
   wire n_0_617;
   wire n_0_1_484;
   wire n_0_618;
   wire n_0_1_485;
   wire n_0_619;
   wire n_0_1_486;
   wire n_0_620;
   wire n_0_1_487;
   wire n_0_621;
   wire n_0_1_488;
   wire n_0_622;
   wire n_0_1_489;
   wire n_0_623;
   wire n_0_1_490;
   wire n_0_624;
   wire n_0_1_491;
   wire n_0_625;
   wire n_0_1_492;
   wire n_0_626;
   wire n_0_1_493;
   wire n_0_627;
   wire n_0_1_494;
   wire n_0_628;
   wire n_0_1_495;
   wire n_0_629;
   wire n_0_1_496;
   wire n_0_630;
   wire n_0_1_497;
   wire n_0_631;
   wire n_0_1_498;
   wire n_0_632;
   wire n_0_1_499;
   wire n_0_633;
   wire n_0_1_500;
   wire n_0_634;
   wire n_0_1_501;
   wire n_0_635;
   wire n_0_1_502;
   wire n_0_636;
   wire n_0_1_503;
   wire n_0_637;
   wire n_0_1_504;
   wire n_0_638;
   wire n_0_1_505;
   wire n_0_639;
   wire n_0_1_506;
   wire n_0_640;
   wire n_0_1_507;
   wire n_0_641;
   wire n_0_1_508;
   wire n_0_642;
   wire n_0_1_509;
   wire n_0_643;
   wire n_0_1_510;
   wire n_0_644;
   wire n_0_1_511;
   wire n_0_645;
   wire n_0_1_512;
   wire n_0_1_513;
   wire n_0_1_514;
   wire n_0_1_515;
   wire n_0_1_516;
   wire n_0_1_517;
   wire n_0_646;
   wire n_0_1_518;
   wire n_0_1_519;
   wire n_0_1_520;
   wire n_0_1_521;
   wire n_0_1_522;
   wire n_0_1_523;
   wire n_0_647;
   wire n_0_648;
   wire n_0_1_524;
   wire n_0_1_525;
   wire n_0_649;
   wire n_0_1_526;
   wire n_0_650;
   wire n_0_1_527;
   wire n_0_651;
   wire n_0_1_528;
   wire n_0_652;
   wire n_0_1_529;
   wire n_0_653;
   wire n_0_1_530;
   wire n_0_654;
   wire n_0_1_531;
   wire n_0_655;
   wire n_0_1_532;
   wire n_0_656;
   wire n_0_1_533;
   wire n_0_657;
   wire n_0_1_534;
   wire n_0_658;
   wire n_0_1_535;
   wire n_0_659;
   wire n_0_1_536;
   wire n_0_660;
   wire n_0_1_537;
   wire n_0_661;
   wire n_0_1_538;
   wire n_0_662;
   wire n_0_1_539;
   wire n_0_663;
   wire n_0_1_540;
   wire n_0_664;
   wire n_0_1_541;
   wire n_0_665;
   wire n_0_1_542;
   wire n_0_666;
   wire n_0_1_543;
   wire n_0_667;
   wire n_0_1_544;
   wire n_0_668;
   wire n_0_1_545;
   wire n_0_669;
   wire n_0_1_546;
   wire n_0_670;
   wire n_0_1_547;
   wire n_0_671;
   wire n_0_1_548;
   wire n_0_672;
   wire n_0_1_549;
   wire n_0_673;
   wire n_0_1_550;
   wire n_0_674;
   wire n_0_1_551;
   wire n_0_675;
   wire n_0_1_552;
   wire n_0_676;
   wire n_0_1_553;
   wire n_0_1_560;
   wire n_0_679;
   wire n_0_1_561;
   wire n_0_1_562;
   wire n_0_1_563;
   wire n_0_1_564;
   wire n_0_1_565;
   wire n_0_1_566;
   wire n_0_680;
   wire n_0_681;
   wire n_0_1_567;
   wire n_0_1_568;
   wire n_0_682;
   wire n_0_1_569;
   wire n_0_683;
   wire n_0_1_570;
   wire n_0_684;
   wire n_0_1_571;
   wire n_0_685;
   wire n_0_1_572;
   wire n_0_686;
   wire n_0_1_573;
   wire n_0_687;
   wire n_0_1_574;
   wire n_0_688;
   wire n_0_1_575;
   wire n_0_689;
   wire n_0_1_576;
   wire n_0_690;
   wire n_0_1_577;
   wire n_0_691;
   wire n_0_1_578;
   wire n_0_692;
   wire n_0_1_579;
   wire n_0_693;
   wire n_0_1_580;
   wire n_0_694;
   wire n_0_1_581;
   wire n_0_695;
   wire n_0_1_582;
   wire n_0_696;
   wire n_0_1_583;
   wire n_0_697;
   wire n_0_1_584;
   wire n_0_698;
   wire n_0_1_585;
   wire n_0_699;
   wire n_0_1_586;
   wire n_0_700;
   wire n_0_1_587;
   wire n_0_701;
   wire n_0_1_588;
   wire n_0_703;
   wire n_0_1_590;
   wire n_0_704;
   wire n_0_1_591;
   wire n_0_705;
   wire n_0_1_592;
   wire n_0_706;
   wire n_0_1_593;
   wire n_0_707;
   wire n_0_1_594;
   wire n_0_708;
   wire n_0_1_595;
   wire n_0_709;
   wire n_0_1_596;
   wire n_0_711;
   wire n_0_1_598;
   wire n_0_1_603;
   wire n_0_712;
   wire n_0_1_604;
   wire n_0_1_605;
   wire n_0_1_606;
   wire n_0_1_607;
   wire n_0_1_608;
   wire n_0_1_609;
   wire n_0_713;
   wire n_0_714;
   wire n_0_1_610;
   wire n_0_1_611;
   wire n_0_715;
   wire n_0_1_612;
   wire n_0_716;
   wire n_0_1_613;
   wire n_0_717;
   wire n_0_1_614;
   wire n_0_718;
   wire n_0_1_615;
   wire n_0_719;
   wire n_0_1_616;
   wire n_0_720;
   wire n_0_1_617;
   wire n_0_721;
   wire n_0_1_618;
   wire n_0_722;
   wire n_0_1_619;
   wire n_0_723;
   wire n_0_1_620;
   wire n_0_724;
   wire n_0_1_621;
   wire n_0_725;
   wire n_0_1_622;
   wire n_0_726;
   wire n_0_1_623;
   wire n_0_727;
   wire n_0_1_624;
   wire n_0_728;
   wire n_0_1_625;
   wire n_0_729;
   wire n_0_1_626;
   wire n_0_730;
   wire n_0_1_627;
   wire n_0_731;
   wire n_0_1_628;
   wire n_0_732;
   wire n_0_1_629;
   wire n_0_733;
   wire n_0_1_630;
   wire n_0_734;
   wire n_0_1_631;
   wire n_0_735;
   wire n_0_1_632;
   wire n_0_736;
   wire n_0_1_633;
   wire n_0_737;
   wire n_0_1_634;
   wire n_0_738;
   wire n_0_1_635;
   wire n_0_740;
   wire n_0_1_637;
   wire n_0_741;
   wire n_0_1_638;
   wire n_0_742;
   wire n_0_1_639;
   wire n_0_744;
   wire n_0_1_641;
   wire n_0_1_646;
   wire n_0_745;
   wire n_0_1_647;
   wire n_0_1_648;
   wire n_0_1_649;
   wire n_0_1_650;
   wire n_0_1_651;
   wire n_0_1_652;
   wire n_0_746;
   wire n_0_747;
   wire n_0_1_653;
   wire n_0_1_654;
   wire n_0_748;
   wire n_0_1_655;
   wire n_0_749;
   wire n_0_1_656;
   wire n_0_750;
   wire n_0_1_657;
   wire n_0_751;
   wire n_0_1_658;
   wire n_0_752;
   wire n_0_1_659;
   wire n_0_753;
   wire n_0_1_660;
   wire n_0_754;
   wire n_0_1_661;
   wire n_0_755;
   wire n_0_1_662;
   wire n_0_756;
   wire n_0_1_663;
   wire n_0_757;
   wire n_0_1_664;
   wire n_0_758;
   wire n_0_1_665;
   wire n_0_759;
   wire n_0_1_666;
   wire n_0_760;
   wire n_0_1_667;
   wire n_0_761;
   wire n_0_1_668;
   wire n_0_762;
   wire n_0_1_669;
   wire n_0_763;
   wire n_0_1_670;
   wire n_0_764;
   wire n_0_1_671;
   wire n_0_765;
   wire n_0_1_672;
   wire n_0_766;
   wire n_0_1_673;
   wire n_0_767;
   wire n_0_1_674;
   wire n_0_768;
   wire n_0_1_675;
   wire n_0_769;
   wire n_0_1_676;
   wire n_0_770;
   wire n_0_1_677;
   wire n_0_771;
   wire n_0_1_678;
   wire n_0_773;
   wire n_0_1_680;
   wire n_0_774;
   wire n_0_1_681;
   wire n_0_775;
   wire n_0_1_682;
   wire n_0_776;
   wire n_0_1_683;
   wire n_0_777;
   wire n_0_1_684;
   wire n_0_1_689;
   wire n_0_778;
   wire n_0_1_690;
   wire n_0_1_691;
   wire n_0_1_692;
   wire n_0_1_693;
   wire n_0_1_694;
   wire n_0_1_695;
   wire n_0_779;
   wire n_0_780;
   wire n_0_1_696;
   wire n_0_1_697;
   wire n_0_781;
   wire n_0_1_698;
   wire n_0_782;
   wire n_0_1_699;
   wire n_0_783;
   wire n_0_1_700;
   wire n_0_784;
   wire n_0_1_701;
   wire n_0_786;
   wire n_0_1_703;
   wire n_0_787;
   wire n_0_1_704;
   wire n_0_788;
   wire n_0_1_705;
   wire n_0_789;
   wire n_0_1_706;
   wire n_0_790;
   wire n_0_1_707;
   wire n_0_791;
   wire n_0_1_708;
   wire n_0_792;
   wire n_0_1_709;
   wire n_0_793;
   wire n_0_1_710;
   wire n_0_794;
   wire n_0_1_711;
   wire n_0_795;
   wire n_0_1_712;
   wire n_0_796;
   wire n_0_1_713;
   wire n_0_798;
   wire n_0_1_715;
   wire n_0_799;
   wire n_0_1_716;
   wire n_0_800;
   wire n_0_1_717;
   wire n_0_802;
   wire n_0_1_719;
   wire n_0_803;
   wire n_0_1_720;
   wire n_0_804;
   wire n_0_1_721;
   wire n_0_805;
   wire n_0_1_722;
   wire n_0_808;
   wire n_0_1_725;
   wire n_0_1_732;
   wire n_0_811;
   wire n_0_1_733;
   wire n_0_1_734;
   wire n_0_1_735;
   wire n_0_1_736;
   wire n_0_1_737;
   wire n_0_1_738;
   wire n_0_812;
   wire n_0_1_739;
   wire n_0_814;
   wire n_0_1_740;
   wire n_0_815;
   wire n_0_1_741;
   wire n_0_816;
   wire n_0_1_742;
   wire n_0_817;
   wire n_0_1_743;
   wire n_0_818;
   wire n_0_1_744;
   wire n_0_819;
   wire n_0_1_745;
   wire n_0_820;
   wire n_0_1_746;
   wire n_0_821;
   wire n_0_1_747;
   wire n_0_822;
   wire n_0_1_748;
   wire n_0_824;
   wire n_0_1_750;
   wire n_0_825;
   wire n_0_1_751;
   wire n_0_830;
   wire n_0_1_756;
   wire n_0_831;
   wire n_0_1_757;
   wire n_0_832;
   wire n_0_1_758;
   wire n_0_833;
   wire n_0_1_759;
   wire n_0_834;
   wire n_0_1_760;
   wire n_0_835;
   wire n_0_1_761;
   wire n_0_836;
   wire n_0_1_762;
   wire n_0_837;
   wire n_0_1_763;
   wire n_0_838;
   wire n_0_1_764;
   wire n_0_839;
   wire n_0_1_765;
   wire n_0_840;
   wire n_0_1_766;
   wire n_0_842;
   wire n_0_1_768;
   wire n_0_1_774;
   wire [31:0]A_imm;
   wire n_0_1_780;
   wire n_0_1_781;
   wire n_0_1_782;
   wire n_0_1_783;
   wire n_0_1_787;
   wire n_0_1_788;
   wire n_0_1_789;
   wire n_0_1_790;
   wire n_0_1_791;
   wire n_0_1_792;
   wire n_0_1_793;
   wire n_0_1_794;
   wire n_0_1_795;
   wire n_0_1_797;
   wire n_0_1_798;
   wire n_0_1_799;
   wire n_0_1_800;
   wire n_0_1_801;
   wire n_0_1_803;
   wire n_0_1_805;
   wire n_0_1_807;
   wire n_0_1_809;
   wire n_0_1_811;
   wire n_0_1_812;
   wire n_0_1_813;
   wire n_0_1_814;
   wire n_0_1_815;
   wire n_0_1_816;
   wire n_0_1_817;
   wire n_0_1_819;
   wire n_0_1_820;
   wire n_0_1_821;
   wire n_0_1_822;
   wire n_0_1_823;
   wire n_0_1_824;
   wire n_0_1_825;
   wire n_0_1_827;
   wire n_0_1_829;
   wire n_0_1_831;
   wire n_0_1_833;
   wire n_0_1_835;
   wire n_0_1_839;
   wire n_0_1_840;
   wire n_0_1_841;
   wire n_0_1_842;
   wire n_0_1_843;
   wire n_0_1_844;
   wire n_0_1_845;
   wire n_0_1_846;
   wire n_0_1_847;
   wire n_0_1_848;
   wire n_0_1_849;
   wire n_0_1_850;
   wire n_0_1_851;
   wire n_0_1_852;
   wire n_0_1_853;
   wire n_0_1_854;
   wire n_0_1_855;
   wire n_0_1_856;
   wire n_0_1_857;
   wire n_0_1_858;
   wire n_0_1_859;
   wire n_0_1_860;
   wire n_0_1_861;
   wire n_0_1_862;
   wire n_0_1_863;
   wire n_0_1_864;
   wire n_0_1_865;
   wire n_0_1_866;
   wire n_0_1_867;
   wire n_0_1_868;
   wire n_0_1_784;
   wire n_0_1_776;
   wire n_0_188;
   wire n_0_1_0;
   wire n_0_189;
   wire n_0_1_1;
   wire n_0_1_2;
   wire n_0_190;
   wire n_0_1_3;
   wire n_0_191;
   wire n_0_1_4;
   wire n_0_192;
   wire n_0_1_5;
   wire n_0_193;
   wire n_0_1_6;
   wire n_0_194;
   wire n_0_1_7;
   wire n_0_195;
   wire n_0_1_8;
   wire n_0_196;
   wire n_0_1_9;
   wire n_0_197;
   wire n_0_1_10;
   wire n_0_198;
   wire n_0_1_11;
   wire n_0_199;
   wire n_0_1_12;
   wire n_0_200;
   wire n_0_1_13;
   wire n_0_201;
   wire n_0_1_14;
   wire n_0_202;
   wire n_0_1_15;
   wire n_0_203;
   wire n_0_1_16;
   wire n_0_1_17;
   wire n_0_204;
   wire n_0_1_18;
   wire n_0_1_19;
   wire n_0_205;
   wire n_0_1_20;
   wire n_0_1_21;
   wire n_0_206;
   wire n_0_1_22;
   wire n_0_1_23;
   wire n_0_207;
   wire n_0_1_24;
   wire n_0_1_25;
   wire n_0_208;
   wire n_0_1_26;
   wire n_0_1_27;
   wire n_0_209;
   wire n_0_1_28;
   wire n_0_1_29;
   wire n_0_210;
   wire n_0_1_30;
   wire n_0_1_31;
   wire n_0_211;
   wire n_0_1_32;
   wire n_0_1_33;
   wire n_0_212;
   wire n_0_1_34;
   wire n_0_1_35;
   wire n_0_213;
   wire n_0_1_36;
   wire n_0_1_37;
   wire n_0_214;
   wire n_0_1_38;
   wire n_0_1_39;
   wire n_0_215;
   wire n_0_1_40;
   wire n_0_1_41;
   wire n_0_216;
   wire n_0_1_42;
   wire n_0_1_43;
   wire n_0_217;
   wire n_0_1_44;
   wire n_0_1_45;
   wire n_0_218;
   wire n_0_1_46;
   wire n_0_219;
   wire n_0_1_47;
   wire n_0_220;
   wire n_0_1_48;
   wire n_0_1_49;
   wire n_0_221;
   wire n_0_1_50;
   wire n_0_1_51;
   wire n_0_222;
   wire n_0_1_52;
   wire n_0_1_53;
   wire n_0_223;
   wire n_0_1_54;
   wire n_0_1_55;
   wire n_0_224;
   wire n_0_1_56;
   wire n_0_1_57;
   wire n_0_225;
   wire n_0_1_58;
   wire n_0_1_59;
   wire n_0_226;
   wire n_0_1_60;
   wire n_0_1_61;
   wire n_0_227;
   wire n_0_1_62;
   wire n_0_1_63;
   wire n_0_228;
   wire n_0_1_64;
   wire n_0_1_65;
   wire n_0_229;
   wire n_0_1_66;
   wire n_0_1_67;
   wire n_0_230;
   wire n_0_1_68;
   wire n_0_1_69;
   wire n_0_231;
   wire n_0_1_70;
   wire n_0_1_71;
   wire n_0_232;
   wire n_0_1_72;
   wire n_0_1_73;
   wire n_0_233;
   wire n_0_1_78;
   wire n_0_1_83;
   wire n_0_234;
   wire n_0_1_84;
   wire n_0_235;
   wire n_0_1_85;
   wire n_0_236;
   wire n_0_1_86;
   wire n_0_237;
   wire n_0_1_87;
   wire n_0_238;
   wire n_0_1_88;
   wire n_0_1_89;
   wire n_0_239;
   wire n_0_1_554;
   wire n_0_1_555;
   wire n_0_240;
   wire n_0_1_589;
   wire n_0_1_597;
   wire n_0_241;
   wire n_0_1_636;
   wire n_0_1_640;
   wire n_0_242;
   wire n_0_1_679;
   wire n_0_1_702;
   wire n_0_243;
   wire n_0_1_714;
   wire n_0_244;
   wire n_0_1_718;
   wire n_0_245;
   wire n_0_1_723;
   wire n_0_246;
   wire n_0_1_724;
   wire n_0_1_726;
   wire n_0_247;
   wire n_0_1_727;
   wire n_0_248;
   wire n_0_1_749;
   wire n_0_249;
   wire n_0_1_752;
   wire n_0_1_753;
   wire n_0_250;
   wire n_0_1_754;
   wire n_0_1_755;
   wire n_0_1_767;
   wire n_0_1_769;
   wire n_0_1_773;
   wire n_0_1_777;
   wire n_0_1_779;
   wire n_0_1_785;
   wire n_0_1_838;
   wire n_0_1_869;
   wire n_0_1_870;
   wire n_0_1_871;
   wire n_0_1_872;
   wire n_0_1_873;
   wire n_0_1_874;
   wire n_0_1_875;
   wire n_0_1_876;
   wire n_0_1_877;
   wire n_0_1_878;
   wire n_0_1_879;
   wire n_0_1_880;
   wire n_0_1_881;
   wire n_0_1_882;
   wire n_0_1_883;
   wire n_0_1_884;
   wire n_0_1_885;
   wire n_0_1_886;
   wire n_0_1_887;
   wire n_0_1_888;
   wire n_0_1_889;
   wire n_0_1_890;
   wire n_0_1_891;
   wire n_0_1_892;
   wire n_0_1_893;
   wire n_0_1_894;
   wire n_0_1_895;
   wire n_0_1_896;
   wire n_0_1_897;
   wire n_0_1_898;
   wire n_0_1_899;
   wire n_0_1_900;
   wire n_0_1_901;
   wire n_0_1_902;
   wire n_0_1_903;
   wire n_0_1_904;
   wire n_0_1_905;
   wire n_0_1_906;
   wire n_0_1_907;
   wire n_0_1_908;
   wire n_0_1_909;
   wire n_0_283;
   wire n_0_1_910;
   wire n_0_677;
   wire n_0_1_911;
   wire n_0_1_912;
   wire n_0_678;
   wire n_0_1_913;
   wire n_0_1_559;
   wire n_0_1_914;
   wire n_0_1_558;
   wire n_0_1_557;
   wire n_0_1_915;
   wire n_0_1_556;
   wire n_0_702;
   wire n_0_1_916;
   wire n_0_1_917;
   wire n_0_710;
   wire n_0_1_918;
   wire n_0_1_601;
   wire n_0_1_600;
   wire n_0_1_919;
   wire n_0_1_602;
   wire n_0_1_920;
   wire n_0_1_599;
   wire n_0_1_921;
   wire n_0_739;
   wire n_0_1_922;
   wire n_0_1_923;
   wire n_0_743;
   wire n_0_1_924;
   wire n_0_1_642;
   wire n_0_1_643;
   wire n_0_1_925;
   wire n_0_1_645;
   wire n_0_1_926;
   wire n_0_1_644;
   wire n_0_772;
   wire n_0_1_927;
   wire n_0_1_688;
   wire n_0_1_928;
   wire n_0_1_687;
   wire n_0_1_686;
   wire n_0_1_929;
   wire n_0_1_685;
   wire n_0_1_930;
   wire n_0_785;
   wire n_0_1_931;
   wire n_0_1_786;
   wire n_0_1_932;
   wire n_0_797;
   wire n_0_1_933;
   wire n_0_1_810;
   wire n_0_1_934;
   wire n_0_801;
   wire n_0_1_935;
   wire n_0_1_818;
   wire n_0_1_936;
   wire n_0_806;
   wire n_0_1_937;
   wire n_0_1_938;
   wire n_0_807;
   wire n_0_1_939;
   wire n_0_1_830;
   wire n_0_1_940;
   wire n_0_809;
   wire n_0_1_941;
   wire n_0_1_942;
   wire n_0_810;
   wire n_0_1_943;
   wire n_0_1_731;
   wire n_0_1_944;
   wire n_0_1_945;
   wire n_0_1_729;
   wire n_0_1_836;
   wire n_0_1_946;
   wire n_0_1_730;
   wire n_0_1_947;
   wire n_0_1_728;
   wire n_0_1_948;
   wire n_0_813;
   wire n_0_1_949;
   wire n_0_823;
   wire n_0_1_950;
   wire n_0_1_796;
   wire n_0_826;
   wire n_0_1_951;
   wire n_0_1_802;
   wire n_0_827;
   wire n_0_1_952;
   wire n_0_1_804;
   wire n_0_828;
   wire n_0_1_953;
   wire n_0_1_806;
   wire n_0_829;
   wire n_0_1_954;
   wire n_0_841;
   wire n_0_1_955;
   wire n_0_1_770;
   wire n_0_843;
   wire n_0_1_956;
   wire n_0_1_771;
   wire n_0_1_957;
   wire n_0_844;
   wire n_0_1_958;
   wire n_0_1_959;
   wire n_0_1_772;
   wire n_0_1_960;
   wire n_0_1_775;
   wire n_0_1_961;
   wire n_0_1_962;
   wire n_0_1_963;
   wire n_0_1_964;
   wire n_0_1_965;
   wire n_0_1_966;
   wire n_0_1_778;
   wire n_0_1_967;
   wire n_0_1_968;
   wire n_0_1_969;
   wire n_0_1_808;
   wire n_0_1_826;
   wire n_0_1_828;
   wire n_0_1_832;
   wire n_0_1_834;
   wire n_0_1_970;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_1_837;

   datapath i_0_0 (.A_in({A_in, n_0_125, n_0_126, n_0_127, n_0_128, n_0_129, 
      n_0_130, n_0_131, n_0_132, n_0_133, n_0_134, n_0_135, n_0_136, n_0_137, 
      n_0_138, n_0_139, n_0_140, n_0_141, n_0_142, n_0_143, n_0_144, n_0_145, 
      n_0_146, n_0_147, n_0_148, n_0_149, n_0_150, n_0_151, n_0_152, n_0_153, 
      n_0_154, n_0_155}), .p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, uc_0}));
   datapath__0_0 i_0_2 (.A_imm({A_imm[31], A_imm[30], A_imm[29], A_imm[28], 
      A_imm[27], A_imm[26], A_imm[25], A_imm[24], A_imm[23], A_imm[22], 
      A_imm[21], A_imm[20], A_imm[19], A_imm[18], A_imm[17], A_imm[16], 
      A_imm[15], A_imm[14], A_imm[13], A_imm[12], A_imm[11], A_imm[10], A_imm[9], 
      A_imm[8], A_imm[7], A_imm[6], A_imm[5], A_imm[4], A_imm[3], A_imm[2], 
      A_imm[1], n_0_155}), .A_imm_2s_complement({A_imm_2s_complement[31], 
      A_imm_2s_complement[30], A_imm_2s_complement[29], A_imm_2s_complement[28], 
      A_imm_2s_complement[27], A_imm_2s_complement[26], A_imm_2s_complement[25], 
      A_imm_2s_complement[24], A_imm_2s_complement[23], A_imm_2s_complement[22], 
      A_imm_2s_complement[21], A_imm_2s_complement[20], A_imm_2s_complement[19], 
      A_imm_2s_complement[18], A_imm_2s_complement[17], A_imm_2s_complement[16], 
      A_imm_2s_complement[15], A_imm_2s_complement[14], A_imm_2s_complement[13], 
      A_imm_2s_complement[12], A_imm_2s_complement[11], A_imm_2s_complement[10], 
      A_imm_2s_complement[9], A_imm_2s_complement[8], A_imm_2s_complement[7], 
      A_imm_2s_complement[6], A_imm_2s_complement[5], A_imm_2s_complement[4], 
      A_imm_2s_complement[3], A_imm_2s_complement[2], A_imm_2s_complement[1], 
      uc_1}));
   datapath__0_1 i_0_3 (.B_in({B_in, n_0_156, n_0_157, n_0_158, n_0_159, n_0_160, 
      n_0_161, n_0_162, n_0_163, n_0_164, n_0_165, n_0_166, n_0_167, n_0_168, 
      n_0_169, n_0_170, n_0_171, n_0_172, n_0_173, n_0_174, n_0_175, n_0_176, 
      n_0_177, n_0_178, n_0_179, n_0_180, n_0_181, n_0_182, n_0_183, n_0_184, 
      n_0_185, n_0_186}), .p_0({n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, 
      n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, 
      n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, 
      n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, uc_2}));
   datapath__0_67 i_0_5 (.p_0({uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, 
      uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, 
      uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, 
      uc_31, n_0_811, n_0_810, n_0_809, n_0_808, n_0_807, n_0_806, n_0_805, 
      n_0_804, n_0_803, n_0_802, n_0_801, n_0_800, n_0_799, n_0_798, n_0_797, 
      n_0_796, n_0_795, n_0_794, n_0_793, n_0_792, n_0_791, n_0_790, n_0_789, 
      n_0_788, n_0_787, n_0_786, n_0_785, n_0_784, n_0_783, n_0_782, n_0_781, 
      n_0_780, n_0_779, uc_32, uc_33}), .p_1({uc_34, uc_35, uc_36, uc_37, uc_38, 
      uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, 
      uc_49, uc_50, uc_51, uc_52, uc_53, uc_54, uc_55, uc_56, uc_57, uc_58, 
      uc_59, uc_60, n_0_778, n_0_777, n_0_776, n_0_775, n_0_774, n_0_773, 
      n_0_772, n_0_771, n_0_770, n_0_769, n_0_768, n_0_767, n_0_766, n_0_765, 
      n_0_764, n_0_763, n_0_762, n_0_761, n_0_760, n_0_759, n_0_758, n_0_757, 
      n_0_756, n_0_755, n_0_754, n_0_753, n_0_752, n_0_751, n_0_750, n_0_749, 
      n_0_748, n_0_747, n_0_746, uc_61, uc_62, uc_63, uc_64}), .p_2({uc_65, 
      uc_66, uc_67, uc_68, uc_69, uc_70, uc_71, uc_72, uc_73, uc_74, uc_75, 
      uc_76, uc_77, uc_78, uc_79, uc_80, uc_81, uc_82, uc_83, uc_84, uc_85, 
      uc_86, uc_87, uc_88, uc_89, n_0_745, n_0_744, n_0_743, n_0_742, n_0_741, 
      n_0_740, n_0_739, n_0_738, n_0_737, n_0_736, n_0_735, n_0_734, n_0_733, 
      n_0_732, n_0_731, n_0_730, n_0_729, n_0_728, n_0_727, n_0_726, n_0_725, 
      n_0_724, n_0_723, n_0_722, n_0_721, n_0_720, n_0_719, n_0_718, n_0_717, 
      n_0_716, n_0_715, n_0_714, n_0_713, uc_90, uc_91, uc_92, uc_93, uc_94, 
      uc_95}), .p_3({uc_96, uc_97, uc_98, uc_99, uc_100, uc_101, uc_102, uc_103, 
      uc_104, uc_105, uc_106, uc_107, uc_108, uc_109, uc_110, uc_111, uc_112, 
      uc_113, uc_114, uc_115, uc_116, uc_117, uc_118, n_0_712, n_0_711, n_0_710, 
      n_0_709, n_0_708, n_0_707, n_0_706, n_0_705, n_0_704, n_0_703, n_0_702, 
      n_0_701, n_0_700, n_0_699, n_0_698, n_0_697, n_0_696, n_0_695, n_0_694, 
      n_0_693, n_0_692, n_0_691, n_0_690, n_0_689, n_0_688, n_0_687, n_0_686, 
      n_0_685, n_0_684, n_0_683, n_0_682, n_0_681, n_0_680, uc_119, uc_120, 
      uc_121, uc_122, uc_123, uc_124, uc_125, uc_126}), .p_4({uc_127, uc_128, 
      uc_129, uc_130, uc_131, uc_132, uc_133, uc_134, uc_135, uc_136, uc_137, 
      uc_138, uc_139, uc_140, uc_141, uc_142, uc_143, uc_144, uc_145, uc_146, 
      uc_147, n_0_679, n_0_678, n_0_677, n_0_676, n_0_675, n_0_674, n_0_673, 
      n_0_672, n_0_671, n_0_670, n_0_669, n_0_668, n_0_667, n_0_666, n_0_665, 
      n_0_664, n_0_663, n_0_662, n_0_661, n_0_660, n_0_659, n_0_658, n_0_657, 
      n_0_656, n_0_655, n_0_654, n_0_653, n_0_652, n_0_651, n_0_650, n_0_649, 
      n_0_648, n_0_647, uc_148, uc_149, uc_150, uc_151, uc_152, uc_153, uc_154, 
      uc_155, uc_156, uc_157}), .p_5({uc_158, uc_159, uc_160, uc_161, uc_162, 
      uc_163, uc_164, uc_165, uc_166, uc_167, uc_168, uc_169, uc_170, uc_171, 
      uc_172, uc_173, uc_174, uc_175, uc_176, n_0_646, n_0_645, n_0_644, n_0_643, 
      n_0_642, n_0_641, n_0_640, n_0_639, n_0_638, n_0_637, n_0_636, n_0_635, 
      n_0_634, n_0_633, n_0_632, n_0_631, n_0_630, n_0_629, n_0_628, n_0_627, 
      n_0_626, n_0_625, n_0_624, n_0_623, n_0_622, n_0_621, n_0_620, n_0_619, 
      n_0_618, n_0_617, n_0_616, n_0_615, n_0_614, uc_177, uc_178, uc_179, 
      uc_180, uc_181, uc_182, uc_183, uc_184, uc_185, uc_186, uc_187, uc_188}), 
      .p_6({uc_189, uc_190, uc_191, uc_192, uc_193, uc_194, uc_195, uc_196, 
      uc_197, uc_198, uc_199, uc_200, uc_201, uc_202, uc_203, uc_204, uc_205, 
      n_0_613, n_0_612, n_0_611, n_0_610, n_0_609, n_0_608, n_0_607, n_0_606, 
      n_0_605, n_0_604, n_0_603, n_0_602, n_0_601, n_0_600, n_0_599, n_0_598, 
      n_0_597, n_0_596, n_0_595, n_0_594, n_0_593, n_0_592, n_0_591, n_0_590, 
      n_0_589, n_0_588, n_0_587, n_0_586, n_0_585, n_0_584, n_0_583, n_0_582, 
      n_0_581, uc_206, uc_207, uc_208, uc_209, uc_210, uc_211, uc_212, uc_213, 
      uc_214, uc_215, uc_216, uc_217, uc_218, uc_219}), .p_7({uc_220, uc_221, 
      uc_222, uc_223, uc_224, uc_225, uc_226, uc_227, uc_228, uc_229, uc_230, 
      uc_231, uc_232, uc_233, uc_234, n_0_580, n_0_579, n_0_578, n_0_577, 
      n_0_576, n_0_575, n_0_574, n_0_573, n_0_572, n_0_571, n_0_570, n_0_569, 
      n_0_568, n_0_567, n_0_566, n_0_565, n_0_564, n_0_563, n_0_562, n_0_561, 
      n_0_560, n_0_559, n_0_558, n_0_557, n_0_556, n_0_555, n_0_554, n_0_553, 
      n_0_552, n_0_551, n_0_550, n_0_549, n_0_548, uc_235, uc_236, uc_237, 
      uc_238, uc_239, uc_240, uc_241, uc_242, uc_243, uc_244, uc_245, uc_246, 
      uc_247, uc_248, uc_249, uc_250}), .p_8({uc_251, uc_252, uc_253, uc_254, 
      uc_255, uc_256, uc_257, uc_258, uc_259, uc_260, uc_261, uc_262, uc_263, 
      n_0_547, n_0_546, n_0_545, n_0_544, n_0_543, n_0_542, n_0_541, n_0_540, 
      n_0_539, n_0_538, n_0_537, n_0_536, n_0_535, n_0_534, n_0_533, n_0_532, 
      n_0_531, n_0_530, n_0_529, n_0_528, n_0_527, n_0_526, n_0_525, n_0_524, 
      n_0_523, n_0_522, n_0_521, n_0_520, n_0_519, n_0_518, n_0_517, n_0_516, 
      n_0_515, uc_264, uc_265, uc_266, uc_267, uc_268, uc_269, uc_270, uc_271, 
      uc_272, uc_273, uc_274, uc_275, uc_276, uc_277, uc_278, uc_279, uc_280, 
      uc_281}), .p_9({uc_282, uc_283, uc_284, uc_285, uc_286, uc_287, uc_288, 
      uc_289, uc_290, uc_291, uc_292, n_0_514, n_0_513, n_0_512, n_0_511, 
      n_0_510, n_0_509, n_0_508, n_0_507, n_0_506, n_0_505, n_0_504, n_0_503, 
      n_0_502, n_0_501, n_0_500, n_0_499, n_0_498, n_0_497, n_0_496, n_0_495, 
      n_0_494, n_0_493, n_0_492, n_0_491, n_0_490, n_0_489, n_0_488, n_0_487, 
      n_0_486, n_0_485, n_0_484, n_0_483, n_0_482, uc_293, uc_294, uc_295, 
      uc_296, uc_297, uc_298, uc_299, uc_300, uc_301, uc_302, uc_303, uc_304, 
      uc_305, uc_306, uc_307, uc_308, uc_309, uc_310, uc_311, uc_312}), .p_10({
      uc_313, uc_314, uc_315, uc_316, uc_317, uc_318, uc_319, uc_320, uc_321, 
      n_0_481, n_0_480, n_0_479, n_0_478, n_0_477, n_0_476, n_0_475, n_0_474, 
      n_0_473, n_0_472, n_0_471, n_0_470, n_0_469, n_0_468, n_0_467, n_0_466, 
      n_0_465, n_0_464, n_0_463, n_0_462, n_0_461, n_0_460, n_0_459, n_0_458, 
      n_0_457, n_0_456, n_0_455, n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, 
      n_0_449, uc_322, uc_323, uc_324, uc_325, uc_326, uc_327, uc_328, uc_329, 
      uc_330, uc_331, uc_332, uc_333, uc_334, uc_335, uc_336, uc_337, uc_338, 
      uc_339, uc_340, uc_341, uc_342, uc_343}), .p_11({uc_344, uc_345, uc_346, 
      uc_347, uc_348, uc_349, uc_350, n_0_448, n_0_447, n_0_446, n_0_445, 
      n_0_444, n_0_443, n_0_442, n_0_441, n_0_440, n_0_439, n_0_438, n_0_437, 
      n_0_436, n_0_435, n_0_434, n_0_433, n_0_432, n_0_431, n_0_430, n_0_429, 
      n_0_428, n_0_427, n_0_426, n_0_425, n_0_424, n_0_423, n_0_422, n_0_421, 
      n_0_420, n_0_419, n_0_418, n_0_417, n_0_416, uc_351, uc_352, uc_353, 
      uc_354, uc_355, uc_356, uc_357, uc_358, uc_359, uc_360, uc_361, uc_362, 
      uc_363, uc_364, uc_365, uc_366, uc_367, uc_368, uc_369, uc_370, uc_371, 
      uc_372, uc_373, uc_374}), .p_12({uc_375, uc_376, uc_377, uc_378, uc_379, 
      n_0_415, n_0_414, n_0_413, n_0_412, n_0_411, n_0_410, n_0_409, n_0_408, 
      n_0_407, n_0_406, n_0_405, n_0_404, n_0_403, n_0_402, n_0_401, n_0_400, 
      n_0_399, n_0_398, n_0_397, n_0_396, n_0_395, n_0_394, n_0_393, n_0_392, 
      n_0_391, n_0_390, n_0_389, n_0_388, n_0_387, n_0_386, n_0_385, n_0_384, 
      n_0_383, uc_380, uc_381, uc_382, uc_383, uc_384, uc_385, uc_386, uc_387, 
      uc_388, uc_389, uc_390, uc_391, uc_392, uc_393, uc_394, uc_395, uc_396, 
      uc_397, uc_398, uc_399, uc_400, uc_401, uc_402, uc_403, uc_404, uc_405}), 
      .p_13({uc_406, uc_407, uc_408, n_0_382, n_0_381, n_0_380, n_0_379, n_0_378, 
      n_0_377, n_0_376, n_0_375, n_0_374, n_0_373, n_0_372, n_0_371, n_0_370, 
      n_0_369, n_0_368, n_0_367, n_0_366, n_0_365, n_0_364, n_0_363, n_0_362, 
      n_0_361, n_0_360, n_0_359, n_0_358, n_0_357, n_0_356, n_0_355, n_0_354, 
      n_0_353, n_0_352, n_0_351, n_0_350, uc_409, uc_410, uc_411, uc_412, uc_413, 
      uc_414, uc_415, uc_416, uc_417, uc_418, uc_419, uc_420, uc_421, uc_422, 
      uc_423, uc_424, uc_425, uc_426, uc_427, uc_428, uc_429, uc_430, uc_431, 
      uc_432, uc_433, uc_434, uc_435, uc_436}), .p_14({uc_437, n_0_349, n_0_348, 
      n_0_347, n_0_346, n_0_345, n_0_344, n_0_343, n_0_342, n_0_341, n_0_340, 
      n_0_339, n_0_338, n_0_337, n_0_336, n_0_335, n_0_334, n_0_333, n_0_332, 
      n_0_331, n_0_330, n_0_329, n_0_328, n_0_327, n_0_326, n_0_325, n_0_324, 
      n_0_323, n_0_322, n_0_321, n_0_320, n_0_319, n_0_318, n_0_317, uc_438, 
      uc_439, uc_440, uc_441, uc_442, uc_443, uc_444, uc_445, uc_446, uc_447, 
      uc_448, uc_449, uc_450, uc_451, uc_452, uc_453, uc_454, uc_455, uc_456, 
      uc_457, uc_458, uc_459, uc_460, uc_461, uc_462, uc_463, uc_464, uc_465, 
      uc_466, uc_467}), .p_15({uc_468, uc_469, uc_470, uc_471, uc_472, uc_473, 
      uc_474, uc_475, uc_476, uc_477, uc_478, uc_479, uc_480, uc_481, uc_482, 
      uc_483, uc_484, uc_485, uc_486, uc_487, uc_488, uc_489, uc_490, uc_491, 
      uc_492, uc_493, uc_494, uc_495, uc_496, uc_497, uc_498, n_0_844, n_0_843, 
      n_0_842, n_0_841, n_0_840, n_0_839, n_0_838, n_0_837, n_0_836, n_0_835, 
      n_0_834, n_0_833, n_0_832, n_0_831, n_0_830, n_0_829, n_0_828, n_0_827, 
      n_0_826, n_0_825, n_0_824, n_0_823, n_0_822, n_0_821, n_0_820, n_0_819, 
      n_0_818, n_0_817, n_0_816, n_0_815, n_0_814, uc_499, uc_500}), 
      .\aggregated_res[14] ({\aggregated_res[14] [63], \aggregated_res[14] [62], 
      \aggregated_res[14] [61], \aggregated_res[14] [60], 
      \aggregated_res[14] [59], \aggregated_res[14] [58], 
      \aggregated_res[14] [57], \aggregated_res[14] [56], 
      \aggregated_res[14] [55], \aggregated_res[14] [54], 
      \aggregated_res[14] [53], \aggregated_res[14] [52], 
      \aggregated_res[14] [51], \aggregated_res[14] [50], 
      \aggregated_res[14] [49], \aggregated_res[14] [48], 
      \aggregated_res[14] [47], \aggregated_res[14] [46], 
      \aggregated_res[14] [45], \aggregated_res[14] [44], 
      \aggregated_res[14] [43], \aggregated_res[14] [42], 
      \aggregated_res[14] [41], \aggregated_res[14] [40], 
      \aggregated_res[14] [39], \aggregated_res[14] [38], 
      \aggregated_res[14] [37], \aggregated_res[14] [36], 
      \aggregated_res[14] [35], \aggregated_res[14] [34], 
      \aggregated_res[14] [33], \aggregated_res[14] [32], 
      \aggregated_res[14] [31], \aggregated_res[14] [30], 
      \aggregated_res[14] [29], \aggregated_res[14] [28], 
      \aggregated_res[14] [27], \aggregated_res[14] [26], 
      \aggregated_res[14] [25], \aggregated_res[14] [24], 
      \aggregated_res[14] [23], \aggregated_res[14] [22], 
      \aggregated_res[14] [21], \aggregated_res[14] [20], 
      \aggregated_res[14] [19], \aggregated_res[14] [18], 
      \aggregated_res[14] [17], \aggregated_res[14] [16], 
      \aggregated_res[14] [15], \aggregated_res[14] [14], 
      \aggregated_res[14] [13], \aggregated_res[14] [12], 
      \aggregated_res[14] [11], \aggregated_res[14] [10], 
      \aggregated_res[14] [9], \aggregated_res[14] [8], \aggregated_res[14] [7], 
      \aggregated_res[14] [6], \aggregated_res[14] [5], \aggregated_res[14] [4], 
      \aggregated_res[14] [3], \aggregated_res[14] [2], uc_501, uc_502}));
   datapath__0_68 i_0_6 (.\aggregated_res[14] ({\aggregated_res[14] [63], 
      \aggregated_res[14] [62], \aggregated_res[14] [61], 
      \aggregated_res[14] [60], \aggregated_res[14] [59], 
      \aggregated_res[14] [58], \aggregated_res[14] [57], 
      \aggregated_res[14] [56], \aggregated_res[14] [55], 
      \aggregated_res[14] [54], \aggregated_res[14] [53], 
      \aggregated_res[14] [52], \aggregated_res[14] [51], 
      \aggregated_res[14] [50], \aggregated_res[14] [49], 
      \aggregated_res[14] [48], \aggregated_res[14] [47], 
      \aggregated_res[14] [46], \aggregated_res[14] [45], 
      \aggregated_res[14] [44], \aggregated_res[14] [43], 
      \aggregated_res[14] [42], \aggregated_res[14] [41], 
      \aggregated_res[14] [40], \aggregated_res[14] [39], 
      \aggregated_res[14] [38], \aggregated_res[14] [37], 
      \aggregated_res[14] [36], \aggregated_res[14] [35], 
      \aggregated_res[14] [34], \aggregated_res[14] [33], 
      \aggregated_res[14] [32], \aggregated_res[14] [31], 
      \aggregated_res[14] [30], \aggregated_res[14] [29], 
      \aggregated_res[14] [28], \aggregated_res[14] [27], 
      \aggregated_res[14] [26], \aggregated_res[14] [25], 
      \aggregated_res[14] [24], \aggregated_res[14] [23], 
      \aggregated_res[14] [22], \aggregated_res[14] [21], 
      \aggregated_res[14] [20], \aggregated_res[14] [19], 
      \aggregated_res[14] [18], \aggregated_res[14] [17], 
      \aggregated_res[14] [16], \aggregated_res[14] [15], 
      \aggregated_res[14] [14], \aggregated_res[14] [13], 
      \aggregated_res[14] [12], \aggregated_res[14] [11], 
      \aggregated_res[14] [10], \aggregated_res[14] [9], \aggregated_res[14] [8], 
      \aggregated_res[14] [7], \aggregated_res[14] [6], \aggregated_res[14] [5], 
      \aggregated_res[14] [4], \aggregated_res[14] [3], \aggregated_res[14] [2], 
      n_0_813, n_0_812}), .p_0({n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, 
      n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, 
      n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, 
      n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, 
      n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, 
      n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, 
      n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, 
      n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, uc_503}));
   DLH_X1 \Res_reg[63]  (.D(n_0_250), .G(n_0_316), .Q(Res[63]));
   DLH_X1 \Res_reg[62]  (.D(n_0_249), .G(n_0_316), .Q(Res[62]));
   DLH_X1 \Res_reg[61]  (.D(n_0_248), .G(n_0_316), .Q(Res[61]));
   DLH_X1 \Res_reg[60]  (.D(n_0_247), .G(n_0_316), .Q(Res[60]));
   DLH_X1 \Res_reg[59]  (.D(n_0_246), .G(n_0_316), .Q(Res[59]));
   DLH_X1 \Res_reg[58]  (.D(n_0_245), .G(n_0_316), .Q(Res[58]));
   DLH_X1 \Res_reg[57]  (.D(n_0_244), .G(n_0_316), .Q(Res[57]));
   DLH_X1 \Res_reg[56]  (.D(n_0_243), .G(n_0_316), .Q(Res[56]));
   DLH_X1 \Res_reg[55]  (.D(n_0_242), .G(n_0_316), .Q(Res[55]));
   DLH_X1 \Res_reg[54]  (.D(n_0_241), .G(n_0_316), .Q(Res[54]));
   DLH_X1 \Res_reg[53]  (.D(n_0_240), .G(n_0_316), .Q(Res[53]));
   DLH_X1 \Res_reg[52]  (.D(n_0_239), .G(n_0_316), .Q(Res[52]));
   DLH_X1 \Res_reg[51]  (.D(n_0_238), .G(n_0_316), .Q(Res[51]));
   DLH_X1 \Res_reg[50]  (.D(n_0_237), .G(n_0_316), .Q(Res[50]));
   DLH_X1 \Res_reg[49]  (.D(n_0_236), .G(n_0_316), .Q(Res[49]));
   DLH_X1 \Res_reg[48]  (.D(n_0_235), .G(n_0_316), .Q(Res[48]));
   DLH_X1 \Res_reg[47]  (.D(n_0_234), .G(n_0_316), .Q(Res[47]));
   DLH_X1 \Res_reg[46]  (.D(n_0_233), .G(n_0_316), .Q(Res[46]));
   DLH_X1 \Res_reg[45]  (.D(n_0_232), .G(n_0_316), .Q(Res[45]));
   DLH_X1 \Res_reg[44]  (.D(n_0_231), .G(n_0_316), .Q(Res[44]));
   DLH_X1 \Res_reg[43]  (.D(n_0_230), .G(n_0_316), .Q(Res[43]));
   DLH_X1 \Res_reg[42]  (.D(n_0_229), .G(n_0_316), .Q(Res[42]));
   DLH_X1 \Res_reg[41]  (.D(n_0_228), .G(n_0_316), .Q(Res[41]));
   DLH_X1 \Res_reg[40]  (.D(n_0_227), .G(n_0_316), .Q(Res[40]));
   DLH_X1 \Res_reg[39]  (.D(n_0_226), .G(n_0_316), .Q(Res[39]));
   DLH_X1 \Res_reg[38]  (.D(n_0_225), .G(n_0_316), .Q(Res[38]));
   DLH_X1 \Res_reg[37]  (.D(n_0_224), .G(n_0_316), .Q(Res[37]));
   DLH_X1 \Res_reg[36]  (.D(n_0_223), .G(n_0_316), .Q(Res[36]));
   DLH_X1 \Res_reg[35]  (.D(n_0_222), .G(n_0_316), .Q(Res[35]));
   DLH_X1 \Res_reg[34]  (.D(n_0_221), .G(n_0_316), .Q(Res[34]));
   DLH_X1 \Res_reg[33]  (.D(n_0_220), .G(n_0_316), .Q(Res[33]));
   DLH_X1 \Res_reg[32]  (.D(n_0_219), .G(n_0_316), .Q(Res[32]));
   DLH_X1 \Res_reg[31]  (.D(n_0_218), .G(n_0_316), .Q(Res[31]));
   DLH_X1 \Res_reg[30]  (.D(n_0_217), .G(n_0_316), .Q(Res[30]));
   DLH_X1 \Res_reg[29]  (.D(n_0_216), .G(n_0_316), .Q(Res[29]));
   DLH_X1 \Res_reg[28]  (.D(n_0_215), .G(n_0_316), .Q(Res[28]));
   DLH_X1 \Res_reg[27]  (.D(n_0_214), .G(n_0_316), .Q(Res[27]));
   DLH_X1 \Res_reg[26]  (.D(n_0_213), .G(n_0_316), .Q(Res[26]));
   DLH_X1 \Res_reg[25]  (.D(n_0_212), .G(n_0_316), .Q(Res[25]));
   DLH_X1 \Res_reg[24]  (.D(n_0_211), .G(n_0_316), .Q(Res[24]));
   DLH_X1 \Res_reg[23]  (.D(n_0_210), .G(n_0_316), .Q(Res[23]));
   DLH_X1 \Res_reg[22]  (.D(n_0_209), .G(n_0_316), .Q(Res[22]));
   DLH_X1 \Res_reg[21]  (.D(n_0_208), .G(n_0_316), .Q(Res[21]));
   DLH_X1 \Res_reg[20]  (.D(n_0_207), .G(n_0_316), .Q(Res[20]));
   DLH_X1 \Res_reg[19]  (.D(n_0_206), .G(n_0_316), .Q(Res[19]));
   DLH_X1 \Res_reg[18]  (.D(n_0_205), .G(n_0_316), .Q(Res[18]));
   DLH_X1 \Res_reg[17]  (.D(n_0_204), .G(n_0_316), .Q(Res[17]));
   DLH_X1 \Res_reg[16]  (.D(n_0_203), .G(n_0_316), .Q(Res[16]));
   DLH_X1 \Res_reg[15]  (.D(n_0_202), .G(n_0_316), .Q(Res[15]));
   DLH_X1 \Res_reg[14]  (.D(n_0_201), .G(n_0_316), .Q(Res[14]));
   DLH_X1 \Res_reg[13]  (.D(n_0_200), .G(n_0_316), .Q(Res[13]));
   DLH_X1 \Res_reg[12]  (.D(n_0_199), .G(n_0_316), .Q(Res[12]));
   DLH_X1 \Res_reg[11]  (.D(n_0_198), .G(n_0_316), .Q(Res[11]));
   DLH_X1 \Res_reg[10]  (.D(n_0_197), .G(n_0_316), .Q(Res[10]));
   DLH_X1 \Res_reg[9]  (.D(n_0_196), .G(n_0_316), .Q(Res[9]));
   DLH_X1 \Res_reg[8]  (.D(n_0_195), .G(n_0_316), .Q(Res[8]));
   DLH_X1 \Res_reg[7]  (.D(n_0_194), .G(n_0_316), .Q(Res[7]));
   DLH_X1 \Res_reg[6]  (.D(n_0_193), .G(n_0_316), .Q(Res[6]));
   DLH_X1 \Res_reg[5]  (.D(n_0_192), .G(n_0_316), .Q(Res[5]));
   DLH_X1 \Res_reg[4]  (.D(n_0_191), .G(n_0_316), .Q(Res[4]));
   DLH_X1 \Res_reg[3]  (.D(n_0_190), .G(n_0_316), .Q(Res[3]));
   DLH_X1 \Res_reg[2]  (.D(n_0_189), .G(n_0_316), .Q(Res[2]));
   DLH_X1 \Res_reg[1]  (.D(n_0_188), .G(n_0_316), .Q(Res[1]));
   DLH_X1 \Res_reg[0]  (.D(n_0_187), .G(n_0_316), .Q(Res[0]));
   DLH_X1 \A_in_reg[31]  (.D(n_0_315), .G(n_0_283), .Q(A_in));
   DLH_X1 \A_in_reg[30]  (.D(n_0_314), .G(n_0_283), .Q(n_0_125));
   DLH_X1 \A_in_reg[29]  (.D(n_0_313), .G(n_0_283), .Q(n_0_126));
   DLH_X1 \A_in_reg[28]  (.D(n_0_312), .G(n_0_283), .Q(n_0_127));
   DLH_X1 \A_in_reg[27]  (.D(n_0_311), .G(n_0_283), .Q(n_0_128));
   DLH_X1 \A_in_reg[26]  (.D(n_0_310), .G(n_0_283), .Q(n_0_129));
   DLH_X1 \A_in_reg[25]  (.D(n_0_309), .G(n_0_283), .Q(n_0_130));
   DLH_X1 \A_in_reg[24]  (.D(n_0_308), .G(n_0_283), .Q(n_0_131));
   DLH_X1 \A_in_reg[23]  (.D(n_0_307), .G(n_0_283), .Q(n_0_132));
   DLH_X1 \A_in_reg[22]  (.D(n_0_306), .G(n_0_283), .Q(n_0_133));
   DLH_X1 \A_in_reg[21]  (.D(n_0_305), .G(n_0_283), .Q(n_0_134));
   DLH_X1 \A_in_reg[20]  (.D(n_0_304), .G(n_0_283), .Q(n_0_135));
   DLH_X1 \A_in_reg[19]  (.D(n_0_303), .G(n_0_283), .Q(n_0_136));
   DLH_X1 \A_in_reg[18]  (.D(n_0_302), .G(n_0_283), .Q(n_0_137));
   DLH_X1 \A_in_reg[17]  (.D(n_0_301), .G(n_0_283), .Q(n_0_138));
   DLH_X1 \A_in_reg[16]  (.D(n_0_300), .G(n_0_283), .Q(n_0_139));
   DLH_X1 \A_in_reg[15]  (.D(n_0_299), .G(n_0_283), .Q(n_0_140));
   DLH_X1 \A_in_reg[14]  (.D(n_0_298), .G(n_0_283), .Q(n_0_141));
   DLH_X1 \A_in_reg[13]  (.D(n_0_297), .G(n_0_283), .Q(n_0_142));
   DLH_X1 \A_in_reg[12]  (.D(n_0_296), .G(n_0_283), .Q(n_0_143));
   DLH_X1 \A_in_reg[11]  (.D(n_0_295), .G(n_0_283), .Q(n_0_144));
   DLH_X1 \A_in_reg[10]  (.D(n_0_294), .G(n_0_283), .Q(n_0_145));
   DLH_X1 \A_in_reg[9]  (.D(n_0_293), .G(n_0_283), .Q(n_0_146));
   DLH_X1 \A_in_reg[8]  (.D(n_0_292), .G(n_0_283), .Q(n_0_147));
   DLH_X1 \A_in_reg[7]  (.D(n_0_291), .G(n_0_283), .Q(n_0_148));
   DLH_X1 \A_in_reg[6]  (.D(n_0_290), .G(n_0_283), .Q(n_0_149));
   DLH_X1 \A_in_reg[5]  (.D(n_0_289), .G(n_0_283), .Q(n_0_150));
   DLH_X1 \A_in_reg[4]  (.D(n_0_288), .G(n_0_283), .Q(n_0_151));
   DLH_X1 \A_in_reg[3]  (.D(n_0_287), .G(n_0_283), .Q(n_0_152));
   DLH_X1 \A_in_reg[2]  (.D(n_0_286), .G(n_0_283), .Q(n_0_153));
   DLH_X1 \A_in_reg[1]  (.D(n_0_285), .G(n_0_283), .Q(n_0_154));
   DLH_X1 \A_in_reg[0]  (.D(n_0_284), .G(n_0_283), .Q(n_0_155));
   DLH_X1 \B_in_reg[31]  (.D(n_0_282), .G(n_0_283), .Q(B_in));
   DLH_X1 \B_in_reg[30]  (.D(n_0_281), .G(n_0_283), .Q(n_0_156));
   DLH_X1 \B_in_reg[29]  (.D(n_0_280), .G(n_0_283), .Q(n_0_157));
   DLH_X1 \B_in_reg[28]  (.D(n_0_279), .G(n_0_283), .Q(n_0_158));
   DLH_X1 \B_in_reg[27]  (.D(n_0_278), .G(n_0_283), .Q(n_0_159));
   DLH_X1 \B_in_reg[26]  (.D(n_0_277), .G(n_0_283), .Q(n_0_160));
   DLH_X1 \B_in_reg[25]  (.D(n_0_276), .G(n_0_283), .Q(n_0_161));
   DLH_X1 \B_in_reg[24]  (.D(n_0_275), .G(n_0_283), .Q(n_0_162));
   DLH_X1 \B_in_reg[23]  (.D(n_0_274), .G(n_0_283), .Q(n_0_163));
   DLH_X1 \B_in_reg[22]  (.D(n_0_273), .G(n_0_283), .Q(n_0_164));
   DLH_X1 \B_in_reg[21]  (.D(n_0_272), .G(n_0_283), .Q(n_0_165));
   DLH_X1 \B_in_reg[20]  (.D(n_0_271), .G(n_0_283), .Q(n_0_166));
   DLH_X1 \B_in_reg[19]  (.D(n_0_270), .G(n_0_283), .Q(n_0_167));
   DLH_X1 \B_in_reg[18]  (.D(n_0_269), .G(n_0_283), .Q(n_0_168));
   DLH_X1 \B_in_reg[17]  (.D(n_0_268), .G(n_0_283), .Q(n_0_169));
   DLH_X1 \B_in_reg[16]  (.D(n_0_267), .G(n_0_283), .Q(n_0_170));
   DLH_X1 \B_in_reg[15]  (.D(n_0_266), .G(n_0_283), .Q(n_0_171));
   DLH_X1 \B_in_reg[14]  (.D(n_0_265), .G(n_0_283), .Q(n_0_172));
   DLH_X1 \B_in_reg[13]  (.D(n_0_264), .G(n_0_283), .Q(n_0_173));
   DLH_X1 \B_in_reg[12]  (.D(n_0_263), .G(n_0_283), .Q(n_0_174));
   DLH_X1 \B_in_reg[11]  (.D(n_0_262), .G(n_0_283), .Q(n_0_175));
   DLH_X1 \B_in_reg[10]  (.D(n_0_261), .G(n_0_283), .Q(n_0_176));
   DLH_X1 \B_in_reg[9]  (.D(n_0_260), .G(n_0_283), .Q(n_0_177));
   DLH_X1 \B_in_reg[8]  (.D(n_0_259), .G(n_0_283), .Q(n_0_178));
   DLH_X1 \B_in_reg[7]  (.D(n_0_258), .G(n_0_283), .Q(n_0_179));
   DLH_X1 \B_in_reg[6]  (.D(n_0_257), .G(n_0_283), .Q(n_0_180));
   DLH_X1 \B_in_reg[5]  (.D(n_0_256), .G(n_0_283), .Q(n_0_181));
   DLH_X1 \B_in_reg[4]  (.D(n_0_255), .G(n_0_283), .Q(n_0_182));
   DLH_X1 \B_in_reg[3]  (.D(n_0_254), .G(n_0_283), .Q(n_0_183));
   DLH_X1 \B_in_reg[2]  (.D(n_0_253), .G(n_0_283), .Q(n_0_184));
   DLH_X1 \B_in_reg[1]  (.D(n_0_252), .G(n_0_283), .Q(n_0_185));
   DLH_X1 \B_in_reg[0]  (.D(n_0_251), .G(n_0_283), .Q(n_0_186));
   AND2_X1 i_0_1_0 (.A1(n_0_812), .A2(n_0_1_837), .ZN(n_0_187));
   NOR4_X1 i_0_1_138 (.A1(\aggregated_res[14] [28]), .A2(
      \aggregated_res[14] [27]), .A3(\aggregated_res[14] [26]), .A4(
      \aggregated_res[14] [25]), .ZN(n_0_1_74));
   NOR4_X1 i_0_1_139 (.A1(\aggregated_res[14] [63]), .A2(
      \aggregated_res[14] [30]), .A3(\aggregated_res[14] [29]), .A4(
      \aggregated_res[14] [23]), .ZN(n_0_1_75));
   NOR4_X1 i_0_1_140 (.A1(\aggregated_res[14] [20]), .A2(
      \aggregated_res[14] [19]), .A3(\aggregated_res[14] [18]), .A4(
      \aggregated_res[14] [17]), .ZN(n_0_1_76));
   NOR4_X1 i_0_1_141 (.A1(\aggregated_res[14] [24]), .A2(
      \aggregated_res[14] [22]), .A3(\aggregated_res[14] [21]), .A4(
      \aggregated_res[14] [16]), .ZN(n_0_1_77));
   NOR3_X1 i_0_1_143 (.A1(\aggregated_res[14] [45]), .A2(
      \aggregated_res[14] [39]), .A3(n_0_812), .ZN(n_0_1_79));
   NOR4_X1 i_0_1_144 (.A1(\aggregated_res[14] [44]), .A2(
      \aggregated_res[14] [43]), .A3(\aggregated_res[14] [42]), .A4(
      \aggregated_res[14] [41]), .ZN(n_0_1_80));
   NOR4_X1 i_0_1_145 (.A1(\aggregated_res[14] [36]), .A2(
      \aggregated_res[14] [35]), .A3(\aggregated_res[14] [34]), .A4(
      \aggregated_res[14] [33]), .ZN(n_0_1_81));
   NOR4_X1 i_0_1_146 (.A1(\aggregated_res[14] [46]), .A2(
      \aggregated_res[14] [40]), .A3(\aggregated_res[14] [38]), .A4(
      \aggregated_res[14] [37]), .ZN(n_0_1_82));
   AND2_X1 i_0_1_220 (.A1(n_0_1_131), .A2(n_0_155), .ZN(n_0_317));
   OAI211_X1 i_0_1_221 (.A(n_0_1_91), .B(n_0_1_90), .C1(n_0_1_776), .C2(
      n_0_1_129), .ZN(n_0_318));
   NAND2_X1 i_0_1_222 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_127), .ZN(n_0_1_90));
   OAI21_X1 i_0_1_223 (.A(n_0_155), .B1(n_0_1_124), .B2(n_0_1_123), .ZN(n_0_1_91));
   OAI221_X1 i_0_1_224 (.A(n_0_1_92), .B1(n_0_1_125), .B2(n_0_1_776), .C1(
      n_0_1_778), .C2(n_0_1_129), .ZN(n_0_319));
   AOI22_X1 i_0_1_225 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[1]), .ZN(n_0_1_92));
   OAI221_X1 i_0_1_226 (.A(n_0_1_93), .B1(n_0_1_125), .B2(n_0_1_778), .C1(
      n_0_1_780), .C2(n_0_1_129), .ZN(n_0_320));
   AOI22_X1 i_0_1_227 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[2]), .ZN(n_0_1_93));
   OAI221_X1 i_0_1_228 (.A(n_0_1_94), .B1(n_0_1_125), .B2(n_0_1_780), .C1(
      n_0_1_782), .C2(n_0_1_129), .ZN(n_0_321));
   AOI22_X1 i_0_1_229 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[3]), .ZN(n_0_1_94));
   OAI221_X1 i_0_1_230 (.A(n_0_1_95), .B1(n_0_1_125), .B2(n_0_1_782), .C1(
      n_0_1_784), .C2(n_0_1_129), .ZN(n_0_322));
   AOI22_X1 i_0_1_231 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[4]), .ZN(n_0_1_95));
   OAI221_X1 i_0_1_232 (.A(n_0_1_96), .B1(n_0_1_125), .B2(n_0_1_784), .C1(
      n_0_1_786), .C2(n_0_1_129), .ZN(n_0_323));
   AOI22_X1 i_0_1_233 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[5]), .ZN(n_0_1_96));
   OAI221_X1 i_0_1_234 (.A(n_0_1_97), .B1(n_0_1_125), .B2(n_0_1_786), .C1(
      n_0_1_788), .C2(n_0_1_129), .ZN(n_0_324));
   AOI22_X1 i_0_1_235 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[6]), .ZN(n_0_1_97));
   OAI221_X1 i_0_1_236 (.A(n_0_1_98), .B1(n_0_1_125), .B2(n_0_1_788), .C1(
      n_0_1_790), .C2(n_0_1_129), .ZN(n_0_325));
   AOI22_X1 i_0_1_237 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[7]), .ZN(n_0_1_98));
   OAI221_X1 i_0_1_238 (.A(n_0_1_99), .B1(n_0_1_125), .B2(n_0_1_790), .C1(
      n_0_1_792), .C2(n_0_1_129), .ZN(n_0_326));
   AOI22_X1 i_0_1_239 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[8]), .ZN(n_0_1_99));
   OAI221_X1 i_0_1_240 (.A(n_0_1_100), .B1(n_0_1_125), .B2(n_0_1_792), .C1(
      n_0_1_794), .C2(n_0_1_129), .ZN(n_0_327));
   AOI22_X1 i_0_1_241 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[9]), .ZN(n_0_1_100));
   OAI221_X1 i_0_1_242 (.A(n_0_1_101), .B1(n_0_1_125), .B2(n_0_1_794), .C1(
      n_0_1_796), .C2(n_0_1_129), .ZN(n_0_328));
   AOI22_X1 i_0_1_243 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[10]), .ZN(n_0_1_101));
   OAI221_X1 i_0_1_244 (.A(n_0_1_102), .B1(n_0_1_125), .B2(n_0_1_796), .C1(
      n_0_1_798), .C2(n_0_1_129), .ZN(n_0_329));
   AOI22_X1 i_0_1_245 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[11]), .ZN(n_0_1_102));
   OAI221_X1 i_0_1_246 (.A(n_0_1_103), .B1(n_0_1_125), .B2(n_0_1_798), .C1(
      n_0_1_800), .C2(n_0_1_129), .ZN(n_0_330));
   AOI22_X1 i_0_1_247 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[12]), .ZN(n_0_1_103));
   OAI221_X1 i_0_1_248 (.A(n_0_1_104), .B1(n_0_1_125), .B2(n_0_1_800), .C1(
      n_0_1_802), .C2(n_0_1_129), .ZN(n_0_331));
   AOI22_X1 i_0_1_249 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[13]), .ZN(n_0_1_104));
   OAI221_X1 i_0_1_250 (.A(n_0_1_105), .B1(n_0_1_125), .B2(n_0_1_802), .C1(
      n_0_1_804), .C2(n_0_1_129), .ZN(n_0_332));
   AOI22_X1 i_0_1_251 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[14]), .ZN(n_0_1_105));
   OAI221_X1 i_0_1_252 (.A(n_0_1_106), .B1(n_0_1_125), .B2(n_0_1_804), .C1(
      n_0_1_806), .C2(n_0_1_129), .ZN(n_0_333));
   AOI22_X1 i_0_1_253 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[15]), .ZN(n_0_1_106));
   OAI221_X1 i_0_1_254 (.A(n_0_1_107), .B1(n_0_1_125), .B2(n_0_1_806), .C1(
      n_0_1_808), .C2(n_0_1_129), .ZN(n_0_334));
   AOI22_X1 i_0_1_255 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[16]), .ZN(n_0_1_107));
   OAI221_X1 i_0_1_256 (.A(n_0_1_108), .B1(n_0_1_125), .B2(n_0_1_808), .C1(
      n_0_1_810), .C2(n_0_1_129), .ZN(n_0_335));
   AOI22_X1 i_0_1_257 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[17]), .ZN(n_0_1_108));
   OAI221_X1 i_0_1_258 (.A(n_0_1_109), .B1(n_0_1_125), .B2(n_0_1_810), .C1(
      n_0_1_812), .C2(n_0_1_129), .ZN(n_0_336));
   AOI22_X1 i_0_1_259 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[18]), .ZN(n_0_1_109));
   OAI221_X1 i_0_1_260 (.A(n_0_1_110), .B1(n_0_1_125), .B2(n_0_1_812), .C1(
      n_0_1_814), .C2(n_0_1_129), .ZN(n_0_337));
   AOI22_X1 i_0_1_261 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[19]), .ZN(n_0_1_110));
   OAI221_X1 i_0_1_262 (.A(n_0_1_111), .B1(n_0_1_125), .B2(n_0_1_814), .C1(
      n_0_1_816), .C2(n_0_1_129), .ZN(n_0_338));
   AOI22_X1 i_0_1_263 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[20]), .ZN(n_0_1_111));
   OAI221_X1 i_0_1_264 (.A(n_0_1_112), .B1(n_0_1_125), .B2(n_0_1_816), .C1(
      n_0_1_818), .C2(n_0_1_129), .ZN(n_0_339));
   AOI22_X1 i_0_1_265 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[21]), .ZN(n_0_1_112));
   OAI221_X1 i_0_1_266 (.A(n_0_1_113), .B1(n_0_1_125), .B2(n_0_1_818), .C1(
      n_0_1_820), .C2(n_0_1_129), .ZN(n_0_340));
   AOI22_X1 i_0_1_267 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[22]), .ZN(n_0_1_113));
   OAI221_X1 i_0_1_268 (.A(n_0_1_114), .B1(n_0_1_125), .B2(n_0_1_820), .C1(
      n_0_1_822), .C2(n_0_1_129), .ZN(n_0_341));
   AOI22_X1 i_0_1_269 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[23]), .ZN(n_0_1_114));
   OAI221_X1 i_0_1_270 (.A(n_0_1_115), .B1(n_0_1_125), .B2(n_0_1_822), .C1(
      n_0_1_824), .C2(n_0_1_129), .ZN(n_0_342));
   AOI22_X1 i_0_1_271 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[24]), .ZN(n_0_1_115));
   OAI221_X1 i_0_1_272 (.A(n_0_1_116), .B1(n_0_1_125), .B2(n_0_1_824), .C1(
      n_0_1_826), .C2(n_0_1_129), .ZN(n_0_343));
   AOI22_X1 i_0_1_273 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[25]), .ZN(n_0_1_116));
   OAI221_X1 i_0_1_274 (.A(n_0_1_117), .B1(n_0_1_125), .B2(n_0_1_826), .C1(
      n_0_1_828), .C2(n_0_1_129), .ZN(n_0_344));
   AOI22_X1 i_0_1_275 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[26]), .ZN(n_0_1_117));
   OAI221_X1 i_0_1_276 (.A(n_0_1_118), .B1(n_0_1_125), .B2(n_0_1_828), .C1(
      n_0_1_830), .C2(n_0_1_129), .ZN(n_0_345));
   AOI22_X1 i_0_1_277 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[27]), .ZN(n_0_1_118));
   OAI221_X1 i_0_1_278 (.A(n_0_1_119), .B1(n_0_1_125), .B2(n_0_1_830), .C1(
      n_0_1_832), .C2(n_0_1_129), .ZN(n_0_346));
   AOI22_X1 i_0_1_279 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[28]), .ZN(n_0_1_119));
   OAI221_X1 i_0_1_280 (.A(n_0_1_120), .B1(n_0_1_125), .B2(n_0_1_832), .C1(
      n_0_1_834), .C2(n_0_1_129), .ZN(n_0_347));
   AOI22_X1 i_0_1_281 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_127), .B1(
      n_0_1_123), .B2(A_imm_2s_complement[29]), .ZN(n_0_1_120));
   NAND2_X1 i_0_1_282 (.A1(n_0_1_126), .A2(n_0_1_121), .ZN(n_0_348));
   AOI22_X1 i_0_1_283 (.A1(n_0_1_124), .A2(A_imm[30]), .B1(
      A_imm_2s_complement[30]), .B2(n_0_1_123), .ZN(n_0_1_121));
   OAI211_X1 i_0_1_284 (.A(n_0_1_126), .B(n_0_1_122), .C1(n_0_1_125), .C2(
      n_0_1_836), .ZN(n_0_349));
   NAND2_X1 i_0_1_285 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_123), .ZN(
      n_0_1_122));
   NOR3_X1 i_0_1_286 (.A1(n_0_1_133), .A2(n_0_59), .A3(n_0_60), .ZN(n_0_1_123));
   INV_X1 i_0_1_287 (.A(n_0_1_125), .ZN(n_0_1_124));
   NAND3_X1 i_0_1_288 (.A1(n_0_1_174), .A2(n_0_1_133), .A3(n_0_1_132), .ZN(
      n_0_1_125));
   AOI21_X1 i_0_1_289 (.A(n_0_1_128), .B1(n_0_1_127), .B2(
      A_imm_2s_complement[31]), .ZN(n_0_1_126));
   NOR2_X1 i_0_1_290 (.A1(n_0_1_130), .A2(n_0_1_133), .ZN(n_0_1_127));
   NOR2_X1 i_0_1_291 (.A1(n_0_1_129), .A2(n_0_1_836), .ZN(n_0_1_128));
   NAND2_X1 i_0_1_292 (.A1(n_0_1_133), .A2(n_0_1_131), .ZN(n_0_1_129));
   INV_X1 i_0_1_293 (.A(n_0_1_131), .ZN(n_0_1_130));
   XNOR2_X1 i_0_1_294 (.A(n_0_1_175), .B(n_0_1_132), .ZN(n_0_1_131));
   MUX2_X1 i_0_1_295 (.A(n_0_156), .B(n_0_60), .S(B_in), .Z(n_0_1_132));
   NAND2_X1 i_0_1_296 (.A1(B_in), .A2(n_0_61), .ZN(n_0_1_133));
   AND2_X1 i_0_1_297 (.A1(n_0_1_169), .A2(n_0_155), .ZN(n_0_350));
   OAI211_X1 i_0_1_298 (.A(n_0_1_135), .B(n_0_1_134), .C1(n_0_1_776), .C2(
      n_0_1_165), .ZN(n_0_351));
   OAI21_X1 i_0_1_299 (.A(n_0_155), .B1(n_0_1_170), .B2(n_0_1_167), .ZN(
      n_0_1_134));
   NAND2_X1 i_0_1_300 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_168), .ZN(
      n_0_1_135));
   OAI21_X1 i_0_1_301 (.A(n_0_1_136), .B1(n_0_1_165), .B2(n_0_1_778), .ZN(
      n_0_352));
   AOI222_X1 i_0_1_302 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[1]), .C1(A_imm[1]), .C2(n_0_1_170), 
      .ZN(n_0_1_136));
   OAI21_X1 i_0_1_303 (.A(n_0_1_137), .B1(n_0_1_165), .B2(n_0_1_780), .ZN(
      n_0_353));
   AOI222_X1 i_0_1_304 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[2]), .C1(A_imm[2]), .C2(n_0_1_170), 
      .ZN(n_0_1_137));
   OAI21_X1 i_0_1_305 (.A(n_0_1_138), .B1(n_0_1_165), .B2(n_0_1_782), .ZN(
      n_0_354));
   AOI222_X1 i_0_1_306 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[3]), .C1(A_imm[3]), .C2(n_0_1_170), 
      .ZN(n_0_1_138));
   OAI21_X1 i_0_1_307 (.A(n_0_1_139), .B1(n_0_1_165), .B2(n_0_1_784), .ZN(
      n_0_355));
   AOI222_X1 i_0_1_308 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[4]), .C1(A_imm[4]), .C2(n_0_1_170), 
      .ZN(n_0_1_139));
   OAI21_X1 i_0_1_309 (.A(n_0_1_140), .B1(n_0_1_165), .B2(n_0_1_786), .ZN(
      n_0_356));
   AOI222_X1 i_0_1_310 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[5]), .C1(A_imm[5]), .C2(n_0_1_170), 
      .ZN(n_0_1_140));
   OAI21_X1 i_0_1_311 (.A(n_0_1_141), .B1(n_0_1_165), .B2(n_0_1_788), .ZN(
      n_0_357));
   AOI222_X1 i_0_1_312 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[6]), .C1(A_imm[6]), .C2(n_0_1_170), 
      .ZN(n_0_1_141));
   OAI21_X1 i_0_1_313 (.A(n_0_1_142), .B1(n_0_1_165), .B2(n_0_1_790), .ZN(
      n_0_358));
   AOI222_X1 i_0_1_314 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[7]), .C1(A_imm[7]), .C2(n_0_1_170), 
      .ZN(n_0_1_142));
   OAI21_X1 i_0_1_315 (.A(n_0_1_143), .B1(n_0_1_165), .B2(n_0_1_792), .ZN(
      n_0_359));
   AOI222_X1 i_0_1_316 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[8]), .C1(A_imm[8]), .C2(n_0_1_170), 
      .ZN(n_0_1_143));
   OAI21_X1 i_0_1_317 (.A(n_0_1_144), .B1(n_0_1_165), .B2(n_0_1_794), .ZN(
      n_0_360));
   AOI222_X1 i_0_1_318 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[9]), .C1(A_imm[9]), .C2(n_0_1_170), 
      .ZN(n_0_1_144));
   OAI21_X1 i_0_1_319 (.A(n_0_1_145), .B1(n_0_1_165), .B2(n_0_1_796), .ZN(
      n_0_361));
   AOI222_X1 i_0_1_320 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[10]), .C1(A_imm[10]), .C2(n_0_1_170), 
      .ZN(n_0_1_145));
   OAI21_X1 i_0_1_321 (.A(n_0_1_146), .B1(n_0_1_165), .B2(n_0_1_798), .ZN(
      n_0_362));
   AOI222_X1 i_0_1_322 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[11]), .C1(A_imm[11]), .C2(n_0_1_170), 
      .ZN(n_0_1_146));
   OAI21_X1 i_0_1_323 (.A(n_0_1_147), .B1(n_0_1_165), .B2(n_0_1_800), .ZN(
      n_0_363));
   AOI222_X1 i_0_1_324 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[12]), .C1(A_imm[12]), .C2(n_0_1_170), 
      .ZN(n_0_1_147));
   OAI21_X1 i_0_1_325 (.A(n_0_1_148), .B1(n_0_1_165), .B2(n_0_1_802), .ZN(
      n_0_364));
   AOI222_X1 i_0_1_326 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[13]), .C1(A_imm[13]), .C2(n_0_1_170), 
      .ZN(n_0_1_148));
   OAI21_X1 i_0_1_327 (.A(n_0_1_149), .B1(n_0_1_165), .B2(n_0_1_804), .ZN(
      n_0_365));
   AOI222_X1 i_0_1_328 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[14]), .C1(A_imm[14]), .C2(n_0_1_170), 
      .ZN(n_0_1_149));
   OAI21_X1 i_0_1_329 (.A(n_0_1_150), .B1(n_0_1_165), .B2(n_0_1_806), .ZN(
      n_0_366));
   AOI222_X1 i_0_1_330 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[15]), .C1(A_imm[15]), .C2(n_0_1_170), 
      .ZN(n_0_1_150));
   OAI21_X1 i_0_1_331 (.A(n_0_1_151), .B1(n_0_1_165), .B2(n_0_1_808), .ZN(
      n_0_367));
   AOI222_X1 i_0_1_332 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[16]), .C1(A_imm[16]), .C2(n_0_1_170), 
      .ZN(n_0_1_151));
   OAI21_X1 i_0_1_333 (.A(n_0_1_152), .B1(n_0_1_165), .B2(n_0_1_810), .ZN(
      n_0_368));
   AOI222_X1 i_0_1_334 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[17]), .C1(A_imm[17]), .C2(n_0_1_170), 
      .ZN(n_0_1_152));
   OAI21_X1 i_0_1_335 (.A(n_0_1_153), .B1(n_0_1_165), .B2(n_0_1_812), .ZN(
      n_0_369));
   AOI222_X1 i_0_1_336 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[18]), .C1(A_imm[18]), .C2(n_0_1_170), 
      .ZN(n_0_1_153));
   OAI21_X1 i_0_1_337 (.A(n_0_1_154), .B1(n_0_1_165), .B2(n_0_1_814), .ZN(
      n_0_370));
   AOI222_X1 i_0_1_338 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[19]), .C1(A_imm[19]), .C2(n_0_1_170), 
      .ZN(n_0_1_154));
   OAI21_X1 i_0_1_339 (.A(n_0_1_155), .B1(n_0_1_165), .B2(n_0_1_816), .ZN(
      n_0_371));
   AOI222_X1 i_0_1_340 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[20]), .C1(A_imm[20]), .C2(n_0_1_170), 
      .ZN(n_0_1_155));
   OAI21_X1 i_0_1_341 (.A(n_0_1_156), .B1(n_0_1_165), .B2(n_0_1_818), .ZN(
      n_0_372));
   AOI222_X1 i_0_1_342 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[21]), .C1(A_imm[21]), .C2(n_0_1_170), 
      .ZN(n_0_1_156));
   OAI21_X1 i_0_1_343 (.A(n_0_1_157), .B1(n_0_1_165), .B2(n_0_1_820), .ZN(
      n_0_373));
   AOI222_X1 i_0_1_344 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[22]), .C1(A_imm[22]), .C2(n_0_1_170), 
      .ZN(n_0_1_157));
   OAI21_X1 i_0_1_345 (.A(n_0_1_158), .B1(n_0_1_165), .B2(n_0_1_822), .ZN(
      n_0_374));
   AOI222_X1 i_0_1_346 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[23]), .C1(A_imm[23]), .C2(n_0_1_170), 
      .ZN(n_0_1_158));
   OAI21_X1 i_0_1_347 (.A(n_0_1_159), .B1(n_0_1_165), .B2(n_0_1_824), .ZN(
      n_0_375));
   AOI222_X1 i_0_1_348 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[24]), .C1(A_imm[24]), .C2(n_0_1_170), 
      .ZN(n_0_1_159));
   OAI21_X1 i_0_1_349 (.A(n_0_1_160), .B1(n_0_1_165), .B2(n_0_1_826), .ZN(
      n_0_376));
   AOI222_X1 i_0_1_350 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[25]), .C1(A_imm[25]), .C2(n_0_1_170), 
      .ZN(n_0_1_160));
   OAI21_X1 i_0_1_351 (.A(n_0_1_161), .B1(n_0_1_165), .B2(n_0_1_828), .ZN(
      n_0_377));
   AOI222_X1 i_0_1_352 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[26]), .C1(A_imm[26]), .C2(n_0_1_170), 
      .ZN(n_0_1_161));
   OAI21_X1 i_0_1_353 (.A(n_0_1_162), .B1(n_0_1_165), .B2(n_0_1_830), .ZN(
      n_0_378));
   AOI222_X1 i_0_1_354 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[27]), .C1(A_imm[27]), .C2(n_0_1_170), 
      .ZN(n_0_1_162));
   OAI21_X1 i_0_1_355 (.A(n_0_1_163), .B1(n_0_1_165), .B2(n_0_1_832), .ZN(
      n_0_379));
   AOI222_X1 i_0_1_356 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[28]), .C1(A_imm[28]), .C2(n_0_1_170), 
      .ZN(n_0_1_163));
   OAI21_X1 i_0_1_357 (.A(n_0_1_164), .B1(n_0_1_165), .B2(n_0_1_834), .ZN(
      n_0_380));
   AOI222_X1 i_0_1_358 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[29]), .C1(A_imm[29]), .C2(n_0_1_170), 
      .ZN(n_0_1_164));
   OAI21_X1 i_0_1_359 (.A(n_0_1_166), .B1(n_0_1_165), .B2(n_0_1_836), .ZN(
      n_0_381));
   NAND2_X1 i_0_1_360 (.A1(n_0_1_169), .A2(n_0_1_175), .ZN(n_0_1_165));
   AOI222_X1 i_0_1_361 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_168), .B1(
      n_0_1_167), .B2(A_imm_2s_complement[30]), .C1(A_imm[30]), .C2(n_0_1_170), 
      .ZN(n_0_1_166));
   NOR2_X1 i_0_1_362 (.A1(n_0_1_172), .A2(n_0_1_175), .ZN(n_0_1_167));
   AND2_X1 i_0_1_363 (.A1(n_0_1_174), .A2(n_0_1_169), .ZN(n_0_1_168));
   XNOR2_X1 i_0_1_364 (.A(n_0_1_219), .B(n_0_1_179), .ZN(n_0_1_169));
   NOR2_X1 i_0_1_365 (.A1(n_0_1_178), .A2(n_0_1_174), .ZN(n_0_1_170));
   NAND2_X1 i_0_1_366 (.A1(n_0_1_173), .A2(n_0_1_171), .ZN(n_0_382));
   NAND3_X1 i_0_1_367 (.A1(n_0_1_172), .A2(n_0_1_175), .A3(A_imm[31]), .ZN(
      n_0_1_171));
   OR2_X1 i_0_1_368 (.A1(n_0_1_220), .A2(n_0_1_179), .ZN(n_0_1_172));
   NAND3_X1 i_0_1_369 (.A1(n_0_1_178), .A2(n_0_1_174), .A3(
      A_imm_2s_complement[31]), .ZN(n_0_1_173));
   OAI21_X1 i_0_1_370 (.A(n_0_1_177), .B1(n_0_1_868), .B2(B_in), .ZN(n_0_1_174));
   AOI21_X1 i_0_1_371 (.A(n_0_1_176), .B1(n_0_59), .B2(B_in), .ZN(n_0_1_175));
   NOR2_X1 i_0_1_372 (.A1(n_0_1_868), .A2(B_in), .ZN(n_0_1_176));
   NAND2_X1 i_0_1_373 (.A1(B_in), .A2(n_0_59), .ZN(n_0_1_177));
   NAND2_X1 i_0_1_374 (.A1(n_0_1_220), .A2(n_0_1_179), .ZN(n_0_1_178));
   MUX2_X1 i_0_1_375 (.A(n_0_158), .B(n_0_58), .S(B_in), .Z(n_0_1_179));
   AND2_X1 i_0_1_376 (.A1(n_0_1_216), .A2(n_0_155), .ZN(n_0_383));
   OAI211_X1 i_0_1_377 (.A(n_0_1_181), .B(n_0_1_180), .C1(n_0_1_776), .C2(
      n_0_1_213), .ZN(n_0_384));
   OAI21_X1 i_0_1_378 (.A(n_0_155), .B1(n_0_1_214), .B2(n_0_1_212), .ZN(
      n_0_1_180));
   NAND2_X1 i_0_1_379 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_215), .ZN(
      n_0_1_181));
   OAI21_X1 i_0_1_380 (.A(n_0_1_182), .B1(n_0_1_213), .B2(n_0_1_778), .ZN(
      n_0_385));
   AOI222_X1 i_0_1_381 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[1]), .C1(n_0_1_212), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_182));
   OAI21_X1 i_0_1_382 (.A(n_0_1_183), .B1(n_0_1_213), .B2(n_0_1_780), .ZN(
      n_0_386));
   AOI222_X1 i_0_1_383 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[2]), .C1(n_0_1_212), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_183));
   OAI21_X1 i_0_1_384 (.A(n_0_1_184), .B1(n_0_1_213), .B2(n_0_1_782), .ZN(
      n_0_387));
   AOI222_X1 i_0_1_385 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[3]), .C1(n_0_1_212), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_184));
   OAI21_X1 i_0_1_386 (.A(n_0_1_185), .B1(n_0_1_213), .B2(n_0_1_784), .ZN(
      n_0_388));
   AOI222_X1 i_0_1_387 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[4]), .C1(n_0_1_212), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_185));
   OAI21_X1 i_0_1_388 (.A(n_0_1_186), .B1(n_0_1_213), .B2(n_0_1_786), .ZN(
      n_0_389));
   AOI222_X1 i_0_1_389 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[5]), .C1(n_0_1_212), .C2(A_imm_2s_complement[5]), 
      .ZN(n_0_1_186));
   OAI21_X1 i_0_1_390 (.A(n_0_1_187), .B1(n_0_1_213), .B2(n_0_1_788), .ZN(
      n_0_390));
   AOI222_X1 i_0_1_391 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[6]), .C1(n_0_1_212), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_187));
   OAI21_X1 i_0_1_392 (.A(n_0_1_188), .B1(n_0_1_213), .B2(n_0_1_790), .ZN(
      n_0_391));
   AOI222_X1 i_0_1_393 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[7]), .C1(n_0_1_212), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_188));
   OAI21_X1 i_0_1_394 (.A(n_0_1_189), .B1(n_0_1_213), .B2(n_0_1_792), .ZN(
      n_0_392));
   AOI222_X1 i_0_1_395 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[8]), .C1(n_0_1_212), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_189));
   OAI21_X1 i_0_1_396 (.A(n_0_1_190), .B1(n_0_1_213), .B2(n_0_1_794), .ZN(
      n_0_393));
   AOI222_X1 i_0_1_397 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[9]), .C1(n_0_1_212), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_190));
   OAI21_X1 i_0_1_398 (.A(n_0_1_191), .B1(n_0_1_213), .B2(n_0_1_796), .ZN(
      n_0_394));
   AOI222_X1 i_0_1_399 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[10]), .C1(n_0_1_212), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_191));
   OAI21_X1 i_0_1_400 (.A(n_0_1_192), .B1(n_0_1_213), .B2(n_0_1_798), .ZN(
      n_0_395));
   AOI222_X1 i_0_1_401 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[11]), .C1(n_0_1_212), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_192));
   OAI21_X1 i_0_1_402 (.A(n_0_1_193), .B1(n_0_1_213), .B2(n_0_1_800), .ZN(
      n_0_396));
   AOI222_X1 i_0_1_403 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[12]), .C1(n_0_1_212), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_193));
   OAI21_X1 i_0_1_404 (.A(n_0_1_194), .B1(n_0_1_213), .B2(n_0_1_802), .ZN(
      n_0_397));
   AOI222_X1 i_0_1_405 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[13]), .C1(n_0_1_212), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_194));
   OAI21_X1 i_0_1_406 (.A(n_0_1_195), .B1(n_0_1_213), .B2(n_0_1_804), .ZN(
      n_0_398));
   AOI222_X1 i_0_1_407 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[14]), .C1(n_0_1_212), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_195));
   OAI21_X1 i_0_1_408 (.A(n_0_1_196), .B1(n_0_1_213), .B2(n_0_1_806), .ZN(
      n_0_399));
   AOI222_X1 i_0_1_409 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[15]), .C1(n_0_1_212), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_196));
   OAI21_X1 i_0_1_410 (.A(n_0_1_197), .B1(n_0_1_213), .B2(n_0_1_808), .ZN(
      n_0_400));
   AOI222_X1 i_0_1_411 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[16]), .C1(n_0_1_212), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_197));
   OAI21_X1 i_0_1_412 (.A(n_0_1_198), .B1(n_0_1_213), .B2(n_0_1_810), .ZN(
      n_0_401));
   AOI222_X1 i_0_1_413 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[17]), .C1(n_0_1_212), .C2(A_imm_2s_complement[17]), 
      .ZN(n_0_1_198));
   OAI21_X1 i_0_1_414 (.A(n_0_1_199), .B1(n_0_1_213), .B2(n_0_1_812), .ZN(
      n_0_402));
   AOI222_X1 i_0_1_415 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[18]), .C1(n_0_1_212), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_199));
   OAI21_X1 i_0_1_416 (.A(n_0_1_200), .B1(n_0_1_213), .B2(n_0_1_814), .ZN(
      n_0_403));
   AOI222_X1 i_0_1_417 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[19]), .C1(n_0_1_212), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_200));
   OAI21_X1 i_0_1_418 (.A(n_0_1_201), .B1(n_0_1_213), .B2(n_0_1_816), .ZN(
      n_0_404));
   AOI222_X1 i_0_1_419 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[20]), .C1(n_0_1_212), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_201));
   OAI21_X1 i_0_1_420 (.A(n_0_1_202), .B1(n_0_1_213), .B2(n_0_1_818), .ZN(
      n_0_405));
   AOI222_X1 i_0_1_421 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[21]), .C1(n_0_1_212), .C2(A_imm_2s_complement[21]), 
      .ZN(n_0_1_202));
   OAI21_X1 i_0_1_422 (.A(n_0_1_203), .B1(n_0_1_213), .B2(n_0_1_820), .ZN(
      n_0_406));
   AOI222_X1 i_0_1_423 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[22]), .C1(n_0_1_212), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_203));
   OAI21_X1 i_0_1_424 (.A(n_0_1_204), .B1(n_0_1_213), .B2(n_0_1_822), .ZN(
      n_0_407));
   AOI222_X1 i_0_1_425 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[23]), .C1(n_0_1_212), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_204));
   OAI21_X1 i_0_1_426 (.A(n_0_1_205), .B1(n_0_1_213), .B2(n_0_1_824), .ZN(
      n_0_408));
   AOI222_X1 i_0_1_427 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[24]), .C1(n_0_1_212), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_205));
   OAI21_X1 i_0_1_428 (.A(n_0_1_206), .B1(n_0_1_213), .B2(n_0_1_826), .ZN(
      n_0_409));
   AOI222_X1 i_0_1_429 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[25]), .C1(n_0_1_212), .C2(A_imm_2s_complement[25]), 
      .ZN(n_0_1_206));
   OAI21_X1 i_0_1_430 (.A(n_0_1_207), .B1(n_0_1_213), .B2(n_0_1_828), .ZN(
      n_0_410));
   AOI222_X1 i_0_1_431 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[26]), .C1(n_0_1_212), .C2(A_imm_2s_complement[26]), 
      .ZN(n_0_1_207));
   OAI21_X1 i_0_1_432 (.A(n_0_1_208), .B1(n_0_1_213), .B2(n_0_1_830), .ZN(
      n_0_411));
   AOI222_X1 i_0_1_433 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[27]), .C1(n_0_1_212), .C2(A_imm_2s_complement[27]), 
      .ZN(n_0_1_208));
   OAI21_X1 i_0_1_434 (.A(n_0_1_209), .B1(n_0_1_213), .B2(n_0_1_832), .ZN(
      n_0_412));
   AOI222_X1 i_0_1_435 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[28]), .C1(n_0_1_212), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_209));
   OAI21_X1 i_0_1_436 (.A(n_0_1_210), .B1(n_0_1_213), .B2(n_0_1_834), .ZN(
      n_0_413));
   AOI222_X1 i_0_1_437 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[29]), .C1(n_0_1_212), .C2(A_imm_2s_complement[29]), 
      .ZN(n_0_1_210));
   OAI21_X1 i_0_1_438 (.A(n_0_1_211), .B1(n_0_1_213), .B2(n_0_1_836), .ZN(
      n_0_414));
   AOI222_X1 i_0_1_439 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_215), .B1(
      n_0_1_214), .B2(A_imm[30]), .C1(n_0_1_212), .C2(A_imm_2s_complement[30]), 
      .ZN(n_0_1_211));
   NOR3_X1 i_0_1_440 (.A1(n_0_1_219), .A2(n_0_1_222), .A3(n_0_1_263), .ZN(
      n_0_1_212));
   NAND2_X1 i_0_1_441 (.A1(n_0_1_216), .A2(n_0_1_219), .ZN(n_0_1_213));
   NOR2_X1 i_0_1_442 (.A1(n_0_1_221), .A2(n_0_1_220), .ZN(n_0_1_214));
   AND2_X1 i_0_1_443 (.A1(n_0_1_220), .A2(n_0_1_216), .ZN(n_0_1_215));
   XNOR2_X1 i_0_1_444 (.A(n_0_1_262), .B(n_0_1_222), .ZN(n_0_1_216));
   OAI21_X1 i_0_1_445 (.A(n_0_1_218), .B1(n_0_1_217), .B2(n_0_1_220), .ZN(
      n_0_415));
   OAI21_X1 i_0_1_446 (.A(A_imm[31]), .B1(n_0_1_263), .B2(n_0_1_222), .ZN(
      n_0_1_217));
   NAND3_X1 i_0_1_447 (.A1(n_0_1_221), .A2(n_0_1_220), .A3(
      A_imm_2s_complement[31]), .ZN(n_0_1_218));
   INV_X1 i_0_1_448 (.A(n_0_1_220), .ZN(n_0_1_219));
   MUX2_X1 i_0_1_449 (.A(n_0_159), .B(n_0_57), .S(B_in), .Z(n_0_1_220));
   NAND2_X1 i_0_1_450 (.A1(n_0_1_263), .A2(n_0_1_222), .ZN(n_0_1_221));
   MUX2_X1 i_0_1_451 (.A(n_0_160), .B(n_0_56), .S(B_in), .Z(n_0_1_222));
   AND2_X1 i_0_1_452 (.A1(n_0_1_259), .A2(n_0_155), .ZN(n_0_416));
   OAI211_X1 i_0_1_453 (.A(n_0_1_224), .B(n_0_1_223), .C1(n_0_1_776), .C2(
      n_0_1_256), .ZN(n_0_417));
   OAI21_X1 i_0_1_454 (.A(n_0_155), .B1(n_0_1_257), .B2(n_0_1_255), .ZN(
      n_0_1_223));
   NAND2_X1 i_0_1_455 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_258), .ZN(
      n_0_1_224));
   OAI21_X1 i_0_1_456 (.A(n_0_1_225), .B1(n_0_1_256), .B2(n_0_1_778), .ZN(
      n_0_418));
   AOI222_X1 i_0_1_457 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[1]), .C1(n_0_1_255), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_225));
   OAI21_X1 i_0_1_458 (.A(n_0_1_226), .B1(n_0_1_256), .B2(n_0_1_780), .ZN(
      n_0_419));
   AOI222_X1 i_0_1_459 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[2]), .C1(n_0_1_255), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_226));
   OAI21_X1 i_0_1_460 (.A(n_0_1_227), .B1(n_0_1_256), .B2(n_0_1_782), .ZN(
      n_0_420));
   AOI222_X1 i_0_1_461 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[3]), .C1(n_0_1_255), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_227));
   OAI21_X1 i_0_1_462 (.A(n_0_1_228), .B1(n_0_1_256), .B2(n_0_1_784), .ZN(
      n_0_421));
   AOI222_X1 i_0_1_463 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[4]), .C1(n_0_1_255), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_228));
   OAI21_X1 i_0_1_464 (.A(n_0_1_229), .B1(n_0_1_256), .B2(n_0_1_786), .ZN(
      n_0_422));
   AOI222_X1 i_0_1_465 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[5]), .C1(n_0_1_255), .C2(A_imm_2s_complement[5]), 
      .ZN(n_0_1_229));
   OAI21_X1 i_0_1_466 (.A(n_0_1_230), .B1(n_0_1_256), .B2(n_0_1_788), .ZN(
      n_0_423));
   AOI222_X1 i_0_1_467 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[6]), .C1(n_0_1_255), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_230));
   OAI21_X1 i_0_1_468 (.A(n_0_1_231), .B1(n_0_1_256), .B2(n_0_1_790), .ZN(
      n_0_424));
   AOI222_X1 i_0_1_469 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[7]), .C1(n_0_1_255), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_231));
   OAI21_X1 i_0_1_470 (.A(n_0_1_232), .B1(n_0_1_256), .B2(n_0_1_792), .ZN(
      n_0_425));
   AOI222_X1 i_0_1_471 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[8]), .C1(n_0_1_255), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_232));
   OAI21_X1 i_0_1_472 (.A(n_0_1_233), .B1(n_0_1_256), .B2(n_0_1_794), .ZN(
      n_0_426));
   AOI222_X1 i_0_1_473 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[9]), .C1(n_0_1_255), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_233));
   OAI21_X1 i_0_1_474 (.A(n_0_1_234), .B1(n_0_1_256), .B2(n_0_1_796), .ZN(
      n_0_427));
   AOI222_X1 i_0_1_475 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[10]), .C1(n_0_1_255), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_234));
   OAI21_X1 i_0_1_476 (.A(n_0_1_235), .B1(n_0_1_256), .B2(n_0_1_798), .ZN(
      n_0_428));
   AOI222_X1 i_0_1_477 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[11]), .C1(n_0_1_255), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_235));
   OAI21_X1 i_0_1_478 (.A(n_0_1_236), .B1(n_0_1_256), .B2(n_0_1_800), .ZN(
      n_0_429));
   AOI222_X1 i_0_1_479 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[12]), .C1(n_0_1_255), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_236));
   OAI21_X1 i_0_1_480 (.A(n_0_1_237), .B1(n_0_1_256), .B2(n_0_1_802), .ZN(
      n_0_430));
   AOI222_X1 i_0_1_481 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[13]), .C1(n_0_1_255), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_237));
   OAI21_X1 i_0_1_482 (.A(n_0_1_238), .B1(n_0_1_256), .B2(n_0_1_804), .ZN(
      n_0_431));
   AOI222_X1 i_0_1_483 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[14]), .C1(n_0_1_255), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_238));
   OAI21_X1 i_0_1_484 (.A(n_0_1_239), .B1(n_0_1_256), .B2(n_0_1_806), .ZN(
      n_0_432));
   AOI222_X1 i_0_1_485 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[15]), .C1(n_0_1_255), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_239));
   OAI21_X1 i_0_1_486 (.A(n_0_1_240), .B1(n_0_1_256), .B2(n_0_1_808), .ZN(
      n_0_433));
   AOI222_X1 i_0_1_487 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[16]), .C1(n_0_1_255), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_240));
   OAI21_X1 i_0_1_488 (.A(n_0_1_241), .B1(n_0_1_256), .B2(n_0_1_810), .ZN(
      n_0_434));
   AOI222_X1 i_0_1_489 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[17]), .C1(n_0_1_255), .C2(A_imm_2s_complement[17]), 
      .ZN(n_0_1_241));
   OAI21_X1 i_0_1_490 (.A(n_0_1_242), .B1(n_0_1_256), .B2(n_0_1_812), .ZN(
      n_0_435));
   AOI222_X1 i_0_1_491 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[18]), .C1(n_0_1_255), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_242));
   OAI21_X1 i_0_1_492 (.A(n_0_1_243), .B1(n_0_1_256), .B2(n_0_1_814), .ZN(
      n_0_436));
   AOI222_X1 i_0_1_493 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[19]), .C1(n_0_1_255), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_243));
   OAI21_X1 i_0_1_494 (.A(n_0_1_244), .B1(n_0_1_256), .B2(n_0_1_816), .ZN(
      n_0_437));
   AOI222_X1 i_0_1_495 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[20]), .C1(n_0_1_255), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_244));
   OAI21_X1 i_0_1_496 (.A(n_0_1_245), .B1(n_0_1_256), .B2(n_0_1_818), .ZN(
      n_0_438));
   AOI222_X1 i_0_1_497 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[21]), .C1(n_0_1_255), .C2(A_imm_2s_complement[21]), 
      .ZN(n_0_1_245));
   OAI21_X1 i_0_1_498 (.A(n_0_1_246), .B1(n_0_1_256), .B2(n_0_1_820), .ZN(
      n_0_439));
   AOI222_X1 i_0_1_499 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[22]), .C1(n_0_1_255), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_246));
   OAI21_X1 i_0_1_500 (.A(n_0_1_247), .B1(n_0_1_256), .B2(n_0_1_822), .ZN(
      n_0_440));
   AOI222_X1 i_0_1_501 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[23]), .C1(n_0_1_255), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_247));
   OAI21_X1 i_0_1_502 (.A(n_0_1_248), .B1(n_0_1_256), .B2(n_0_1_824), .ZN(
      n_0_441));
   AOI222_X1 i_0_1_503 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[24]), .C1(n_0_1_255), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_248));
   OAI21_X1 i_0_1_504 (.A(n_0_1_249), .B1(n_0_1_256), .B2(n_0_1_826), .ZN(
      n_0_442));
   AOI222_X1 i_0_1_505 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[25]), .C1(n_0_1_255), .C2(A_imm_2s_complement[25]), 
      .ZN(n_0_1_249));
   OAI21_X1 i_0_1_506 (.A(n_0_1_250), .B1(n_0_1_256), .B2(n_0_1_828), .ZN(
      n_0_443));
   AOI222_X1 i_0_1_507 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[26]), .C1(n_0_1_255), .C2(A_imm_2s_complement[26]), 
      .ZN(n_0_1_250));
   OAI21_X1 i_0_1_508 (.A(n_0_1_251), .B1(n_0_1_256), .B2(n_0_1_830), .ZN(
      n_0_444));
   AOI222_X1 i_0_1_509 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[27]), .C1(n_0_1_255), .C2(A_imm_2s_complement[27]), 
      .ZN(n_0_1_251));
   OAI21_X1 i_0_1_510 (.A(n_0_1_252), .B1(n_0_1_256), .B2(n_0_1_832), .ZN(
      n_0_445));
   AOI222_X1 i_0_1_511 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[28]), .C1(n_0_1_255), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_252));
   OAI21_X1 i_0_1_512 (.A(n_0_1_253), .B1(n_0_1_256), .B2(n_0_1_834), .ZN(
      n_0_446));
   AOI222_X1 i_0_1_513 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[29]), .C1(n_0_1_255), .C2(A_imm_2s_complement[29]), 
      .ZN(n_0_1_253));
   OAI21_X1 i_0_1_514 (.A(n_0_1_254), .B1(n_0_1_256), .B2(n_0_1_836), .ZN(
      n_0_447));
   AOI222_X1 i_0_1_515 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_258), .B1(
      n_0_1_257), .B2(A_imm[30]), .C1(n_0_1_255), .C2(A_imm_2s_complement[30]), 
      .ZN(n_0_1_254));
   NOR3_X1 i_0_1_516 (.A1(n_0_1_262), .A2(n_0_1_265), .A3(n_0_1_306), .ZN(
      n_0_1_255));
   NAND2_X1 i_0_1_517 (.A1(n_0_1_259), .A2(n_0_1_262), .ZN(n_0_1_256));
   NOR2_X1 i_0_1_518 (.A1(n_0_1_264), .A2(n_0_1_263), .ZN(n_0_1_257));
   AND2_X1 i_0_1_519 (.A1(n_0_1_263), .A2(n_0_1_259), .ZN(n_0_1_258));
   XNOR2_X1 i_0_1_520 (.A(n_0_1_305), .B(n_0_1_265), .ZN(n_0_1_259));
   OAI21_X1 i_0_1_521 (.A(n_0_1_261), .B1(n_0_1_260), .B2(n_0_1_263), .ZN(
      n_0_448));
   OAI21_X1 i_0_1_522 (.A(A_imm[31]), .B1(n_0_1_306), .B2(n_0_1_265), .ZN(
      n_0_1_260));
   NAND3_X1 i_0_1_523 (.A1(n_0_1_264), .A2(n_0_1_263), .A3(
      A_imm_2s_complement[31]), .ZN(n_0_1_261));
   INV_X1 i_0_1_524 (.A(n_0_1_263), .ZN(n_0_1_262));
   MUX2_X1 i_0_1_525 (.A(n_0_161), .B(n_0_55), .S(B_in), .Z(n_0_1_263));
   NAND2_X1 i_0_1_526 (.A1(n_0_1_306), .A2(n_0_1_265), .ZN(n_0_1_264));
   MUX2_X1 i_0_1_527 (.A(n_0_162), .B(n_0_54), .S(B_in), .Z(n_0_1_265));
   AND2_X1 i_0_1_528 (.A1(n_0_1_302), .A2(n_0_155), .ZN(n_0_449));
   OAI211_X1 i_0_1_529 (.A(n_0_1_267), .B(n_0_1_266), .C1(n_0_1_776), .C2(
      n_0_1_299), .ZN(n_0_450));
   OAI21_X1 i_0_1_530 (.A(n_0_155), .B1(n_0_1_300), .B2(n_0_1_298), .ZN(
      n_0_1_266));
   NAND2_X1 i_0_1_531 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_301), .ZN(
      n_0_1_267));
   OAI21_X1 i_0_1_532 (.A(n_0_1_268), .B1(n_0_1_299), .B2(n_0_1_778), .ZN(
      n_0_451));
   AOI222_X1 i_0_1_533 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[1]), .C1(n_0_1_298), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_268));
   OAI21_X1 i_0_1_534 (.A(n_0_1_269), .B1(n_0_1_299), .B2(n_0_1_780), .ZN(
      n_0_452));
   AOI222_X1 i_0_1_535 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[2]), .C1(n_0_1_298), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_269));
   OAI21_X1 i_0_1_536 (.A(n_0_1_270), .B1(n_0_1_299), .B2(n_0_1_782), .ZN(
      n_0_453));
   AOI222_X1 i_0_1_537 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[3]), .C1(n_0_1_298), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_270));
   OAI21_X1 i_0_1_538 (.A(n_0_1_271), .B1(n_0_1_299), .B2(n_0_1_784), .ZN(
      n_0_454));
   AOI222_X1 i_0_1_539 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[4]), .C1(n_0_1_298), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_271));
   OAI21_X1 i_0_1_540 (.A(n_0_1_272), .B1(n_0_1_299), .B2(n_0_1_786), .ZN(
      n_0_455));
   AOI222_X1 i_0_1_541 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[5]), .C1(n_0_1_298), .C2(A_imm_2s_complement[5]), 
      .ZN(n_0_1_272));
   OAI21_X1 i_0_1_542 (.A(n_0_1_273), .B1(n_0_1_299), .B2(n_0_1_788), .ZN(
      n_0_456));
   AOI222_X1 i_0_1_543 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[6]), .C1(n_0_1_298), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_273));
   OAI21_X1 i_0_1_544 (.A(n_0_1_274), .B1(n_0_1_299), .B2(n_0_1_790), .ZN(
      n_0_457));
   AOI222_X1 i_0_1_545 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[7]), .C1(n_0_1_298), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_274));
   OAI21_X1 i_0_1_546 (.A(n_0_1_275), .B1(n_0_1_299), .B2(n_0_1_792), .ZN(
      n_0_458));
   AOI222_X1 i_0_1_547 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[8]), .C1(n_0_1_298), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_275));
   OAI21_X1 i_0_1_548 (.A(n_0_1_276), .B1(n_0_1_299), .B2(n_0_1_794), .ZN(
      n_0_459));
   AOI222_X1 i_0_1_549 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[9]), .C1(n_0_1_298), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_276));
   OAI21_X1 i_0_1_550 (.A(n_0_1_277), .B1(n_0_1_299), .B2(n_0_1_796), .ZN(
      n_0_460));
   AOI222_X1 i_0_1_551 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[10]), .C1(n_0_1_298), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_277));
   OAI21_X1 i_0_1_552 (.A(n_0_1_278), .B1(n_0_1_299), .B2(n_0_1_798), .ZN(
      n_0_461));
   AOI222_X1 i_0_1_553 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[11]), .C1(n_0_1_298), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_278));
   OAI21_X1 i_0_1_554 (.A(n_0_1_279), .B1(n_0_1_299), .B2(n_0_1_800), .ZN(
      n_0_462));
   AOI222_X1 i_0_1_555 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[12]), .C1(n_0_1_298), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_279));
   OAI21_X1 i_0_1_556 (.A(n_0_1_280), .B1(n_0_1_299), .B2(n_0_1_802), .ZN(
      n_0_463));
   AOI222_X1 i_0_1_557 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[13]), .C1(n_0_1_298), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_280));
   OAI21_X1 i_0_1_558 (.A(n_0_1_281), .B1(n_0_1_299), .B2(n_0_1_804), .ZN(
      n_0_464));
   AOI222_X1 i_0_1_559 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[14]), .C1(n_0_1_298), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_281));
   OAI21_X1 i_0_1_560 (.A(n_0_1_282), .B1(n_0_1_299), .B2(n_0_1_806), .ZN(
      n_0_465));
   AOI222_X1 i_0_1_561 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[15]), .C1(n_0_1_298), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_282));
   OAI21_X1 i_0_1_562 (.A(n_0_1_283), .B1(n_0_1_299), .B2(n_0_1_808), .ZN(
      n_0_466));
   AOI222_X1 i_0_1_563 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[16]), .C1(n_0_1_298), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_283));
   OAI21_X1 i_0_1_564 (.A(n_0_1_284), .B1(n_0_1_299), .B2(n_0_1_810), .ZN(
      n_0_467));
   AOI222_X1 i_0_1_565 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[17]), .C1(n_0_1_298), .C2(A_imm_2s_complement[17]), 
      .ZN(n_0_1_284));
   OAI21_X1 i_0_1_566 (.A(n_0_1_285), .B1(n_0_1_299), .B2(n_0_1_812), .ZN(
      n_0_468));
   AOI222_X1 i_0_1_567 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[18]), .C1(n_0_1_298), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_285));
   OAI21_X1 i_0_1_568 (.A(n_0_1_286), .B1(n_0_1_299), .B2(n_0_1_814), .ZN(
      n_0_469));
   AOI222_X1 i_0_1_569 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[19]), .C1(n_0_1_298), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_286));
   OAI21_X1 i_0_1_570 (.A(n_0_1_287), .B1(n_0_1_299), .B2(n_0_1_816), .ZN(
      n_0_470));
   AOI222_X1 i_0_1_571 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[20]), .C1(n_0_1_298), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_287));
   OAI21_X1 i_0_1_572 (.A(n_0_1_288), .B1(n_0_1_299), .B2(n_0_1_818), .ZN(
      n_0_471));
   AOI222_X1 i_0_1_573 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[21]), .C1(n_0_1_298), .C2(A_imm_2s_complement[21]), 
      .ZN(n_0_1_288));
   OAI21_X1 i_0_1_574 (.A(n_0_1_289), .B1(n_0_1_299), .B2(n_0_1_820), .ZN(
      n_0_472));
   AOI222_X1 i_0_1_575 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[22]), .C1(n_0_1_298), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_289));
   OAI21_X1 i_0_1_576 (.A(n_0_1_290), .B1(n_0_1_299), .B2(n_0_1_822), .ZN(
      n_0_473));
   AOI222_X1 i_0_1_577 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[23]), .C1(n_0_1_298), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_290));
   OAI21_X1 i_0_1_578 (.A(n_0_1_291), .B1(n_0_1_299), .B2(n_0_1_824), .ZN(
      n_0_474));
   AOI222_X1 i_0_1_579 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[24]), .C1(n_0_1_298), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_291));
   OAI21_X1 i_0_1_580 (.A(n_0_1_292), .B1(n_0_1_299), .B2(n_0_1_826), .ZN(
      n_0_475));
   AOI222_X1 i_0_1_581 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[25]), .C1(n_0_1_298), .C2(A_imm_2s_complement[25]), 
      .ZN(n_0_1_292));
   OAI21_X1 i_0_1_582 (.A(n_0_1_293), .B1(n_0_1_299), .B2(n_0_1_828), .ZN(
      n_0_476));
   AOI222_X1 i_0_1_583 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[26]), .C1(n_0_1_298), .C2(A_imm_2s_complement[26]), 
      .ZN(n_0_1_293));
   OAI21_X1 i_0_1_584 (.A(n_0_1_294), .B1(n_0_1_299), .B2(n_0_1_830), .ZN(
      n_0_477));
   AOI222_X1 i_0_1_585 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[27]), .C1(n_0_1_298), .C2(A_imm_2s_complement[27]), 
      .ZN(n_0_1_294));
   OAI21_X1 i_0_1_586 (.A(n_0_1_295), .B1(n_0_1_299), .B2(n_0_1_832), .ZN(
      n_0_478));
   AOI222_X1 i_0_1_587 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[28]), .C1(n_0_1_298), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_295));
   OAI21_X1 i_0_1_588 (.A(n_0_1_296), .B1(n_0_1_299), .B2(n_0_1_834), .ZN(
      n_0_479));
   AOI222_X1 i_0_1_589 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[29]), .C1(n_0_1_298), .C2(A_imm_2s_complement[29]), 
      .ZN(n_0_1_296));
   OAI21_X1 i_0_1_590 (.A(n_0_1_297), .B1(n_0_1_299), .B2(n_0_1_836), .ZN(
      n_0_480));
   AOI222_X1 i_0_1_591 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_301), .B1(
      n_0_1_300), .B2(A_imm[30]), .C1(n_0_1_298), .C2(A_imm_2s_complement[30]), 
      .ZN(n_0_1_297));
   NOR3_X1 i_0_1_592 (.A1(n_0_1_305), .A2(n_0_1_308), .A3(n_0_1_349), .ZN(
      n_0_1_298));
   NAND2_X1 i_0_1_593 (.A1(n_0_1_302), .A2(n_0_1_305), .ZN(n_0_1_299));
   NOR2_X1 i_0_1_594 (.A1(n_0_1_307), .A2(n_0_1_306), .ZN(n_0_1_300));
   AND2_X1 i_0_1_595 (.A1(n_0_1_306), .A2(n_0_1_302), .ZN(n_0_1_301));
   XNOR2_X1 i_0_1_596 (.A(n_0_1_348), .B(n_0_1_308), .ZN(n_0_1_302));
   OAI21_X1 i_0_1_597 (.A(n_0_1_304), .B1(n_0_1_303), .B2(n_0_1_306), .ZN(
      n_0_481));
   OAI21_X1 i_0_1_598 (.A(A_imm[31]), .B1(n_0_1_349), .B2(n_0_1_308), .ZN(
      n_0_1_303));
   NAND3_X1 i_0_1_599 (.A1(n_0_1_307), .A2(n_0_1_306), .A3(
      A_imm_2s_complement[31]), .ZN(n_0_1_304));
   INV_X1 i_0_1_600 (.A(n_0_1_306), .ZN(n_0_1_305));
   MUX2_X1 i_0_1_601 (.A(n_0_163), .B(n_0_53), .S(B_in), .Z(n_0_1_306));
   NAND2_X1 i_0_1_602 (.A1(n_0_1_349), .A2(n_0_1_308), .ZN(n_0_1_307));
   MUX2_X1 i_0_1_603 (.A(n_0_164), .B(n_0_52), .S(B_in), .Z(n_0_1_308));
   AND2_X1 i_0_1_604 (.A1(n_0_1_345), .A2(n_0_155), .ZN(n_0_482));
   OAI211_X1 i_0_1_605 (.A(n_0_1_310), .B(n_0_1_309), .C1(n_0_1_776), .C2(
      n_0_1_342), .ZN(n_0_483));
   OAI21_X1 i_0_1_606 (.A(n_0_155), .B1(n_0_1_343), .B2(n_0_1_341), .ZN(
      n_0_1_309));
   NAND2_X1 i_0_1_607 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_344), .ZN(
      n_0_1_310));
   OAI21_X1 i_0_1_608 (.A(n_0_1_311), .B1(n_0_1_342), .B2(n_0_1_778), .ZN(
      n_0_484));
   AOI222_X1 i_0_1_609 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[1]), .C1(n_0_1_341), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_311));
   OAI21_X1 i_0_1_610 (.A(n_0_1_312), .B1(n_0_1_342), .B2(n_0_1_780), .ZN(
      n_0_485));
   AOI222_X1 i_0_1_611 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[2]), .C1(n_0_1_341), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_312));
   OAI21_X1 i_0_1_612 (.A(n_0_1_313), .B1(n_0_1_342), .B2(n_0_1_782), .ZN(
      n_0_486));
   AOI222_X1 i_0_1_613 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[3]), .C1(n_0_1_341), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_313));
   OAI21_X1 i_0_1_614 (.A(n_0_1_314), .B1(n_0_1_342), .B2(n_0_1_784), .ZN(
      n_0_487));
   AOI222_X1 i_0_1_615 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[4]), .C1(n_0_1_341), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_314));
   OAI21_X1 i_0_1_616 (.A(n_0_1_315), .B1(n_0_1_342), .B2(n_0_1_786), .ZN(
      n_0_488));
   AOI222_X1 i_0_1_617 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[5]), .C1(n_0_1_341), .C2(A_imm_2s_complement[5]), 
      .ZN(n_0_1_315));
   OAI21_X1 i_0_1_618 (.A(n_0_1_316), .B1(n_0_1_342), .B2(n_0_1_788), .ZN(
      n_0_489));
   AOI222_X1 i_0_1_619 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[6]), .C1(n_0_1_341), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_316));
   OAI21_X1 i_0_1_620 (.A(n_0_1_317), .B1(n_0_1_342), .B2(n_0_1_790), .ZN(
      n_0_490));
   AOI222_X1 i_0_1_621 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[7]), .C1(n_0_1_341), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_317));
   OAI21_X1 i_0_1_622 (.A(n_0_1_318), .B1(n_0_1_342), .B2(n_0_1_792), .ZN(
      n_0_491));
   AOI222_X1 i_0_1_623 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[8]), .C1(n_0_1_341), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_318));
   OAI21_X1 i_0_1_624 (.A(n_0_1_319), .B1(n_0_1_342), .B2(n_0_1_794), .ZN(
      n_0_492));
   AOI222_X1 i_0_1_625 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[9]), .C1(n_0_1_341), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_319));
   OAI21_X1 i_0_1_626 (.A(n_0_1_320), .B1(n_0_1_342), .B2(n_0_1_796), .ZN(
      n_0_493));
   AOI222_X1 i_0_1_627 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[10]), .C1(n_0_1_341), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_320));
   OAI21_X1 i_0_1_628 (.A(n_0_1_321), .B1(n_0_1_342), .B2(n_0_1_798), .ZN(
      n_0_494));
   AOI222_X1 i_0_1_629 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[11]), .C1(n_0_1_341), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_321));
   OAI21_X1 i_0_1_630 (.A(n_0_1_322), .B1(n_0_1_342), .B2(n_0_1_800), .ZN(
      n_0_495));
   AOI222_X1 i_0_1_631 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[12]), .C1(n_0_1_341), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_322));
   OAI21_X1 i_0_1_632 (.A(n_0_1_323), .B1(n_0_1_342), .B2(n_0_1_802), .ZN(
      n_0_496));
   AOI222_X1 i_0_1_633 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[13]), .C1(n_0_1_341), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_323));
   OAI21_X1 i_0_1_634 (.A(n_0_1_324), .B1(n_0_1_342), .B2(n_0_1_804), .ZN(
      n_0_497));
   AOI222_X1 i_0_1_635 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[14]), .C1(n_0_1_341), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_324));
   OAI21_X1 i_0_1_636 (.A(n_0_1_325), .B1(n_0_1_342), .B2(n_0_1_806), .ZN(
      n_0_498));
   AOI222_X1 i_0_1_637 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[15]), .C1(n_0_1_341), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_325));
   OAI21_X1 i_0_1_638 (.A(n_0_1_326), .B1(n_0_1_342), .B2(n_0_1_808), .ZN(
      n_0_499));
   AOI222_X1 i_0_1_639 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[16]), .C1(n_0_1_341), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_326));
   OAI21_X1 i_0_1_640 (.A(n_0_1_327), .B1(n_0_1_342), .B2(n_0_1_810), .ZN(
      n_0_500));
   AOI222_X1 i_0_1_641 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[17]), .C1(n_0_1_341), .C2(A_imm_2s_complement[17]), 
      .ZN(n_0_1_327));
   OAI21_X1 i_0_1_642 (.A(n_0_1_328), .B1(n_0_1_342), .B2(n_0_1_812), .ZN(
      n_0_501));
   AOI222_X1 i_0_1_643 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[18]), .C1(n_0_1_341), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_328));
   OAI21_X1 i_0_1_644 (.A(n_0_1_329), .B1(n_0_1_342), .B2(n_0_1_814), .ZN(
      n_0_502));
   AOI222_X1 i_0_1_645 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[19]), .C1(n_0_1_341), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_329));
   OAI21_X1 i_0_1_646 (.A(n_0_1_330), .B1(n_0_1_342), .B2(n_0_1_816), .ZN(
      n_0_503));
   AOI222_X1 i_0_1_647 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[20]), .C1(n_0_1_341), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_330));
   OAI21_X1 i_0_1_648 (.A(n_0_1_331), .B1(n_0_1_342), .B2(n_0_1_818), .ZN(
      n_0_504));
   AOI222_X1 i_0_1_649 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[21]), .C1(n_0_1_341), .C2(A_imm_2s_complement[21]), 
      .ZN(n_0_1_331));
   OAI21_X1 i_0_1_650 (.A(n_0_1_332), .B1(n_0_1_342), .B2(n_0_1_820), .ZN(
      n_0_505));
   AOI222_X1 i_0_1_651 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[22]), .C1(n_0_1_341), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_332));
   OAI21_X1 i_0_1_652 (.A(n_0_1_333), .B1(n_0_1_342), .B2(n_0_1_822), .ZN(
      n_0_506));
   AOI222_X1 i_0_1_653 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[23]), .C1(n_0_1_341), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_333));
   OAI21_X1 i_0_1_654 (.A(n_0_1_334), .B1(n_0_1_342), .B2(n_0_1_824), .ZN(
      n_0_507));
   AOI222_X1 i_0_1_655 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[24]), .C1(n_0_1_341), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_334));
   OAI21_X1 i_0_1_656 (.A(n_0_1_335), .B1(n_0_1_342), .B2(n_0_1_826), .ZN(
      n_0_508));
   AOI222_X1 i_0_1_657 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[25]), .C1(n_0_1_341), .C2(A_imm_2s_complement[25]), 
      .ZN(n_0_1_335));
   OAI21_X1 i_0_1_658 (.A(n_0_1_336), .B1(n_0_1_342), .B2(n_0_1_828), .ZN(
      n_0_509));
   AOI222_X1 i_0_1_659 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[26]), .C1(n_0_1_341), .C2(A_imm_2s_complement[26]), 
      .ZN(n_0_1_336));
   OAI21_X1 i_0_1_660 (.A(n_0_1_337), .B1(n_0_1_342), .B2(n_0_1_830), .ZN(
      n_0_510));
   AOI222_X1 i_0_1_661 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[27]), .C1(n_0_1_341), .C2(A_imm_2s_complement[27]), 
      .ZN(n_0_1_337));
   OAI21_X1 i_0_1_662 (.A(n_0_1_338), .B1(n_0_1_342), .B2(n_0_1_832), .ZN(
      n_0_511));
   AOI222_X1 i_0_1_663 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[28]), .C1(n_0_1_341), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_338));
   OAI21_X1 i_0_1_664 (.A(n_0_1_339), .B1(n_0_1_342), .B2(n_0_1_834), .ZN(
      n_0_512));
   AOI222_X1 i_0_1_665 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[29]), .C1(n_0_1_341), .C2(A_imm_2s_complement[29]), 
      .ZN(n_0_1_339));
   OAI21_X1 i_0_1_666 (.A(n_0_1_340), .B1(n_0_1_342), .B2(n_0_1_836), .ZN(
      n_0_513));
   AOI222_X1 i_0_1_667 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_344), .B1(
      n_0_1_343), .B2(A_imm[30]), .C1(n_0_1_341), .C2(A_imm_2s_complement[30]), 
      .ZN(n_0_1_340));
   NOR3_X1 i_0_1_668 (.A1(n_0_1_348), .A2(n_0_1_351), .A3(n_0_1_394), .ZN(
      n_0_1_341));
   NAND2_X1 i_0_1_669 (.A1(n_0_1_345), .A2(n_0_1_348), .ZN(n_0_1_342));
   NOR2_X1 i_0_1_670 (.A1(n_0_1_349), .A2(n_0_1_347), .ZN(n_0_1_343));
   AND2_X1 i_0_1_671 (.A1(n_0_1_349), .A2(n_0_1_345), .ZN(n_0_1_344));
   XNOR2_X1 i_0_1_672 (.A(n_0_1_393), .B(n_0_1_351), .ZN(n_0_1_345));
   OAI21_X1 i_0_1_673 (.A(n_0_1_346), .B1(n_0_1_349), .B2(n_0_1_350), .ZN(
      n_0_514));
   NAND3_X1 i_0_1_674 (.A1(n_0_1_347), .A2(A_imm_2s_complement[31]), .A3(
      n_0_1_349), .ZN(n_0_1_346));
   NAND2_X1 i_0_1_675 (.A1(n_0_1_394), .A2(n_0_1_351), .ZN(n_0_1_347));
   INV_X1 i_0_1_676 (.A(n_0_1_349), .ZN(n_0_1_348));
   MUX2_X1 i_0_1_677 (.A(n_0_165), .B(n_0_51), .S(B_in), .Z(n_0_1_349));
   OAI21_X1 i_0_1_678 (.A(A_imm[31]), .B1(n_0_1_394), .B2(n_0_1_351), .ZN(
      n_0_1_350));
   MUX2_X1 i_0_1_679 (.A(n_0_166), .B(n_0_50), .S(B_in), .Z(n_0_1_351));
   AND2_X1 i_0_1_680 (.A1(n_0_1_388), .A2(n_0_155), .ZN(n_0_515));
   OAI211_X1 i_0_1_681 (.A(n_0_1_353), .B(n_0_1_352), .C1(n_0_1_776), .C2(
      n_0_1_385), .ZN(n_0_516));
   OAI21_X1 i_0_1_682 (.A(n_0_155), .B1(n_0_1_386), .B2(n_0_1_384), .ZN(
      n_0_1_352));
   NAND2_X1 i_0_1_683 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_387), .ZN(
      n_0_1_353));
   OAI21_X1 i_0_1_684 (.A(n_0_1_354), .B1(n_0_1_385), .B2(n_0_1_778), .ZN(
      n_0_517));
   AOI222_X1 i_0_1_685 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[1]), .C1(n_0_1_384), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_354));
   OAI21_X1 i_0_1_686 (.A(n_0_1_355), .B1(n_0_1_385), .B2(n_0_1_780), .ZN(
      n_0_518));
   AOI222_X1 i_0_1_687 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[2]), .C1(n_0_1_384), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_355));
   OAI21_X1 i_0_1_688 (.A(n_0_1_356), .B1(n_0_1_385), .B2(n_0_1_782), .ZN(
      n_0_519));
   AOI222_X1 i_0_1_689 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[3]), .C1(n_0_1_384), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_356));
   OAI21_X1 i_0_1_690 (.A(n_0_1_357), .B1(n_0_1_385), .B2(n_0_1_784), .ZN(
      n_0_520));
   AOI222_X1 i_0_1_691 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[4]), .C1(n_0_1_384), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_357));
   OAI21_X1 i_0_1_692 (.A(n_0_1_358), .B1(n_0_1_385), .B2(n_0_1_786), .ZN(
      n_0_521));
   AOI222_X1 i_0_1_693 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[5]), .C1(n_0_1_384), .C2(A_imm_2s_complement[5]), 
      .ZN(n_0_1_358));
   OAI21_X1 i_0_1_694 (.A(n_0_1_359), .B1(n_0_1_385), .B2(n_0_1_788), .ZN(
      n_0_522));
   AOI222_X1 i_0_1_695 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[6]), .C1(n_0_1_384), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_359));
   OAI21_X1 i_0_1_696 (.A(n_0_1_360), .B1(n_0_1_385), .B2(n_0_1_790), .ZN(
      n_0_523));
   AOI222_X1 i_0_1_697 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[7]), .C1(n_0_1_384), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_360));
   OAI21_X1 i_0_1_698 (.A(n_0_1_361), .B1(n_0_1_385), .B2(n_0_1_792), .ZN(
      n_0_524));
   AOI222_X1 i_0_1_699 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[8]), .C1(n_0_1_384), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_361));
   OAI21_X1 i_0_1_700 (.A(n_0_1_362), .B1(n_0_1_385), .B2(n_0_1_794), .ZN(
      n_0_525));
   AOI222_X1 i_0_1_701 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[9]), .C1(n_0_1_384), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_362));
   OAI21_X1 i_0_1_702 (.A(n_0_1_363), .B1(n_0_1_385), .B2(n_0_1_796), .ZN(
      n_0_526));
   AOI222_X1 i_0_1_703 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[10]), .C1(n_0_1_384), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_363));
   OAI21_X1 i_0_1_704 (.A(n_0_1_364), .B1(n_0_1_385), .B2(n_0_1_798), .ZN(
      n_0_527));
   AOI222_X1 i_0_1_705 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[11]), .C1(n_0_1_384), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_364));
   OAI21_X1 i_0_1_706 (.A(n_0_1_365), .B1(n_0_1_385), .B2(n_0_1_800), .ZN(
      n_0_528));
   AOI222_X1 i_0_1_707 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[12]), .C1(n_0_1_384), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_365));
   OAI21_X1 i_0_1_708 (.A(n_0_1_366), .B1(n_0_1_385), .B2(n_0_1_802), .ZN(
      n_0_529));
   AOI222_X1 i_0_1_709 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[13]), .C1(n_0_1_384), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_366));
   OAI21_X1 i_0_1_710 (.A(n_0_1_367), .B1(n_0_1_385), .B2(n_0_1_804), .ZN(
      n_0_530));
   AOI222_X1 i_0_1_711 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[14]), .C1(n_0_1_384), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_367));
   OAI21_X1 i_0_1_712 (.A(n_0_1_368), .B1(n_0_1_385), .B2(n_0_1_806), .ZN(
      n_0_531));
   AOI222_X1 i_0_1_713 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[15]), .C1(n_0_1_384), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_368));
   OAI21_X1 i_0_1_714 (.A(n_0_1_369), .B1(n_0_1_385), .B2(n_0_1_808), .ZN(
      n_0_532));
   AOI222_X1 i_0_1_715 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[16]), .C1(n_0_1_384), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_369));
   OAI21_X1 i_0_1_716 (.A(n_0_1_370), .B1(n_0_1_385), .B2(n_0_1_810), .ZN(
      n_0_533));
   AOI222_X1 i_0_1_717 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[17]), .C1(n_0_1_384), .C2(A_imm_2s_complement[17]), 
      .ZN(n_0_1_370));
   OAI21_X1 i_0_1_718 (.A(n_0_1_371), .B1(n_0_1_385), .B2(n_0_1_812), .ZN(
      n_0_534));
   AOI222_X1 i_0_1_719 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[18]), .C1(n_0_1_384), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_371));
   OAI21_X1 i_0_1_720 (.A(n_0_1_372), .B1(n_0_1_385), .B2(n_0_1_814), .ZN(
      n_0_535));
   AOI222_X1 i_0_1_721 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[19]), .C1(n_0_1_384), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_372));
   OAI21_X1 i_0_1_722 (.A(n_0_1_373), .B1(n_0_1_385), .B2(n_0_1_816), .ZN(
      n_0_536));
   AOI222_X1 i_0_1_723 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[20]), .C1(n_0_1_384), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_373));
   OAI21_X1 i_0_1_724 (.A(n_0_1_374), .B1(n_0_1_385), .B2(n_0_1_818), .ZN(
      n_0_537));
   AOI222_X1 i_0_1_725 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[21]), .C1(n_0_1_384), .C2(A_imm_2s_complement[21]), 
      .ZN(n_0_1_374));
   OAI21_X1 i_0_1_726 (.A(n_0_1_375), .B1(n_0_1_385), .B2(n_0_1_820), .ZN(
      n_0_538));
   AOI222_X1 i_0_1_727 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[22]), .C1(n_0_1_384), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_375));
   OAI21_X1 i_0_1_728 (.A(n_0_1_376), .B1(n_0_1_385), .B2(n_0_1_822), .ZN(
      n_0_539));
   AOI222_X1 i_0_1_729 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[23]), .C1(n_0_1_384), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_376));
   OAI21_X1 i_0_1_730 (.A(n_0_1_377), .B1(n_0_1_385), .B2(n_0_1_824), .ZN(
      n_0_540));
   AOI222_X1 i_0_1_731 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[24]), .C1(n_0_1_384), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_377));
   OAI21_X1 i_0_1_732 (.A(n_0_1_378), .B1(n_0_1_385), .B2(n_0_1_826), .ZN(
      n_0_541));
   AOI222_X1 i_0_1_733 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[25]), .C1(n_0_1_384), .C2(A_imm_2s_complement[25]), 
      .ZN(n_0_1_378));
   OAI21_X1 i_0_1_734 (.A(n_0_1_379), .B1(n_0_1_385), .B2(n_0_1_828), .ZN(
      n_0_542));
   AOI222_X1 i_0_1_735 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[26]), .C1(n_0_1_384), .C2(A_imm_2s_complement[26]), 
      .ZN(n_0_1_379));
   OAI21_X1 i_0_1_736 (.A(n_0_1_380), .B1(n_0_1_385), .B2(n_0_1_830), .ZN(
      n_0_543));
   AOI222_X1 i_0_1_737 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[27]), .C1(n_0_1_384), .C2(A_imm_2s_complement[27]), 
      .ZN(n_0_1_380));
   OAI21_X1 i_0_1_738 (.A(n_0_1_381), .B1(n_0_1_385), .B2(n_0_1_832), .ZN(
      n_0_544));
   AOI222_X1 i_0_1_739 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[28]), .C1(n_0_1_384), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_381));
   OAI21_X1 i_0_1_740 (.A(n_0_1_382), .B1(n_0_1_385), .B2(n_0_1_834), .ZN(
      n_0_545));
   AOI222_X1 i_0_1_741 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[29]), .C1(n_0_1_384), .C2(A_imm_2s_complement[29]), 
      .ZN(n_0_1_382));
   OAI21_X1 i_0_1_742 (.A(n_0_1_383), .B1(n_0_1_385), .B2(n_0_1_836), .ZN(
      n_0_546));
   AOI222_X1 i_0_1_743 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_387), .B1(
      n_0_1_386), .B2(A_imm[30]), .C1(n_0_1_384), .C2(A_imm_2s_complement[30]), 
      .ZN(n_0_1_383));
   NOR3_X1 i_0_1_744 (.A1(n_0_1_393), .A2(n_0_1_392), .A3(n_0_1_435), .ZN(
      n_0_1_384));
   NAND2_X1 i_0_1_745 (.A1(n_0_1_388), .A2(n_0_1_393), .ZN(n_0_1_385));
   NOR2_X1 i_0_1_746 (.A1(n_0_1_394), .A2(n_0_1_390), .ZN(n_0_1_386));
   AND2_X1 i_0_1_747 (.A1(n_0_1_394), .A2(n_0_1_388), .ZN(n_0_1_387));
   XNOR2_X1 i_0_1_748 (.A(n_0_1_434), .B(n_0_1_392), .ZN(n_0_1_388));
   OAI21_X1 i_0_1_749 (.A(n_0_1_389), .B1(n_0_1_391), .B2(n_0_1_394), .ZN(
      n_0_547));
   NAND3_X1 i_0_1_750 (.A1(n_0_1_390), .A2(A_imm_2s_complement[31]), .A3(
      n_0_1_394), .ZN(n_0_1_389));
   NAND2_X1 i_0_1_751 (.A1(n_0_1_435), .A2(n_0_1_392), .ZN(n_0_1_390));
   OAI21_X1 i_0_1_752 (.A(A_imm[31]), .B1(n_0_1_435), .B2(n_0_1_392), .ZN(
      n_0_1_391));
   MUX2_X1 i_0_1_753 (.A(n_0_168), .B(n_0_48), .S(B_in), .Z(n_0_1_392));
   INV_X1 i_0_1_754 (.A(n_0_1_394), .ZN(n_0_1_393));
   MUX2_X1 i_0_1_755 (.A(n_0_167), .B(n_0_49), .S(B_in), .Z(n_0_1_394));
   AND2_X1 i_0_1_756 (.A1(n_0_1_431), .A2(n_0_155), .ZN(n_0_548));
   OAI211_X1 i_0_1_757 (.A(n_0_1_396), .B(n_0_1_395), .C1(n_0_1_776), .C2(
      n_0_1_428), .ZN(n_0_549));
   OAI21_X1 i_0_1_758 (.A(n_0_155), .B1(n_0_1_429), .B2(n_0_1_427), .ZN(
      n_0_1_395));
   NAND2_X1 i_0_1_759 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_430), .ZN(
      n_0_1_396));
   OAI21_X1 i_0_1_760 (.A(n_0_1_397), .B1(n_0_1_428), .B2(n_0_1_778), .ZN(
      n_0_550));
   AOI222_X1 i_0_1_761 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[1]), .C1(n_0_1_427), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_397));
   OAI21_X1 i_0_1_762 (.A(n_0_1_398), .B1(n_0_1_428), .B2(n_0_1_780), .ZN(
      n_0_551));
   AOI222_X1 i_0_1_763 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[2]), .C1(n_0_1_427), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_398));
   OAI21_X1 i_0_1_764 (.A(n_0_1_399), .B1(n_0_1_428), .B2(n_0_1_782), .ZN(
      n_0_552));
   AOI222_X1 i_0_1_765 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[3]), .C1(n_0_1_427), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_399));
   OAI21_X1 i_0_1_766 (.A(n_0_1_400), .B1(n_0_1_428), .B2(n_0_1_784), .ZN(
      n_0_553));
   AOI222_X1 i_0_1_767 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[4]), .C1(n_0_1_427), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_400));
   OAI21_X1 i_0_1_768 (.A(n_0_1_401), .B1(n_0_1_428), .B2(n_0_1_786), .ZN(
      n_0_554));
   AOI222_X1 i_0_1_769 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[5]), .C1(n_0_1_427), .C2(A_imm_2s_complement[5]), 
      .ZN(n_0_1_401));
   OAI21_X1 i_0_1_770 (.A(n_0_1_402), .B1(n_0_1_428), .B2(n_0_1_788), .ZN(
      n_0_555));
   AOI222_X1 i_0_1_771 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[6]), .C1(n_0_1_427), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_402));
   OAI21_X1 i_0_1_772 (.A(n_0_1_403), .B1(n_0_1_428), .B2(n_0_1_790), .ZN(
      n_0_556));
   AOI222_X1 i_0_1_773 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[7]), .C1(n_0_1_427), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_403));
   OAI21_X1 i_0_1_774 (.A(n_0_1_404), .B1(n_0_1_428), .B2(n_0_1_792), .ZN(
      n_0_557));
   AOI222_X1 i_0_1_775 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[8]), .C1(n_0_1_427), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_404));
   OAI21_X1 i_0_1_776 (.A(n_0_1_405), .B1(n_0_1_428), .B2(n_0_1_794), .ZN(
      n_0_558));
   AOI222_X1 i_0_1_777 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[9]), .C1(n_0_1_427), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_405));
   OAI21_X1 i_0_1_778 (.A(n_0_1_406), .B1(n_0_1_428), .B2(n_0_1_796), .ZN(
      n_0_559));
   AOI222_X1 i_0_1_779 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[10]), .C1(n_0_1_427), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_406));
   OAI21_X1 i_0_1_780 (.A(n_0_1_407), .B1(n_0_1_428), .B2(n_0_1_798), .ZN(
      n_0_560));
   AOI222_X1 i_0_1_781 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[11]), .C1(n_0_1_427), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_407));
   OAI21_X1 i_0_1_782 (.A(n_0_1_408), .B1(n_0_1_428), .B2(n_0_1_800), .ZN(
      n_0_561));
   AOI222_X1 i_0_1_783 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[12]), .C1(n_0_1_427), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_408));
   OAI21_X1 i_0_1_784 (.A(n_0_1_409), .B1(n_0_1_428), .B2(n_0_1_802), .ZN(
      n_0_562));
   AOI222_X1 i_0_1_785 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[13]), .C1(n_0_1_427), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_409));
   OAI21_X1 i_0_1_786 (.A(n_0_1_410), .B1(n_0_1_428), .B2(n_0_1_804), .ZN(
      n_0_563));
   AOI222_X1 i_0_1_787 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[14]), .C1(n_0_1_427), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_410));
   OAI21_X1 i_0_1_788 (.A(n_0_1_411), .B1(n_0_1_428), .B2(n_0_1_806), .ZN(
      n_0_564));
   AOI222_X1 i_0_1_789 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[15]), .C1(n_0_1_427), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_411));
   OAI21_X1 i_0_1_790 (.A(n_0_1_412), .B1(n_0_1_428), .B2(n_0_1_808), .ZN(
      n_0_565));
   AOI222_X1 i_0_1_791 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[16]), .C1(n_0_1_427), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_412));
   OAI21_X1 i_0_1_792 (.A(n_0_1_413), .B1(n_0_1_428), .B2(n_0_1_810), .ZN(
      n_0_566));
   AOI222_X1 i_0_1_793 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[17]), .C1(n_0_1_427), .C2(A_imm_2s_complement[17]), 
      .ZN(n_0_1_413));
   OAI21_X1 i_0_1_794 (.A(n_0_1_414), .B1(n_0_1_428), .B2(n_0_1_812), .ZN(
      n_0_567));
   AOI222_X1 i_0_1_795 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[18]), .C1(n_0_1_427), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_414));
   OAI21_X1 i_0_1_796 (.A(n_0_1_415), .B1(n_0_1_428), .B2(n_0_1_814), .ZN(
      n_0_568));
   AOI222_X1 i_0_1_797 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[19]), .C1(n_0_1_427), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_415));
   OAI21_X1 i_0_1_798 (.A(n_0_1_416), .B1(n_0_1_428), .B2(n_0_1_816), .ZN(
      n_0_569));
   AOI222_X1 i_0_1_799 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[20]), .C1(n_0_1_427), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_416));
   OAI21_X1 i_0_1_800 (.A(n_0_1_417), .B1(n_0_1_428), .B2(n_0_1_818), .ZN(
      n_0_570));
   AOI222_X1 i_0_1_801 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[21]), .C1(n_0_1_427), .C2(A_imm_2s_complement[21]), 
      .ZN(n_0_1_417));
   OAI21_X1 i_0_1_802 (.A(n_0_1_418), .B1(n_0_1_428), .B2(n_0_1_820), .ZN(
      n_0_571));
   AOI222_X1 i_0_1_803 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[22]), .C1(n_0_1_427), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_418));
   OAI21_X1 i_0_1_804 (.A(n_0_1_419), .B1(n_0_1_428), .B2(n_0_1_822), .ZN(
      n_0_572));
   AOI222_X1 i_0_1_805 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[23]), .C1(n_0_1_427), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_419));
   OAI21_X1 i_0_1_806 (.A(n_0_1_420), .B1(n_0_1_428), .B2(n_0_1_824), .ZN(
      n_0_573));
   AOI222_X1 i_0_1_807 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[24]), .C1(n_0_1_427), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_420));
   OAI21_X1 i_0_1_808 (.A(n_0_1_421), .B1(n_0_1_428), .B2(n_0_1_826), .ZN(
      n_0_574));
   AOI222_X1 i_0_1_809 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[25]), .C1(n_0_1_427), .C2(A_imm_2s_complement[25]), 
      .ZN(n_0_1_421));
   OAI21_X1 i_0_1_810 (.A(n_0_1_422), .B1(n_0_1_428), .B2(n_0_1_828), .ZN(
      n_0_575));
   AOI222_X1 i_0_1_811 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[26]), .C1(n_0_1_427), .C2(A_imm_2s_complement[26]), 
      .ZN(n_0_1_422));
   OAI21_X1 i_0_1_812 (.A(n_0_1_423), .B1(n_0_1_428), .B2(n_0_1_830), .ZN(
      n_0_576));
   AOI222_X1 i_0_1_813 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[27]), .C1(n_0_1_427), .C2(A_imm_2s_complement[27]), 
      .ZN(n_0_1_423));
   OAI21_X1 i_0_1_814 (.A(n_0_1_424), .B1(n_0_1_428), .B2(n_0_1_832), .ZN(
      n_0_577));
   AOI222_X1 i_0_1_815 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[28]), .C1(n_0_1_427), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_424));
   OAI21_X1 i_0_1_816 (.A(n_0_1_425), .B1(n_0_1_428), .B2(n_0_1_834), .ZN(
      n_0_578));
   AOI222_X1 i_0_1_817 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[29]), .C1(n_0_1_427), .C2(A_imm_2s_complement[29]), 
      .ZN(n_0_1_425));
   OAI21_X1 i_0_1_818 (.A(n_0_1_426), .B1(n_0_1_428), .B2(n_0_1_836), .ZN(
      n_0_579));
   AOI222_X1 i_0_1_819 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_430), .B1(
      n_0_1_429), .B2(A_imm[30]), .C1(n_0_1_427), .C2(A_imm_2s_complement[30]), 
      .ZN(n_0_1_426));
   NOR3_X1 i_0_1_820 (.A1(n_0_1_434), .A2(n_0_1_437), .A3(n_0_1_478), .ZN(
      n_0_1_427));
   NAND2_X1 i_0_1_821 (.A1(n_0_1_431), .A2(n_0_1_434), .ZN(n_0_1_428));
   NOR2_X1 i_0_1_822 (.A1(n_0_1_436), .A2(n_0_1_435), .ZN(n_0_1_429));
   AND2_X1 i_0_1_823 (.A1(n_0_1_435), .A2(n_0_1_431), .ZN(n_0_1_430));
   XNOR2_X1 i_0_1_824 (.A(n_0_1_477), .B(n_0_1_437), .ZN(n_0_1_431));
   OAI21_X1 i_0_1_825 (.A(n_0_1_433), .B1(n_0_1_432), .B2(n_0_1_435), .ZN(
      n_0_580));
   OAI21_X1 i_0_1_826 (.A(A_imm[31]), .B1(n_0_1_478), .B2(n_0_1_437), .ZN(
      n_0_1_432));
   NAND3_X1 i_0_1_827 (.A1(n_0_1_436), .A2(n_0_1_435), .A3(
      A_imm_2s_complement[31]), .ZN(n_0_1_433));
   INV_X1 i_0_1_828 (.A(n_0_1_435), .ZN(n_0_1_434));
   MUX2_X1 i_0_1_829 (.A(n_0_169), .B(n_0_47), .S(B_in), .Z(n_0_1_435));
   NAND2_X1 i_0_1_830 (.A1(n_0_1_478), .A2(n_0_1_437), .ZN(n_0_1_436));
   MUX2_X1 i_0_1_831 (.A(n_0_170), .B(n_0_46), .S(B_in), .Z(n_0_1_437));
   AND2_X1 i_0_1_832 (.A1(n_0_1_474), .A2(n_0_155), .ZN(n_0_581));
   OAI211_X1 i_0_1_833 (.A(n_0_1_439), .B(n_0_1_438), .C1(n_0_1_776), .C2(
      n_0_1_471), .ZN(n_0_582));
   OAI21_X1 i_0_1_834 (.A(n_0_155), .B1(n_0_1_472), .B2(n_0_1_470), .ZN(
      n_0_1_438));
   NAND2_X1 i_0_1_835 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_473), .ZN(
      n_0_1_439));
   OAI21_X1 i_0_1_836 (.A(n_0_1_440), .B1(n_0_1_471), .B2(n_0_1_778), .ZN(
      n_0_583));
   AOI222_X1 i_0_1_837 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[1]), .C1(n_0_1_470), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_440));
   OAI21_X1 i_0_1_838 (.A(n_0_1_441), .B1(n_0_1_471), .B2(n_0_1_780), .ZN(
      n_0_584));
   AOI222_X1 i_0_1_839 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[2]), .C1(n_0_1_470), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_441));
   OAI21_X1 i_0_1_840 (.A(n_0_1_442), .B1(n_0_1_471), .B2(n_0_1_782), .ZN(
      n_0_585));
   AOI222_X1 i_0_1_841 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[3]), .C1(n_0_1_470), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_442));
   OAI21_X1 i_0_1_842 (.A(n_0_1_443), .B1(n_0_1_471), .B2(n_0_1_784), .ZN(
      n_0_586));
   AOI222_X1 i_0_1_843 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[4]), .C1(n_0_1_470), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_443));
   OAI21_X1 i_0_1_844 (.A(n_0_1_444), .B1(n_0_1_471), .B2(n_0_1_786), .ZN(
      n_0_587));
   AOI222_X1 i_0_1_845 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[5]), .C1(n_0_1_470), .C2(A_imm_2s_complement[5]), 
      .ZN(n_0_1_444));
   OAI21_X1 i_0_1_846 (.A(n_0_1_445), .B1(n_0_1_471), .B2(n_0_1_788), .ZN(
      n_0_588));
   AOI222_X1 i_0_1_847 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[6]), .C1(n_0_1_470), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_445));
   OAI21_X1 i_0_1_848 (.A(n_0_1_446), .B1(n_0_1_471), .B2(n_0_1_790), .ZN(
      n_0_589));
   AOI222_X1 i_0_1_849 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[7]), .C1(n_0_1_470), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_446));
   OAI21_X1 i_0_1_850 (.A(n_0_1_447), .B1(n_0_1_471), .B2(n_0_1_792), .ZN(
      n_0_590));
   AOI222_X1 i_0_1_851 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[8]), .C1(n_0_1_470), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_447));
   OAI21_X1 i_0_1_852 (.A(n_0_1_448), .B1(n_0_1_471), .B2(n_0_1_794), .ZN(
      n_0_591));
   AOI222_X1 i_0_1_853 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[9]), .C1(n_0_1_470), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_448));
   OAI21_X1 i_0_1_854 (.A(n_0_1_449), .B1(n_0_1_471), .B2(n_0_1_796), .ZN(
      n_0_592));
   AOI222_X1 i_0_1_855 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[10]), .C1(n_0_1_470), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_449));
   OAI21_X1 i_0_1_856 (.A(n_0_1_450), .B1(n_0_1_471), .B2(n_0_1_798), .ZN(
      n_0_593));
   AOI222_X1 i_0_1_857 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[11]), .C1(n_0_1_470), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_450));
   OAI21_X1 i_0_1_858 (.A(n_0_1_451), .B1(n_0_1_471), .B2(n_0_1_800), .ZN(
      n_0_594));
   AOI222_X1 i_0_1_859 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[12]), .C1(n_0_1_470), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_451));
   OAI21_X1 i_0_1_860 (.A(n_0_1_452), .B1(n_0_1_471), .B2(n_0_1_802), .ZN(
      n_0_595));
   AOI222_X1 i_0_1_861 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[13]), .C1(n_0_1_470), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_452));
   OAI21_X1 i_0_1_862 (.A(n_0_1_453), .B1(n_0_1_471), .B2(n_0_1_804), .ZN(
      n_0_596));
   AOI222_X1 i_0_1_863 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[14]), .C1(n_0_1_470), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_453));
   OAI21_X1 i_0_1_864 (.A(n_0_1_454), .B1(n_0_1_471), .B2(n_0_1_806), .ZN(
      n_0_597));
   AOI222_X1 i_0_1_865 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[15]), .C1(n_0_1_470), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_454));
   OAI21_X1 i_0_1_866 (.A(n_0_1_455), .B1(n_0_1_471), .B2(n_0_1_808), .ZN(
      n_0_598));
   AOI222_X1 i_0_1_867 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[16]), .C1(n_0_1_470), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_455));
   OAI21_X1 i_0_1_868 (.A(n_0_1_456), .B1(n_0_1_471), .B2(n_0_1_810), .ZN(
      n_0_599));
   AOI222_X1 i_0_1_869 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[17]), .C1(n_0_1_470), .C2(A_imm_2s_complement[17]), 
      .ZN(n_0_1_456));
   OAI21_X1 i_0_1_870 (.A(n_0_1_457), .B1(n_0_1_471), .B2(n_0_1_812), .ZN(
      n_0_600));
   AOI222_X1 i_0_1_871 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[18]), .C1(n_0_1_470), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_457));
   OAI21_X1 i_0_1_872 (.A(n_0_1_458), .B1(n_0_1_471), .B2(n_0_1_814), .ZN(
      n_0_601));
   AOI222_X1 i_0_1_873 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[19]), .C1(n_0_1_470), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_458));
   OAI21_X1 i_0_1_874 (.A(n_0_1_459), .B1(n_0_1_471), .B2(n_0_1_816), .ZN(
      n_0_602));
   AOI222_X1 i_0_1_875 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[20]), .C1(n_0_1_470), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_459));
   OAI21_X1 i_0_1_876 (.A(n_0_1_460), .B1(n_0_1_471), .B2(n_0_1_818), .ZN(
      n_0_603));
   AOI222_X1 i_0_1_877 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[21]), .C1(n_0_1_470), .C2(A_imm_2s_complement[21]), 
      .ZN(n_0_1_460));
   OAI21_X1 i_0_1_878 (.A(n_0_1_461), .B1(n_0_1_471), .B2(n_0_1_820), .ZN(
      n_0_604));
   AOI222_X1 i_0_1_879 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[22]), .C1(n_0_1_470), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_461));
   OAI21_X1 i_0_1_880 (.A(n_0_1_462), .B1(n_0_1_471), .B2(n_0_1_822), .ZN(
      n_0_605));
   AOI222_X1 i_0_1_881 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[23]), .C1(n_0_1_470), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_462));
   OAI21_X1 i_0_1_882 (.A(n_0_1_463), .B1(n_0_1_471), .B2(n_0_1_824), .ZN(
      n_0_606));
   AOI222_X1 i_0_1_883 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[24]), .C1(n_0_1_470), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_463));
   OAI21_X1 i_0_1_884 (.A(n_0_1_464), .B1(n_0_1_471), .B2(n_0_1_826), .ZN(
      n_0_607));
   AOI222_X1 i_0_1_885 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[25]), .C1(n_0_1_470), .C2(A_imm_2s_complement[25]), 
      .ZN(n_0_1_464));
   OAI21_X1 i_0_1_886 (.A(n_0_1_465), .B1(n_0_1_471), .B2(n_0_1_828), .ZN(
      n_0_608));
   AOI222_X1 i_0_1_887 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[26]), .C1(n_0_1_470), .C2(A_imm_2s_complement[26]), 
      .ZN(n_0_1_465));
   OAI21_X1 i_0_1_888 (.A(n_0_1_466), .B1(n_0_1_471), .B2(n_0_1_830), .ZN(
      n_0_609));
   AOI222_X1 i_0_1_889 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[27]), .C1(n_0_1_470), .C2(A_imm_2s_complement[27]), 
      .ZN(n_0_1_466));
   OAI21_X1 i_0_1_890 (.A(n_0_1_467), .B1(n_0_1_471), .B2(n_0_1_832), .ZN(
      n_0_610));
   AOI222_X1 i_0_1_891 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[28]), .C1(n_0_1_470), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_467));
   OAI21_X1 i_0_1_892 (.A(n_0_1_468), .B1(n_0_1_471), .B2(n_0_1_834), .ZN(
      n_0_611));
   AOI222_X1 i_0_1_893 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[29]), .C1(n_0_1_470), .C2(A_imm_2s_complement[29]), 
      .ZN(n_0_1_468));
   OAI21_X1 i_0_1_894 (.A(n_0_1_469), .B1(n_0_1_471), .B2(n_0_1_836), .ZN(
      n_0_612));
   AOI222_X1 i_0_1_895 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_473), .B1(
      n_0_1_472), .B2(A_imm[30]), .C1(n_0_1_470), .C2(A_imm_2s_complement[30]), 
      .ZN(n_0_1_469));
   NOR3_X1 i_0_1_896 (.A1(n_0_1_477), .A2(n_0_1_480), .A3(n_0_1_523), .ZN(
      n_0_1_470));
   NAND2_X1 i_0_1_897 (.A1(n_0_1_474), .A2(n_0_1_477), .ZN(n_0_1_471));
   NOR2_X1 i_0_1_898 (.A1(n_0_1_479), .A2(n_0_1_478), .ZN(n_0_1_472));
   AND2_X1 i_0_1_899 (.A1(n_0_1_478), .A2(n_0_1_474), .ZN(n_0_1_473));
   XNOR2_X1 i_0_1_900 (.A(n_0_1_522), .B(n_0_1_480), .ZN(n_0_1_474));
   OAI21_X1 i_0_1_901 (.A(n_0_1_476), .B1(n_0_1_475), .B2(n_0_1_478), .ZN(
      n_0_613));
   OAI21_X1 i_0_1_902 (.A(A_imm[31]), .B1(n_0_1_523), .B2(n_0_1_480), .ZN(
      n_0_1_475));
   NAND3_X1 i_0_1_903 (.A1(n_0_1_479), .A2(n_0_1_478), .A3(
      A_imm_2s_complement[31]), .ZN(n_0_1_476));
   INV_X1 i_0_1_904 (.A(n_0_1_478), .ZN(n_0_1_477));
   MUX2_X1 i_0_1_905 (.A(n_0_171), .B(n_0_45), .S(B_in), .Z(n_0_1_478));
   NAND2_X1 i_0_1_906 (.A1(n_0_1_523), .A2(n_0_1_480), .ZN(n_0_1_479));
   MUX2_X1 i_0_1_907 (.A(n_0_172), .B(n_0_44), .S(B_in), .Z(n_0_1_480));
   AND2_X1 i_0_1_908 (.A1(n_0_1_517), .A2(n_0_155), .ZN(n_0_614));
   OAI211_X1 i_0_1_909 (.A(n_0_1_482), .B(n_0_1_481), .C1(n_0_1_776), .C2(
      n_0_1_514), .ZN(n_0_615));
   OAI21_X1 i_0_1_910 (.A(n_0_155), .B1(n_0_1_515), .B2(n_0_1_513), .ZN(
      n_0_1_481));
   NAND2_X1 i_0_1_911 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_516), .ZN(
      n_0_1_482));
   OAI21_X1 i_0_1_912 (.A(n_0_1_483), .B1(n_0_1_514), .B2(n_0_1_778), .ZN(
      n_0_616));
   AOI222_X1 i_0_1_913 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[1]), .C1(n_0_1_513), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_483));
   OAI21_X1 i_0_1_914 (.A(n_0_1_484), .B1(n_0_1_514), .B2(n_0_1_780), .ZN(
      n_0_617));
   AOI222_X1 i_0_1_915 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[2]), .C1(n_0_1_513), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_484));
   OAI21_X1 i_0_1_916 (.A(n_0_1_485), .B1(n_0_1_514), .B2(n_0_1_782), .ZN(
      n_0_618));
   AOI222_X1 i_0_1_917 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[3]), .C1(n_0_1_513), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_485));
   OAI21_X1 i_0_1_918 (.A(n_0_1_486), .B1(n_0_1_514), .B2(n_0_1_784), .ZN(
      n_0_619));
   AOI222_X1 i_0_1_919 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[4]), .C1(n_0_1_513), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_486));
   OAI21_X1 i_0_1_920 (.A(n_0_1_487), .B1(n_0_1_514), .B2(n_0_1_786), .ZN(
      n_0_620));
   AOI222_X1 i_0_1_921 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[5]), .C1(n_0_1_513), .C2(A_imm_2s_complement[5]), 
      .ZN(n_0_1_487));
   OAI21_X1 i_0_1_922 (.A(n_0_1_488), .B1(n_0_1_514), .B2(n_0_1_788), .ZN(
      n_0_621));
   AOI222_X1 i_0_1_923 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[6]), .C1(n_0_1_513), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_488));
   OAI21_X1 i_0_1_924 (.A(n_0_1_489), .B1(n_0_1_514), .B2(n_0_1_790), .ZN(
      n_0_622));
   AOI222_X1 i_0_1_925 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[7]), .C1(n_0_1_513), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_489));
   OAI21_X1 i_0_1_926 (.A(n_0_1_490), .B1(n_0_1_514), .B2(n_0_1_792), .ZN(
      n_0_623));
   AOI222_X1 i_0_1_927 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[8]), .C1(n_0_1_513), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_490));
   OAI21_X1 i_0_1_928 (.A(n_0_1_491), .B1(n_0_1_514), .B2(n_0_1_794), .ZN(
      n_0_624));
   AOI222_X1 i_0_1_929 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[9]), .C1(n_0_1_513), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_491));
   OAI21_X1 i_0_1_930 (.A(n_0_1_492), .B1(n_0_1_514), .B2(n_0_1_796), .ZN(
      n_0_625));
   AOI222_X1 i_0_1_931 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[10]), .C1(n_0_1_513), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_492));
   OAI21_X1 i_0_1_932 (.A(n_0_1_493), .B1(n_0_1_514), .B2(n_0_1_798), .ZN(
      n_0_626));
   AOI222_X1 i_0_1_933 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[11]), .C1(n_0_1_513), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_493));
   OAI21_X1 i_0_1_934 (.A(n_0_1_494), .B1(n_0_1_514), .B2(n_0_1_800), .ZN(
      n_0_627));
   AOI222_X1 i_0_1_935 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[12]), .C1(n_0_1_513), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_494));
   OAI21_X1 i_0_1_936 (.A(n_0_1_495), .B1(n_0_1_514), .B2(n_0_1_802), .ZN(
      n_0_628));
   AOI222_X1 i_0_1_937 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[13]), .C1(n_0_1_513), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_495));
   OAI21_X1 i_0_1_938 (.A(n_0_1_496), .B1(n_0_1_514), .B2(n_0_1_804), .ZN(
      n_0_629));
   AOI222_X1 i_0_1_939 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[14]), .C1(n_0_1_513), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_496));
   OAI21_X1 i_0_1_940 (.A(n_0_1_497), .B1(n_0_1_514), .B2(n_0_1_806), .ZN(
      n_0_630));
   AOI222_X1 i_0_1_941 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[15]), .C1(n_0_1_513), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_497));
   OAI21_X1 i_0_1_942 (.A(n_0_1_498), .B1(n_0_1_514), .B2(n_0_1_808), .ZN(
      n_0_631));
   AOI222_X1 i_0_1_943 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[16]), .C1(n_0_1_513), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_498));
   OAI21_X1 i_0_1_944 (.A(n_0_1_499), .B1(n_0_1_514), .B2(n_0_1_810), .ZN(
      n_0_632));
   AOI222_X1 i_0_1_945 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[17]), .C1(n_0_1_513), .C2(A_imm_2s_complement[17]), 
      .ZN(n_0_1_499));
   OAI21_X1 i_0_1_946 (.A(n_0_1_500), .B1(n_0_1_514), .B2(n_0_1_812), .ZN(
      n_0_633));
   AOI222_X1 i_0_1_947 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[18]), .C1(n_0_1_513), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_500));
   OAI21_X1 i_0_1_948 (.A(n_0_1_501), .B1(n_0_1_514), .B2(n_0_1_814), .ZN(
      n_0_634));
   AOI222_X1 i_0_1_949 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[19]), .C1(n_0_1_513), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_501));
   OAI21_X1 i_0_1_950 (.A(n_0_1_502), .B1(n_0_1_514), .B2(n_0_1_816), .ZN(
      n_0_635));
   AOI222_X1 i_0_1_951 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[20]), .C1(n_0_1_513), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_502));
   OAI21_X1 i_0_1_952 (.A(n_0_1_503), .B1(n_0_1_514), .B2(n_0_1_818), .ZN(
      n_0_636));
   AOI222_X1 i_0_1_953 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[21]), .C1(n_0_1_513), .C2(A_imm_2s_complement[21]), 
      .ZN(n_0_1_503));
   OAI21_X1 i_0_1_954 (.A(n_0_1_504), .B1(n_0_1_514), .B2(n_0_1_820), .ZN(
      n_0_637));
   AOI222_X1 i_0_1_955 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[22]), .C1(n_0_1_513), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_504));
   OAI21_X1 i_0_1_956 (.A(n_0_1_505), .B1(n_0_1_514), .B2(n_0_1_822), .ZN(
      n_0_638));
   AOI222_X1 i_0_1_957 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[23]), .C1(n_0_1_513), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_505));
   OAI21_X1 i_0_1_958 (.A(n_0_1_506), .B1(n_0_1_514), .B2(n_0_1_824), .ZN(
      n_0_639));
   AOI222_X1 i_0_1_959 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[24]), .C1(n_0_1_513), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_506));
   OAI21_X1 i_0_1_960 (.A(n_0_1_507), .B1(n_0_1_514), .B2(n_0_1_826), .ZN(
      n_0_640));
   AOI222_X1 i_0_1_961 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[25]), .C1(n_0_1_513), .C2(A_imm_2s_complement[25]), 
      .ZN(n_0_1_507));
   OAI21_X1 i_0_1_962 (.A(n_0_1_508), .B1(n_0_1_514), .B2(n_0_1_828), .ZN(
      n_0_641));
   AOI222_X1 i_0_1_963 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[26]), .C1(n_0_1_513), .C2(A_imm_2s_complement[26]), 
      .ZN(n_0_1_508));
   OAI21_X1 i_0_1_964 (.A(n_0_1_509), .B1(n_0_1_514), .B2(n_0_1_830), .ZN(
      n_0_642));
   AOI222_X1 i_0_1_965 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[27]), .C1(n_0_1_513), .C2(A_imm_2s_complement[27]), 
      .ZN(n_0_1_509));
   OAI21_X1 i_0_1_966 (.A(n_0_1_510), .B1(n_0_1_514), .B2(n_0_1_832), .ZN(
      n_0_643));
   AOI222_X1 i_0_1_967 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[28]), .C1(n_0_1_513), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_510));
   OAI21_X1 i_0_1_968 (.A(n_0_1_511), .B1(n_0_1_514), .B2(n_0_1_834), .ZN(
      n_0_644));
   AOI222_X1 i_0_1_969 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[29]), .C1(n_0_1_513), .C2(A_imm_2s_complement[29]), 
      .ZN(n_0_1_511));
   OAI21_X1 i_0_1_970 (.A(n_0_1_512), .B1(n_0_1_514), .B2(n_0_1_836), .ZN(
      n_0_645));
   AOI222_X1 i_0_1_971 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_516), .B1(
      n_0_1_515), .B2(A_imm[30]), .C1(n_0_1_513), .C2(A_imm_2s_complement[30]), 
      .ZN(n_0_1_512));
   NOR3_X1 i_0_1_972 (.A1(n_0_1_522), .A2(n_0_1_521), .A3(n_0_1_566), .ZN(
      n_0_1_513));
   NAND2_X1 i_0_1_973 (.A1(n_0_1_517), .A2(n_0_1_522), .ZN(n_0_1_514));
   NOR2_X1 i_0_1_974 (.A1(n_0_1_523), .A2(n_0_1_519), .ZN(n_0_1_515));
   AND2_X1 i_0_1_975 (.A1(n_0_1_523), .A2(n_0_1_517), .ZN(n_0_1_516));
   XNOR2_X1 i_0_1_976 (.A(n_0_1_565), .B(n_0_1_521), .ZN(n_0_1_517));
   OAI21_X1 i_0_1_977 (.A(n_0_1_518), .B1(n_0_1_520), .B2(n_0_1_523), .ZN(
      n_0_646));
   NAND3_X1 i_0_1_978 (.A1(n_0_1_519), .A2(A_imm_2s_complement[31]), .A3(
      n_0_1_523), .ZN(n_0_1_518));
   NAND2_X1 i_0_1_979 (.A1(n_0_1_566), .A2(n_0_1_521), .ZN(n_0_1_519));
   OAI21_X1 i_0_1_980 (.A(A_imm[31]), .B1(n_0_1_566), .B2(n_0_1_521), .ZN(
      n_0_1_520));
   MUX2_X1 i_0_1_981 (.A(n_0_174), .B(n_0_42), .S(B_in), .Z(n_0_1_521));
   INV_X1 i_0_1_982 (.A(n_0_1_523), .ZN(n_0_1_522));
   MUX2_X1 i_0_1_983 (.A(n_0_173), .B(n_0_43), .S(B_in), .Z(n_0_1_523));
   AND2_X1 i_0_1_984 (.A1(n_0_1_560), .A2(n_0_155), .ZN(n_0_647));
   OAI211_X1 i_0_1_985 (.A(n_0_1_525), .B(n_0_1_524), .C1(n_0_1_776), .C2(
      n_0_1_557), .ZN(n_0_648));
   OAI21_X1 i_0_1_986 (.A(n_0_155), .B1(n_0_1_558), .B2(n_0_1_556), .ZN(
      n_0_1_524));
   NAND2_X1 i_0_1_987 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_559), .ZN(
      n_0_1_525));
   OAI21_X1 i_0_1_988 (.A(n_0_1_526), .B1(n_0_1_557), .B2(n_0_1_778), .ZN(
      n_0_649));
   AOI222_X1 i_0_1_989 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[1]), .C1(n_0_1_556), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_526));
   OAI21_X1 i_0_1_990 (.A(n_0_1_527), .B1(n_0_1_557), .B2(n_0_1_780), .ZN(
      n_0_650));
   AOI222_X1 i_0_1_991 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[2]), .C1(n_0_1_556), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_527));
   OAI21_X1 i_0_1_992 (.A(n_0_1_528), .B1(n_0_1_557), .B2(n_0_1_782), .ZN(
      n_0_651));
   AOI222_X1 i_0_1_993 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[3]), .C1(n_0_1_556), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_528));
   OAI21_X1 i_0_1_994 (.A(n_0_1_529), .B1(n_0_1_557), .B2(n_0_1_784), .ZN(
      n_0_652));
   AOI222_X1 i_0_1_995 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[4]), .C1(n_0_1_556), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_529));
   OAI21_X1 i_0_1_996 (.A(n_0_1_530), .B1(n_0_1_557), .B2(n_0_1_786), .ZN(
      n_0_653));
   AOI222_X1 i_0_1_997 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[5]), .C1(n_0_1_556), .C2(A_imm_2s_complement[5]), 
      .ZN(n_0_1_530));
   OAI21_X1 i_0_1_998 (.A(n_0_1_531), .B1(n_0_1_557), .B2(n_0_1_788), .ZN(
      n_0_654));
   AOI222_X1 i_0_1_999 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[6]), .C1(n_0_1_556), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_531));
   OAI21_X1 i_0_1_1000 (.A(n_0_1_532), .B1(n_0_1_557), .B2(n_0_1_790), .ZN(
      n_0_655));
   AOI222_X1 i_0_1_1001 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[7]), .C1(n_0_1_556), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_532));
   OAI21_X1 i_0_1_1002 (.A(n_0_1_533), .B1(n_0_1_557), .B2(n_0_1_792), .ZN(
      n_0_656));
   AOI222_X1 i_0_1_1003 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[8]), .C1(n_0_1_556), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_533));
   OAI21_X1 i_0_1_1004 (.A(n_0_1_534), .B1(n_0_1_557), .B2(n_0_1_794), .ZN(
      n_0_657));
   AOI222_X1 i_0_1_1005 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[9]), .C1(n_0_1_556), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_534));
   OAI21_X1 i_0_1_1006 (.A(n_0_1_535), .B1(n_0_1_557), .B2(n_0_1_796), .ZN(
      n_0_658));
   AOI222_X1 i_0_1_1007 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[10]), .C1(n_0_1_556), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_535));
   OAI21_X1 i_0_1_1008 (.A(n_0_1_536), .B1(n_0_1_557), .B2(n_0_1_798), .ZN(
      n_0_659));
   AOI222_X1 i_0_1_1009 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[11]), .C1(n_0_1_556), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_536));
   OAI21_X1 i_0_1_1010 (.A(n_0_1_537), .B1(n_0_1_557), .B2(n_0_1_800), .ZN(
      n_0_660));
   AOI222_X1 i_0_1_1011 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[12]), .C1(n_0_1_556), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_537));
   OAI21_X1 i_0_1_1012 (.A(n_0_1_538), .B1(n_0_1_557), .B2(n_0_1_802), .ZN(
      n_0_661));
   AOI222_X1 i_0_1_1013 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[13]), .C1(n_0_1_556), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_538));
   OAI21_X1 i_0_1_1014 (.A(n_0_1_539), .B1(n_0_1_557), .B2(n_0_1_804), .ZN(
      n_0_662));
   AOI222_X1 i_0_1_1015 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[14]), .C1(n_0_1_556), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_539));
   OAI21_X1 i_0_1_1016 (.A(n_0_1_540), .B1(n_0_1_557), .B2(n_0_1_806), .ZN(
      n_0_663));
   AOI222_X1 i_0_1_1017 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[15]), .C1(n_0_1_556), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_540));
   OAI21_X1 i_0_1_1018 (.A(n_0_1_541), .B1(n_0_1_557), .B2(n_0_1_808), .ZN(
      n_0_664));
   AOI222_X1 i_0_1_1019 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[16]), .C1(n_0_1_556), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_541));
   OAI21_X1 i_0_1_1020 (.A(n_0_1_542), .B1(n_0_1_557), .B2(n_0_1_810), .ZN(
      n_0_665));
   AOI222_X1 i_0_1_1021 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[17]), .C1(n_0_1_556), .C2(A_imm_2s_complement[17]), 
      .ZN(n_0_1_542));
   OAI21_X1 i_0_1_1022 (.A(n_0_1_543), .B1(n_0_1_557), .B2(n_0_1_812), .ZN(
      n_0_666));
   AOI222_X1 i_0_1_1023 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[18]), .C1(n_0_1_556), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_543));
   OAI21_X1 i_0_1_1024 (.A(n_0_1_544), .B1(n_0_1_557), .B2(n_0_1_814), .ZN(
      n_0_667));
   AOI222_X1 i_0_1_1025 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[19]), .C1(n_0_1_556), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_544));
   OAI21_X1 i_0_1_1026 (.A(n_0_1_545), .B1(n_0_1_557), .B2(n_0_1_816), .ZN(
      n_0_668));
   AOI222_X1 i_0_1_1027 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[20]), .C1(n_0_1_556), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_545));
   OAI21_X1 i_0_1_1028 (.A(n_0_1_546), .B1(n_0_1_557), .B2(n_0_1_818), .ZN(
      n_0_669));
   AOI222_X1 i_0_1_1029 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[21]), .C1(n_0_1_556), .C2(A_imm_2s_complement[21]), 
      .ZN(n_0_1_546));
   OAI21_X1 i_0_1_1030 (.A(n_0_1_547), .B1(n_0_1_557), .B2(n_0_1_820), .ZN(
      n_0_670));
   AOI222_X1 i_0_1_1031 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[22]), .C1(n_0_1_556), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_547));
   OAI21_X1 i_0_1_1032 (.A(n_0_1_548), .B1(n_0_1_557), .B2(n_0_1_822), .ZN(
      n_0_671));
   AOI222_X1 i_0_1_1033 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[23]), .C1(n_0_1_556), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_548));
   OAI21_X1 i_0_1_1034 (.A(n_0_1_549), .B1(n_0_1_557), .B2(n_0_1_824), .ZN(
      n_0_672));
   AOI222_X1 i_0_1_1035 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[24]), .C1(n_0_1_556), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_549));
   OAI21_X1 i_0_1_1036 (.A(n_0_1_550), .B1(n_0_1_557), .B2(n_0_1_826), .ZN(
      n_0_673));
   AOI222_X1 i_0_1_1037 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[25]), .C1(n_0_1_556), .C2(A_imm_2s_complement[25]), 
      .ZN(n_0_1_550));
   OAI21_X1 i_0_1_1038 (.A(n_0_1_551), .B1(n_0_1_557), .B2(n_0_1_828), .ZN(
      n_0_674));
   AOI222_X1 i_0_1_1039 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[26]), .C1(n_0_1_556), .C2(A_imm_2s_complement[26]), 
      .ZN(n_0_1_551));
   OAI21_X1 i_0_1_1040 (.A(n_0_1_552), .B1(n_0_1_557), .B2(n_0_1_830), .ZN(
      n_0_675));
   AOI222_X1 i_0_1_1041 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[27]), .C1(n_0_1_556), .C2(A_imm_2s_complement[27]), 
      .ZN(n_0_1_552));
   OAI21_X1 i_0_1_1042 (.A(n_0_1_553), .B1(n_0_1_557), .B2(n_0_1_832), .ZN(
      n_0_676));
   AOI222_X1 i_0_1_1043 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_559), .B1(
      n_0_1_558), .B2(A_imm[28]), .C1(n_0_1_556), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_553));
   XNOR2_X1 i_0_1_1052 (.A(n_0_1_606), .B(n_0_1_564), .ZN(n_0_1_560));
   OAI21_X1 i_0_1_1053 (.A(n_0_1_561), .B1(n_0_1_563), .B2(n_0_1_566), .ZN(
      n_0_679));
   NAND3_X1 i_0_1_1054 (.A1(n_0_1_562), .A2(A_imm_2s_complement[31]), .A3(
      n_0_1_566), .ZN(n_0_1_561));
   NAND2_X1 i_0_1_1055 (.A1(n_0_1_607), .A2(n_0_1_564), .ZN(n_0_1_562));
   OAI21_X1 i_0_1_1056 (.A(A_imm[31]), .B1(n_0_1_607), .B2(n_0_1_564), .ZN(
      n_0_1_563));
   MUX2_X1 i_0_1_1057 (.A(n_0_176), .B(n_0_40), .S(B_in), .Z(n_0_1_564));
   INV_X1 i_0_1_1058 (.A(n_0_1_566), .ZN(n_0_1_565));
   MUX2_X1 i_0_1_1059 (.A(n_0_175), .B(n_0_41), .S(B_in), .Z(n_0_1_566));
   AND2_X1 i_0_1_1060 (.A1(n_0_1_603), .A2(n_0_155), .ZN(n_0_680));
   OAI211_X1 i_0_1_1061 (.A(n_0_1_568), .B(n_0_1_567), .C1(n_0_1_776), .C2(
      n_0_1_600), .ZN(n_0_681));
   OAI21_X1 i_0_1_1062 (.A(n_0_155), .B1(n_0_1_601), .B2(n_0_1_599), .ZN(
      n_0_1_567));
   NAND2_X1 i_0_1_1063 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_602), .ZN(
      n_0_1_568));
   OAI21_X1 i_0_1_1064 (.A(n_0_1_569), .B1(n_0_1_600), .B2(n_0_1_778), .ZN(
      n_0_682));
   AOI222_X1 i_0_1_1065 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[1]), .C1(n_0_1_599), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_569));
   OAI21_X1 i_0_1_1066 (.A(n_0_1_570), .B1(n_0_1_600), .B2(n_0_1_780), .ZN(
      n_0_683));
   AOI222_X1 i_0_1_1067 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[2]), .C1(n_0_1_599), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_570));
   OAI21_X1 i_0_1_1068 (.A(n_0_1_571), .B1(n_0_1_600), .B2(n_0_1_782), .ZN(
      n_0_684));
   AOI222_X1 i_0_1_1069 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[3]), .C1(n_0_1_599), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_571));
   OAI21_X1 i_0_1_1070 (.A(n_0_1_572), .B1(n_0_1_600), .B2(n_0_1_784), .ZN(
      n_0_685));
   AOI222_X1 i_0_1_1071 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[4]), .C1(n_0_1_599), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_572));
   OAI21_X1 i_0_1_1072 (.A(n_0_1_573), .B1(n_0_1_600), .B2(n_0_1_786), .ZN(
      n_0_686));
   AOI222_X1 i_0_1_1073 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[5]), .C1(n_0_1_599), .C2(A_imm_2s_complement[5]), 
      .ZN(n_0_1_573));
   OAI21_X1 i_0_1_1074 (.A(n_0_1_574), .B1(n_0_1_600), .B2(n_0_1_788), .ZN(
      n_0_687));
   AOI222_X1 i_0_1_1075 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[6]), .C1(n_0_1_599), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_574));
   OAI21_X1 i_0_1_1076 (.A(n_0_1_575), .B1(n_0_1_600), .B2(n_0_1_790), .ZN(
      n_0_688));
   AOI222_X1 i_0_1_1077 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[7]), .C1(n_0_1_599), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_575));
   OAI21_X1 i_0_1_1078 (.A(n_0_1_576), .B1(n_0_1_600), .B2(n_0_1_792), .ZN(
      n_0_689));
   AOI222_X1 i_0_1_1079 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[8]), .C1(n_0_1_599), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_576));
   OAI21_X1 i_0_1_1080 (.A(n_0_1_577), .B1(n_0_1_600), .B2(n_0_1_794), .ZN(
      n_0_690));
   AOI222_X1 i_0_1_1081 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[9]), .C1(n_0_1_599), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_577));
   OAI21_X1 i_0_1_1082 (.A(n_0_1_578), .B1(n_0_1_600), .B2(n_0_1_796), .ZN(
      n_0_691));
   AOI222_X1 i_0_1_1083 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[10]), .C1(n_0_1_599), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_578));
   OAI21_X1 i_0_1_1084 (.A(n_0_1_579), .B1(n_0_1_600), .B2(n_0_1_798), .ZN(
      n_0_692));
   AOI222_X1 i_0_1_1085 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[11]), .C1(n_0_1_599), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_579));
   OAI21_X1 i_0_1_1086 (.A(n_0_1_580), .B1(n_0_1_600), .B2(n_0_1_800), .ZN(
      n_0_693));
   AOI222_X1 i_0_1_1087 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[12]), .C1(n_0_1_599), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_580));
   OAI21_X1 i_0_1_1088 (.A(n_0_1_581), .B1(n_0_1_600), .B2(n_0_1_802), .ZN(
      n_0_694));
   AOI222_X1 i_0_1_1089 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[13]), .C1(n_0_1_599), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_581));
   OAI21_X1 i_0_1_1090 (.A(n_0_1_582), .B1(n_0_1_600), .B2(n_0_1_804), .ZN(
      n_0_695));
   AOI222_X1 i_0_1_1091 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[14]), .C1(n_0_1_599), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_582));
   OAI21_X1 i_0_1_1092 (.A(n_0_1_583), .B1(n_0_1_600), .B2(n_0_1_806), .ZN(
      n_0_696));
   AOI222_X1 i_0_1_1093 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[15]), .C1(n_0_1_599), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_583));
   OAI21_X1 i_0_1_1094 (.A(n_0_1_584), .B1(n_0_1_600), .B2(n_0_1_808), .ZN(
      n_0_697));
   AOI222_X1 i_0_1_1095 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[16]), .C1(n_0_1_599), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_584));
   OAI21_X1 i_0_1_1096 (.A(n_0_1_585), .B1(n_0_1_600), .B2(n_0_1_810), .ZN(
      n_0_698));
   AOI222_X1 i_0_1_1097 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[17]), .C1(n_0_1_599), .C2(A_imm_2s_complement[17]), 
      .ZN(n_0_1_585));
   OAI21_X1 i_0_1_1098 (.A(n_0_1_586), .B1(n_0_1_600), .B2(n_0_1_812), .ZN(
      n_0_699));
   AOI222_X1 i_0_1_1099 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[18]), .C1(n_0_1_599), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_586));
   OAI21_X1 i_0_1_1100 (.A(n_0_1_587), .B1(n_0_1_600), .B2(n_0_1_814), .ZN(
      n_0_700));
   AOI222_X1 i_0_1_1101 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[19]), .C1(n_0_1_599), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_587));
   OAI21_X1 i_0_1_1102 (.A(n_0_1_588), .B1(n_0_1_600), .B2(n_0_1_816), .ZN(
      n_0_701));
   AOI222_X1 i_0_1_1103 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[20]), .C1(n_0_1_599), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_588));
   OAI21_X1 i_0_1_1106 (.A(n_0_1_590), .B1(n_0_1_600), .B2(n_0_1_820), .ZN(
      n_0_703));
   AOI222_X1 i_0_1_1107 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[22]), .C1(n_0_1_599), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_590));
   OAI21_X1 i_0_1_1108 (.A(n_0_1_591), .B1(n_0_1_600), .B2(n_0_1_822), .ZN(
      n_0_704));
   AOI222_X1 i_0_1_1109 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[23]), .C1(n_0_1_599), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_591));
   OAI21_X1 i_0_1_1110 (.A(n_0_1_592), .B1(n_0_1_600), .B2(n_0_1_824), .ZN(
      n_0_705));
   AOI222_X1 i_0_1_1111 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[24]), .C1(n_0_1_599), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_592));
   OAI21_X1 i_0_1_1112 (.A(n_0_1_593), .B1(n_0_1_600), .B2(n_0_1_826), .ZN(
      n_0_706));
   AOI222_X1 i_0_1_1113 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[25]), .C1(n_0_1_599), .C2(A_imm_2s_complement[25]), 
      .ZN(n_0_1_593));
   OAI21_X1 i_0_1_1114 (.A(n_0_1_594), .B1(n_0_1_600), .B2(n_0_1_828), .ZN(
      n_0_707));
   AOI222_X1 i_0_1_1115 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[26]), .C1(n_0_1_599), .C2(A_imm_2s_complement[26]), 
      .ZN(n_0_1_594));
   OAI21_X1 i_0_1_1116 (.A(n_0_1_595), .B1(n_0_1_600), .B2(n_0_1_830), .ZN(
      n_0_708));
   AOI222_X1 i_0_1_1117 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[27]), .C1(n_0_1_599), .C2(A_imm_2s_complement[27]), 
      .ZN(n_0_1_595));
   OAI21_X1 i_0_1_1118 (.A(n_0_1_596), .B1(n_0_1_600), .B2(n_0_1_832), .ZN(
      n_0_709));
   AOI222_X1 i_0_1_1119 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[28]), .C1(n_0_1_599), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_596));
   OAI21_X1 i_0_1_1122 (.A(n_0_1_598), .B1(n_0_1_600), .B2(n_0_1_836), .ZN(
      n_0_711));
   AOI222_X1 i_0_1_1123 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_602), .B1(
      n_0_1_601), .B2(A_imm[30]), .C1(n_0_1_599), .C2(A_imm_2s_complement[30]), 
      .ZN(n_0_1_598));
   XNOR2_X1 i_0_1_1128 (.A(n_0_1_651), .B(n_0_1_609), .ZN(n_0_1_603));
   OAI21_X1 i_0_1_1129 (.A(n_0_1_605), .B1(n_0_1_604), .B2(n_0_1_607), .ZN(
      n_0_712));
   OAI21_X1 i_0_1_1130 (.A(A_imm[31]), .B1(n_0_1_652), .B2(n_0_1_609), .ZN(
      n_0_1_604));
   NAND3_X1 i_0_1_1131 (.A1(n_0_1_608), .A2(n_0_1_607), .A3(
      A_imm_2s_complement[31]), .ZN(n_0_1_605));
   INV_X1 i_0_1_1132 (.A(n_0_1_607), .ZN(n_0_1_606));
   MUX2_X1 i_0_1_1133 (.A(n_0_177), .B(n_0_39), .S(B_in), .Z(n_0_1_607));
   NAND2_X1 i_0_1_1134 (.A1(n_0_1_652), .A2(n_0_1_609), .ZN(n_0_1_608));
   MUX2_X1 i_0_1_1135 (.A(n_0_178), .B(n_0_38), .S(B_in), .Z(n_0_1_609));
   AND2_X1 i_0_1_1136 (.A1(n_0_1_646), .A2(n_0_155), .ZN(n_0_713));
   OAI211_X1 i_0_1_1137 (.A(n_0_1_611), .B(n_0_1_610), .C1(n_0_1_776), .C2(
      n_0_1_643), .ZN(n_0_714));
   OAI21_X1 i_0_1_1138 (.A(n_0_155), .B1(n_0_1_644), .B2(n_0_1_642), .ZN(
      n_0_1_610));
   NAND2_X1 i_0_1_1139 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_645), .ZN(
      n_0_1_611));
   OAI21_X1 i_0_1_1140 (.A(n_0_1_612), .B1(n_0_1_643), .B2(n_0_1_778), .ZN(
      n_0_715));
   AOI222_X1 i_0_1_1141 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[1]), .C1(n_0_1_642), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_612));
   OAI21_X1 i_0_1_1142 (.A(n_0_1_613), .B1(n_0_1_643), .B2(n_0_1_780), .ZN(
      n_0_716));
   AOI222_X1 i_0_1_1143 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[2]), .C1(n_0_1_642), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_613));
   OAI21_X1 i_0_1_1144 (.A(n_0_1_614), .B1(n_0_1_643), .B2(n_0_1_782), .ZN(
      n_0_717));
   AOI222_X1 i_0_1_1145 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[3]), .C1(n_0_1_642), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_614));
   OAI21_X1 i_0_1_1146 (.A(n_0_1_615), .B1(n_0_1_643), .B2(n_0_1_784), .ZN(
      n_0_718));
   AOI222_X1 i_0_1_1147 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[4]), .C1(n_0_1_642), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_615));
   OAI21_X1 i_0_1_1148 (.A(n_0_1_616), .B1(n_0_1_643), .B2(n_0_1_786), .ZN(
      n_0_719));
   AOI222_X1 i_0_1_1149 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[5]), .C1(n_0_1_642), .C2(A_imm_2s_complement[5]), 
      .ZN(n_0_1_616));
   OAI21_X1 i_0_1_1150 (.A(n_0_1_617), .B1(n_0_1_643), .B2(n_0_1_788), .ZN(
      n_0_720));
   AOI222_X1 i_0_1_1151 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[6]), .C1(n_0_1_642), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_617));
   OAI21_X1 i_0_1_1152 (.A(n_0_1_618), .B1(n_0_1_643), .B2(n_0_1_790), .ZN(
      n_0_721));
   AOI222_X1 i_0_1_1153 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[7]), .C1(n_0_1_642), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_618));
   OAI21_X1 i_0_1_1154 (.A(n_0_1_619), .B1(n_0_1_643), .B2(n_0_1_792), .ZN(
      n_0_722));
   AOI222_X1 i_0_1_1155 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[8]), .C1(n_0_1_642), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_619));
   OAI21_X1 i_0_1_1156 (.A(n_0_1_620), .B1(n_0_1_643), .B2(n_0_1_794), .ZN(
      n_0_723));
   AOI222_X1 i_0_1_1157 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[9]), .C1(n_0_1_642), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_620));
   OAI21_X1 i_0_1_1158 (.A(n_0_1_621), .B1(n_0_1_643), .B2(n_0_1_796), .ZN(
      n_0_724));
   AOI222_X1 i_0_1_1159 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[10]), .C1(n_0_1_642), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_621));
   OAI21_X1 i_0_1_1160 (.A(n_0_1_622), .B1(n_0_1_643), .B2(n_0_1_798), .ZN(
      n_0_725));
   AOI222_X1 i_0_1_1161 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[11]), .C1(n_0_1_642), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_622));
   OAI21_X1 i_0_1_1162 (.A(n_0_1_623), .B1(n_0_1_643), .B2(n_0_1_800), .ZN(
      n_0_726));
   AOI222_X1 i_0_1_1163 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[12]), .C1(n_0_1_642), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_623));
   OAI21_X1 i_0_1_1164 (.A(n_0_1_624), .B1(n_0_1_643), .B2(n_0_1_802), .ZN(
      n_0_727));
   AOI222_X1 i_0_1_1165 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[13]), .C1(n_0_1_642), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_624));
   OAI21_X1 i_0_1_1166 (.A(n_0_1_625), .B1(n_0_1_643), .B2(n_0_1_804), .ZN(
      n_0_728));
   AOI222_X1 i_0_1_1167 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[14]), .C1(n_0_1_642), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_625));
   OAI21_X1 i_0_1_1168 (.A(n_0_1_626), .B1(n_0_1_643), .B2(n_0_1_806), .ZN(
      n_0_729));
   AOI222_X1 i_0_1_1169 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[15]), .C1(n_0_1_642), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_626));
   OAI21_X1 i_0_1_1170 (.A(n_0_1_627), .B1(n_0_1_643), .B2(n_0_1_808), .ZN(
      n_0_730));
   AOI222_X1 i_0_1_1171 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[16]), .C1(n_0_1_642), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_627));
   OAI21_X1 i_0_1_1172 (.A(n_0_1_628), .B1(n_0_1_643), .B2(n_0_1_810), .ZN(
      n_0_731));
   AOI222_X1 i_0_1_1173 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[17]), .C1(n_0_1_642), .C2(A_imm_2s_complement[17]), 
      .ZN(n_0_1_628));
   OAI21_X1 i_0_1_1174 (.A(n_0_1_629), .B1(n_0_1_643), .B2(n_0_1_812), .ZN(
      n_0_732));
   AOI222_X1 i_0_1_1175 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[18]), .C1(n_0_1_642), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_629));
   OAI21_X1 i_0_1_1176 (.A(n_0_1_630), .B1(n_0_1_643), .B2(n_0_1_814), .ZN(
      n_0_733));
   AOI222_X1 i_0_1_1177 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[19]), .C1(n_0_1_642), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_630));
   OAI21_X1 i_0_1_1178 (.A(n_0_1_631), .B1(n_0_1_643), .B2(n_0_1_816), .ZN(
      n_0_734));
   AOI222_X1 i_0_1_1179 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[20]), .C1(n_0_1_642), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_631));
   OAI21_X1 i_0_1_1180 (.A(n_0_1_632), .B1(n_0_1_643), .B2(n_0_1_818), .ZN(
      n_0_735));
   AOI222_X1 i_0_1_1181 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[21]), .C1(n_0_1_642), .C2(A_imm_2s_complement[21]), 
      .ZN(n_0_1_632));
   OAI21_X1 i_0_1_1182 (.A(n_0_1_633), .B1(n_0_1_643), .B2(n_0_1_820), .ZN(
      n_0_736));
   AOI222_X1 i_0_1_1183 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[22]), .C1(n_0_1_642), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_633));
   OAI21_X1 i_0_1_1184 (.A(n_0_1_634), .B1(n_0_1_643), .B2(n_0_1_822), .ZN(
      n_0_737));
   AOI222_X1 i_0_1_1185 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[23]), .C1(n_0_1_642), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_634));
   OAI21_X1 i_0_1_1186 (.A(n_0_1_635), .B1(n_0_1_643), .B2(n_0_1_824), .ZN(
      n_0_738));
   AOI222_X1 i_0_1_1187 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[24]), .C1(n_0_1_642), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_635));
   OAI21_X1 i_0_1_1190 (.A(n_0_1_637), .B1(n_0_1_643), .B2(n_0_1_828), .ZN(
      n_0_740));
   AOI222_X1 i_0_1_1191 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[26]), .C1(n_0_1_642), .C2(A_imm_2s_complement[26]), 
      .ZN(n_0_1_637));
   OAI21_X1 i_0_1_1192 (.A(n_0_1_638), .B1(n_0_1_643), .B2(n_0_1_830), .ZN(
      n_0_741));
   AOI222_X1 i_0_1_1193 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[27]), .C1(n_0_1_642), .C2(A_imm_2s_complement[27]), 
      .ZN(n_0_1_638));
   OAI21_X1 i_0_1_1194 (.A(n_0_1_639), .B1(n_0_1_643), .B2(n_0_1_832), .ZN(
      n_0_742));
   AOI222_X1 i_0_1_1195 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[28]), .C1(n_0_1_642), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_639));
   OAI21_X1 i_0_1_1198 (.A(n_0_1_641), .B1(n_0_1_643), .B2(n_0_1_836), .ZN(
      n_0_744));
   AOI222_X1 i_0_1_1199 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_645), .B1(
      n_0_1_644), .B2(A_imm[30]), .C1(n_0_1_642), .C2(A_imm_2s_complement[30]), 
      .ZN(n_0_1_641));
   XNOR2_X1 i_0_1_1204 (.A(n_0_1_692), .B(n_0_1_650), .ZN(n_0_1_646));
   OAI21_X1 i_0_1_1205 (.A(n_0_1_647), .B1(n_0_1_649), .B2(n_0_1_652), .ZN(
      n_0_745));
   NAND3_X1 i_0_1_1206 (.A1(n_0_1_648), .A2(A_imm_2s_complement[31]), .A3(
      n_0_1_652), .ZN(n_0_1_647));
   NAND2_X1 i_0_1_1207 (.A1(n_0_1_693), .A2(n_0_1_650), .ZN(n_0_1_648));
   OAI21_X1 i_0_1_1208 (.A(A_imm[31]), .B1(n_0_1_693), .B2(n_0_1_650), .ZN(
      n_0_1_649));
   MUX2_X1 i_0_1_1209 (.A(n_0_180), .B(n_0_36), .S(B_in), .Z(n_0_1_650));
   INV_X1 i_0_1_1210 (.A(n_0_1_652), .ZN(n_0_1_651));
   MUX2_X1 i_0_1_1211 (.A(n_0_179), .B(n_0_37), .S(B_in), .Z(n_0_1_652));
   AND2_X1 i_0_1_1212 (.A1(n_0_1_689), .A2(n_0_155), .ZN(n_0_746));
   OAI211_X1 i_0_1_1213 (.A(n_0_1_654), .B(n_0_1_653), .C1(n_0_1_776), .C2(
      n_0_1_686), .ZN(n_0_747));
   OAI21_X1 i_0_1_1214 (.A(n_0_155), .B1(n_0_1_687), .B2(n_0_1_685), .ZN(
      n_0_1_653));
   NAND2_X1 i_0_1_1215 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_688), .ZN(
      n_0_1_654));
   OAI21_X1 i_0_1_1216 (.A(n_0_1_655), .B1(n_0_1_686), .B2(n_0_1_778), .ZN(
      n_0_748));
   AOI222_X1 i_0_1_1217 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[1]), .C1(n_0_1_685), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_655));
   OAI21_X1 i_0_1_1218 (.A(n_0_1_656), .B1(n_0_1_686), .B2(n_0_1_780), .ZN(
      n_0_749));
   AOI222_X1 i_0_1_1219 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[2]), .C1(n_0_1_685), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_656));
   OAI21_X1 i_0_1_1220 (.A(n_0_1_657), .B1(n_0_1_686), .B2(n_0_1_782), .ZN(
      n_0_750));
   AOI222_X1 i_0_1_1221 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[3]), .C1(n_0_1_685), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_657));
   OAI21_X1 i_0_1_1222 (.A(n_0_1_658), .B1(n_0_1_686), .B2(n_0_1_784), .ZN(
      n_0_751));
   AOI222_X1 i_0_1_1223 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[4]), .C1(n_0_1_685), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_658));
   OAI21_X1 i_0_1_1224 (.A(n_0_1_659), .B1(n_0_1_686), .B2(n_0_1_786), .ZN(
      n_0_752));
   AOI222_X1 i_0_1_1225 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[5]), .C1(n_0_1_685), .C2(A_imm_2s_complement[5]), 
      .ZN(n_0_1_659));
   OAI21_X1 i_0_1_1226 (.A(n_0_1_660), .B1(n_0_1_686), .B2(n_0_1_788), .ZN(
      n_0_753));
   AOI222_X1 i_0_1_1227 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[6]), .C1(n_0_1_685), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_660));
   OAI21_X1 i_0_1_1228 (.A(n_0_1_661), .B1(n_0_1_686), .B2(n_0_1_790), .ZN(
      n_0_754));
   AOI222_X1 i_0_1_1229 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[7]), .C1(n_0_1_685), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_661));
   OAI21_X1 i_0_1_1230 (.A(n_0_1_662), .B1(n_0_1_686), .B2(n_0_1_792), .ZN(
      n_0_755));
   AOI222_X1 i_0_1_1231 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[8]), .C1(n_0_1_685), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_662));
   OAI21_X1 i_0_1_1232 (.A(n_0_1_663), .B1(n_0_1_686), .B2(n_0_1_794), .ZN(
      n_0_756));
   AOI222_X1 i_0_1_1233 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[9]), .C1(n_0_1_685), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_663));
   OAI21_X1 i_0_1_1234 (.A(n_0_1_664), .B1(n_0_1_686), .B2(n_0_1_796), .ZN(
      n_0_757));
   AOI222_X1 i_0_1_1235 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[10]), .C1(n_0_1_685), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_664));
   OAI21_X1 i_0_1_1236 (.A(n_0_1_665), .B1(n_0_1_686), .B2(n_0_1_798), .ZN(
      n_0_758));
   AOI222_X1 i_0_1_1237 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[11]), .C1(n_0_1_685), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_665));
   OAI21_X1 i_0_1_1238 (.A(n_0_1_666), .B1(n_0_1_686), .B2(n_0_1_800), .ZN(
      n_0_759));
   AOI222_X1 i_0_1_1239 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[12]), .C1(n_0_1_685), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_666));
   OAI21_X1 i_0_1_1240 (.A(n_0_1_667), .B1(n_0_1_686), .B2(n_0_1_802), .ZN(
      n_0_760));
   AOI222_X1 i_0_1_1241 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[13]), .C1(n_0_1_685), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_667));
   OAI21_X1 i_0_1_1242 (.A(n_0_1_668), .B1(n_0_1_686), .B2(n_0_1_804), .ZN(
      n_0_761));
   AOI222_X1 i_0_1_1243 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[14]), .C1(n_0_1_685), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_668));
   OAI21_X1 i_0_1_1244 (.A(n_0_1_669), .B1(n_0_1_686), .B2(n_0_1_806), .ZN(
      n_0_762));
   AOI222_X1 i_0_1_1245 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[15]), .C1(n_0_1_685), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_669));
   OAI21_X1 i_0_1_1246 (.A(n_0_1_670), .B1(n_0_1_686), .B2(n_0_1_808), .ZN(
      n_0_763));
   AOI222_X1 i_0_1_1247 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[16]), .C1(n_0_1_685), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_670));
   OAI21_X1 i_0_1_1248 (.A(n_0_1_671), .B1(n_0_1_686), .B2(n_0_1_810), .ZN(
      n_0_764));
   AOI222_X1 i_0_1_1249 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[17]), .C1(n_0_1_685), .C2(A_imm_2s_complement[17]), 
      .ZN(n_0_1_671));
   OAI21_X1 i_0_1_1250 (.A(n_0_1_672), .B1(n_0_1_686), .B2(n_0_1_812), .ZN(
      n_0_765));
   AOI222_X1 i_0_1_1251 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[18]), .C1(n_0_1_685), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_672));
   OAI21_X1 i_0_1_1252 (.A(n_0_1_673), .B1(n_0_1_686), .B2(n_0_1_814), .ZN(
      n_0_766));
   AOI222_X1 i_0_1_1253 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[19]), .C1(n_0_1_685), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_673));
   OAI21_X1 i_0_1_1254 (.A(n_0_1_674), .B1(n_0_1_686), .B2(n_0_1_816), .ZN(
      n_0_767));
   AOI222_X1 i_0_1_1255 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[20]), .C1(n_0_1_685), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_674));
   OAI21_X1 i_0_1_1256 (.A(n_0_1_675), .B1(n_0_1_686), .B2(n_0_1_818), .ZN(
      n_0_768));
   AOI222_X1 i_0_1_1257 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[21]), .C1(n_0_1_685), .C2(A_imm_2s_complement[21]), 
      .ZN(n_0_1_675));
   OAI21_X1 i_0_1_1258 (.A(n_0_1_676), .B1(n_0_1_686), .B2(n_0_1_820), .ZN(
      n_0_769));
   AOI222_X1 i_0_1_1259 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[22]), .C1(n_0_1_685), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_676));
   OAI21_X1 i_0_1_1260 (.A(n_0_1_677), .B1(n_0_1_686), .B2(n_0_1_822), .ZN(
      n_0_770));
   AOI222_X1 i_0_1_1261 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[23]), .C1(n_0_1_685), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_677));
   OAI21_X1 i_0_1_1262 (.A(n_0_1_678), .B1(n_0_1_686), .B2(n_0_1_824), .ZN(
      n_0_771));
   AOI222_X1 i_0_1_1263 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[24]), .C1(n_0_1_685), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_678));
   OAI21_X1 i_0_1_1266 (.A(n_0_1_680), .B1(n_0_1_686), .B2(n_0_1_828), .ZN(
      n_0_773));
   AOI222_X1 i_0_1_1267 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[26]), .C1(n_0_1_685), .C2(A_imm_2s_complement[26]), 
      .ZN(n_0_1_680));
   OAI21_X1 i_0_1_1268 (.A(n_0_1_681), .B1(n_0_1_686), .B2(n_0_1_830), .ZN(
      n_0_774));
   AOI222_X1 i_0_1_1269 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[27]), .C1(n_0_1_685), .C2(A_imm_2s_complement[27]), 
      .ZN(n_0_1_681));
   OAI21_X1 i_0_1_1270 (.A(n_0_1_682), .B1(n_0_1_686), .B2(n_0_1_832), .ZN(
      n_0_775));
   AOI222_X1 i_0_1_1271 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[28]), .C1(n_0_1_685), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_682));
   OAI21_X1 i_0_1_1272 (.A(n_0_1_683), .B1(n_0_1_686), .B2(n_0_1_834), .ZN(
      n_0_776));
   AOI222_X1 i_0_1_1273 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[29]), .C1(n_0_1_685), .C2(A_imm_2s_complement[29]), 
      .ZN(n_0_1_683));
   OAI21_X1 i_0_1_1274 (.A(n_0_1_684), .B1(n_0_1_686), .B2(n_0_1_836), .ZN(
      n_0_777));
   AOI222_X1 i_0_1_1275 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_688), .B1(
      n_0_1_687), .B2(A_imm[30]), .C1(n_0_1_685), .C2(A_imm_2s_complement[30]), 
      .ZN(n_0_1_684));
   XNOR2_X1 i_0_1_1280 (.A(n_0_1_735), .B(n_0_1_695), .ZN(n_0_1_689));
   OAI21_X1 i_0_1_1281 (.A(n_0_1_691), .B1(n_0_1_690), .B2(n_0_1_693), .ZN(
      n_0_778));
   OAI21_X1 i_0_1_1282 (.A(A_imm[31]), .B1(n_0_1_736), .B2(n_0_1_695), .ZN(
      n_0_1_690));
   NAND3_X1 i_0_1_1283 (.A1(n_0_1_694), .A2(n_0_1_693), .A3(
      A_imm_2s_complement[31]), .ZN(n_0_1_691));
   INV_X1 i_0_1_1284 (.A(n_0_1_693), .ZN(n_0_1_692));
   MUX2_X1 i_0_1_1285 (.A(n_0_181), .B(n_0_35), .S(B_in), .Z(n_0_1_693));
   NAND2_X1 i_0_1_1286 (.A1(n_0_1_736), .A2(n_0_1_695), .ZN(n_0_1_694));
   MUX2_X1 i_0_1_1287 (.A(n_0_182), .B(n_0_34), .S(B_in), .Z(n_0_1_695));
   AND2_X1 i_0_1_1288 (.A1(n_0_1_732), .A2(n_0_155), .ZN(n_0_779));
   OAI211_X1 i_0_1_1289 (.A(n_0_1_697), .B(n_0_1_696), .C1(n_0_1_776), .C2(
      n_0_1_729), .ZN(n_0_780));
   OAI21_X1 i_0_1_1290 (.A(n_0_155), .B1(n_0_1_730), .B2(n_0_1_728), .ZN(
      n_0_1_696));
   NAND2_X1 i_0_1_1291 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_731), .ZN(
      n_0_1_697));
   OAI21_X1 i_0_1_1292 (.A(n_0_1_698), .B1(n_0_1_729), .B2(n_0_1_778), .ZN(
      n_0_781));
   AOI222_X1 i_0_1_1293 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[1]), .C1(n_0_1_728), .C2(A_imm_2s_complement[1]), 
      .ZN(n_0_1_698));
   OAI21_X1 i_0_1_1294 (.A(n_0_1_699), .B1(n_0_1_729), .B2(n_0_1_780), .ZN(
      n_0_782));
   AOI222_X1 i_0_1_1295 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[2]), .C1(n_0_1_728), .C2(A_imm_2s_complement[2]), 
      .ZN(n_0_1_699));
   OAI21_X1 i_0_1_1296 (.A(n_0_1_700), .B1(n_0_1_729), .B2(n_0_1_782), .ZN(
      n_0_783));
   AOI222_X1 i_0_1_1297 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[3]), .C1(n_0_1_728), .C2(A_imm_2s_complement[3]), 
      .ZN(n_0_1_700));
   OAI21_X1 i_0_1_1298 (.A(n_0_1_701), .B1(n_0_1_729), .B2(n_0_1_784), .ZN(
      n_0_784));
   AOI222_X1 i_0_1_1299 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[4]), .C1(n_0_1_728), .C2(A_imm_2s_complement[4]), 
      .ZN(n_0_1_701));
   OAI21_X1 i_0_1_1302 (.A(n_0_1_703), .B1(n_0_1_729), .B2(n_0_1_788), .ZN(
      n_0_786));
   AOI222_X1 i_0_1_1303 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[6]), .C1(n_0_1_728), .C2(A_imm_2s_complement[6]), 
      .ZN(n_0_1_703));
   OAI21_X1 i_0_1_1304 (.A(n_0_1_704), .B1(n_0_1_729), .B2(n_0_1_790), .ZN(
      n_0_787));
   AOI222_X1 i_0_1_1305 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[7]), .C1(n_0_1_728), .C2(A_imm_2s_complement[7]), 
      .ZN(n_0_1_704));
   OAI21_X1 i_0_1_1306 (.A(n_0_1_705), .B1(n_0_1_729), .B2(n_0_1_792), .ZN(
      n_0_788));
   AOI222_X1 i_0_1_1307 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[8]), .C1(n_0_1_728), .C2(A_imm_2s_complement[8]), 
      .ZN(n_0_1_705));
   OAI21_X1 i_0_1_1308 (.A(n_0_1_706), .B1(n_0_1_729), .B2(n_0_1_794), .ZN(
      n_0_789));
   AOI222_X1 i_0_1_1309 (.A1(A_imm_2s_complement[10]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[9]), .C1(n_0_1_728), .C2(A_imm_2s_complement[9]), 
      .ZN(n_0_1_706));
   OAI21_X1 i_0_1_1310 (.A(n_0_1_707), .B1(n_0_1_729), .B2(n_0_1_796), .ZN(
      n_0_790));
   AOI222_X1 i_0_1_1311 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[10]), .C1(n_0_1_728), .C2(A_imm_2s_complement[10]), 
      .ZN(n_0_1_707));
   OAI21_X1 i_0_1_1312 (.A(n_0_1_708), .B1(n_0_1_729), .B2(n_0_1_798), .ZN(
      n_0_791));
   AOI222_X1 i_0_1_1313 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[11]), .C1(n_0_1_728), .C2(A_imm_2s_complement[11]), 
      .ZN(n_0_1_708));
   OAI21_X1 i_0_1_1314 (.A(n_0_1_709), .B1(n_0_1_729), .B2(n_0_1_800), .ZN(
      n_0_792));
   AOI222_X1 i_0_1_1315 (.A1(A_imm_2s_complement[13]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[12]), .C1(n_0_1_728), .C2(A_imm_2s_complement[12]), 
      .ZN(n_0_1_709));
   OAI21_X1 i_0_1_1316 (.A(n_0_1_710), .B1(n_0_1_729), .B2(n_0_1_802), .ZN(
      n_0_793));
   AOI222_X1 i_0_1_1317 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[13]), .C1(n_0_1_728), .C2(A_imm_2s_complement[13]), 
      .ZN(n_0_1_710));
   OAI21_X1 i_0_1_1318 (.A(n_0_1_711), .B1(n_0_1_729), .B2(n_0_1_804), .ZN(
      n_0_794));
   AOI222_X1 i_0_1_1319 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[14]), .C1(n_0_1_728), .C2(A_imm_2s_complement[14]), 
      .ZN(n_0_1_711));
   OAI21_X1 i_0_1_1320 (.A(n_0_1_712), .B1(n_0_1_729), .B2(n_0_1_806), .ZN(
      n_0_795));
   AOI222_X1 i_0_1_1321 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[15]), .C1(n_0_1_728), .C2(A_imm_2s_complement[15]), 
      .ZN(n_0_1_712));
   OAI21_X1 i_0_1_1322 (.A(n_0_1_713), .B1(n_0_1_729), .B2(n_0_1_808), .ZN(
      n_0_796));
   AOI222_X1 i_0_1_1323 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[16]), .C1(n_0_1_728), .C2(A_imm_2s_complement[16]), 
      .ZN(n_0_1_713));
   OAI21_X1 i_0_1_1326 (.A(n_0_1_715), .B1(n_0_1_729), .B2(n_0_1_812), .ZN(
      n_0_798));
   AOI222_X1 i_0_1_1327 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[18]), .C1(n_0_1_728), .C2(A_imm_2s_complement[18]), 
      .ZN(n_0_1_715));
   OAI21_X1 i_0_1_1328 (.A(n_0_1_716), .B1(n_0_1_729), .B2(n_0_1_814), .ZN(
      n_0_799));
   AOI222_X1 i_0_1_1329 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[19]), .C1(n_0_1_728), .C2(A_imm_2s_complement[19]), 
      .ZN(n_0_1_716));
   OAI21_X1 i_0_1_1330 (.A(n_0_1_717), .B1(n_0_1_729), .B2(n_0_1_816), .ZN(
      n_0_800));
   AOI222_X1 i_0_1_1331 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[20]), .C1(n_0_1_728), .C2(A_imm_2s_complement[20]), 
      .ZN(n_0_1_717));
   OAI21_X1 i_0_1_1334 (.A(n_0_1_719), .B1(n_0_1_729), .B2(n_0_1_820), .ZN(
      n_0_802));
   AOI222_X1 i_0_1_1335 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[22]), .C1(n_0_1_728), .C2(A_imm_2s_complement[22]), 
      .ZN(n_0_1_719));
   OAI21_X1 i_0_1_1336 (.A(n_0_1_720), .B1(n_0_1_729), .B2(n_0_1_822), .ZN(
      n_0_803));
   AOI222_X1 i_0_1_1337 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[23]), .C1(n_0_1_728), .C2(A_imm_2s_complement[23]), 
      .ZN(n_0_1_720));
   OAI21_X1 i_0_1_1338 (.A(n_0_1_721), .B1(n_0_1_729), .B2(n_0_1_824), .ZN(
      n_0_804));
   AOI222_X1 i_0_1_1339 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[24]), .C1(n_0_1_728), .C2(A_imm_2s_complement[24]), 
      .ZN(n_0_1_721));
   OAI21_X1 i_0_1_1340 (.A(n_0_1_722), .B1(n_0_1_729), .B2(n_0_1_826), .ZN(
      n_0_805));
   AOI222_X1 i_0_1_1341 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[25]), .C1(n_0_1_728), .C2(A_imm_2s_complement[25]), 
      .ZN(n_0_1_722));
   OAI21_X1 i_0_1_1346 (.A(n_0_1_725), .B1(n_0_1_729), .B2(n_0_1_832), .ZN(
      n_0_808));
   AOI222_X1 i_0_1_1347 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_731), .B1(
      n_0_1_730), .B2(A_imm[28]), .C1(n_0_1_728), .C2(A_imm_2s_complement[28]), 
      .ZN(n_0_1_725));
   XNOR2_X1 i_0_1_1356 (.A(n_0_1_774), .B(n_0_1_738), .ZN(n_0_1_732));
   OAI21_X1 i_0_1_1357 (.A(n_0_1_734), .B1(n_0_1_733), .B2(n_0_1_736), .ZN(
      n_0_811));
   OAI21_X1 i_0_1_1358 (.A(A_imm[31]), .B1(n_0_1_775), .B2(n_0_1_738), .ZN(
      n_0_1_733));
   NAND3_X1 i_0_1_1359 (.A1(n_0_1_737), .A2(n_0_1_736), .A3(
      A_imm_2s_complement[31]), .ZN(n_0_1_734));
   INV_X1 i_0_1_1360 (.A(n_0_1_736), .ZN(n_0_1_735));
   MUX2_X1 i_0_1_1361 (.A(n_0_183), .B(n_0_33), .S(B_in), .Z(n_0_1_736));
   NAND2_X1 i_0_1_1362 (.A1(n_0_1_775), .A2(n_0_1_738), .ZN(n_0_1_737));
   MUX2_X1 i_0_1_1363 (.A(n_0_184), .B(n_0_32), .S(B_in), .Z(n_0_1_738));
   AND2_X1 i_0_1_1365 (.A1(n_0_186), .A2(n_0_155), .ZN(n_0_812));
   AOI22_X1 i_0_1_1367 (.A1(n_0_155), .A2(n_0_1_771), .B1(n_0_1_770), .B2(
      A_imm_2s_complement[1]), .ZN(n_0_1_739));
   OAI21_X1 i_0_1_1368 (.A(n_0_1_740), .B1(n_0_1_772), .B2(n_0_1_778), .ZN(
      n_0_814));
   AOI22_X1 i_0_1_1369 (.A1(A_imm_2s_complement[1]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[2]), .ZN(n_0_1_740));
   OAI21_X1 i_0_1_1370 (.A(n_0_1_741), .B1(n_0_1_772), .B2(n_0_1_780), .ZN(
      n_0_815));
   AOI22_X1 i_0_1_1371 (.A1(A_imm_2s_complement[2]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[3]), .ZN(n_0_1_741));
   OAI21_X1 i_0_1_1372 (.A(n_0_1_742), .B1(n_0_1_772), .B2(n_0_1_782), .ZN(
      n_0_816));
   AOI22_X1 i_0_1_1373 (.A1(A_imm_2s_complement[3]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[4]), .ZN(n_0_1_742));
   OAI21_X1 i_0_1_1374 (.A(n_0_1_743), .B1(n_0_1_772), .B2(n_0_1_784), .ZN(
      n_0_817));
   AOI22_X1 i_0_1_1375 (.A1(A_imm_2s_complement[4]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[5]), .ZN(n_0_1_743));
   OAI21_X1 i_0_1_1376 (.A(n_0_1_744), .B1(n_0_1_772), .B2(n_0_1_786), .ZN(
      n_0_818));
   AOI22_X1 i_0_1_1377 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[6]), .ZN(n_0_1_744));
   OAI21_X1 i_0_1_1378 (.A(n_0_1_745), .B1(n_0_1_772), .B2(n_0_1_788), .ZN(
      n_0_819));
   AOI22_X1 i_0_1_1379 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[7]), .ZN(n_0_1_745));
   OAI21_X1 i_0_1_1380 (.A(n_0_1_746), .B1(n_0_1_772), .B2(n_0_1_790), .ZN(
      n_0_820));
   AOI22_X1 i_0_1_1381 (.A1(A_imm_2s_complement[7]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[8]), .ZN(n_0_1_746));
   OAI21_X1 i_0_1_1382 (.A(n_0_1_747), .B1(n_0_1_772), .B2(n_0_1_792), .ZN(
      n_0_821));
   AOI22_X1 i_0_1_1383 (.A1(A_imm_2s_complement[8]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[9]), .ZN(n_0_1_747));
   OAI21_X1 i_0_1_1384 (.A(n_0_1_748), .B1(n_0_1_772), .B2(n_0_1_794), .ZN(
      n_0_822));
   AOI22_X1 i_0_1_1385 (.A1(A_imm_2s_complement[9]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[10]), .ZN(n_0_1_748));
   OAI21_X1 i_0_1_1388 (.A(n_0_1_750), .B1(n_0_1_772), .B2(n_0_1_798), .ZN(
      n_0_824));
   AOI22_X1 i_0_1_1389 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[12]), .ZN(n_0_1_750));
   OAI21_X1 i_0_1_1390 (.A(n_0_1_751), .B1(n_0_1_772), .B2(n_0_1_800), .ZN(
      n_0_825));
   AOI22_X1 i_0_1_1391 (.A1(A_imm_2s_complement[12]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[13]), .ZN(n_0_1_751));
   OAI21_X1 i_0_1_1400 (.A(n_0_1_756), .B1(n_0_1_772), .B2(n_0_1_810), .ZN(
      n_0_830));
   AOI22_X1 i_0_1_1401 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[18]), .ZN(n_0_1_756));
   OAI21_X1 i_0_1_1402 (.A(n_0_1_757), .B1(n_0_1_772), .B2(n_0_1_812), .ZN(
      n_0_831));
   AOI22_X1 i_0_1_1403 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[19]), .ZN(n_0_1_757));
   OAI21_X1 i_0_1_1404 (.A(n_0_1_758), .B1(n_0_1_772), .B2(n_0_1_814), .ZN(
      n_0_832));
   AOI22_X1 i_0_1_1405 (.A1(A_imm_2s_complement[19]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[20]), .ZN(n_0_1_758));
   OAI21_X1 i_0_1_1406 (.A(n_0_1_759), .B1(n_0_1_772), .B2(n_0_1_816), .ZN(
      n_0_833));
   AOI22_X1 i_0_1_1407 (.A1(A_imm_2s_complement[20]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[21]), .ZN(n_0_1_759));
   OAI21_X1 i_0_1_1408 (.A(n_0_1_760), .B1(n_0_1_772), .B2(n_0_1_818), .ZN(
      n_0_834));
   AOI22_X1 i_0_1_1409 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[22]), .ZN(n_0_1_760));
   OAI21_X1 i_0_1_1410 (.A(n_0_1_761), .B1(n_0_1_772), .B2(n_0_1_820), .ZN(
      n_0_835));
   AOI22_X1 i_0_1_1411 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[23]), .ZN(n_0_1_761));
   OAI21_X1 i_0_1_1412 (.A(n_0_1_762), .B1(n_0_1_772), .B2(n_0_1_822), .ZN(
      n_0_836));
   AOI22_X1 i_0_1_1413 (.A1(A_imm_2s_complement[23]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[24]), .ZN(n_0_1_762));
   OAI21_X1 i_0_1_1414 (.A(n_0_1_763), .B1(n_0_1_772), .B2(n_0_1_824), .ZN(
      n_0_837));
   AOI22_X1 i_0_1_1415 (.A1(A_imm_2s_complement[24]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[25]), .ZN(n_0_1_763));
   OAI21_X1 i_0_1_1416 (.A(n_0_1_764), .B1(n_0_1_772), .B2(n_0_1_826), .ZN(
      n_0_838));
   AOI22_X1 i_0_1_1417 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[26]), .ZN(n_0_1_764));
   OAI21_X1 i_0_1_1418 (.A(n_0_1_765), .B1(n_0_1_772), .B2(n_0_1_828), .ZN(
      n_0_839));
   AOI22_X1 i_0_1_1419 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[27]), .ZN(n_0_1_765));
   OAI21_X1 i_0_1_1420 (.A(n_0_1_766), .B1(n_0_1_772), .B2(n_0_1_830), .ZN(
      n_0_840));
   AOI22_X1 i_0_1_1421 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[28]), .ZN(n_0_1_766));
   OAI21_X1 i_0_1_1424 (.A(n_0_1_768), .B1(n_0_1_772), .B2(n_0_1_834), .ZN(
      n_0_842));
   AOI22_X1 i_0_1_1425 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_771), .B1(
      n_0_1_770), .B2(A_imm_2s_complement[30]), .ZN(n_0_1_768));
   INV_X1 i_0_1_1433 (.A(n_0_1_775), .ZN(n_0_1_774));
   INV_X1 i_0_1_1441 (.A(n_0_1_780), .ZN(A_imm[3]));
   AOI21_X1 i_0_1_1442 (.A(n_0_1_781), .B1(n_0_2), .B2(A_in), .ZN(n_0_1_780));
   NOR2_X1 i_0_1_1443 (.A1(n_0_1_840), .A2(A_in), .ZN(n_0_1_781));
   INV_X1 i_0_1_1444 (.A(n_0_1_782), .ZN(A_imm[4]));
   AOI21_X1 i_0_1_1445 (.A(n_0_1_783), .B1(n_0_3), .B2(A_in), .ZN(n_0_1_782));
   NOR2_X1 i_0_1_1446 (.A1(n_0_1_841), .A2(A_in), .ZN(n_0_1_783));
   INV_X1 i_0_1_1450 (.A(n_0_1_786), .ZN(A_imm[6]));
   NOR2_X1 i_0_1_1452 (.A1(n_0_1_843), .A2(A_in), .ZN(n_0_1_787));
   INV_X1 i_0_1_1453 (.A(n_0_1_788), .ZN(A_imm[7]));
   AOI21_X1 i_0_1_1454 (.A(n_0_1_789), .B1(n_0_6), .B2(A_in), .ZN(n_0_1_788));
   NOR2_X1 i_0_1_1455 (.A1(n_0_1_844), .A2(A_in), .ZN(n_0_1_789));
   INV_X1 i_0_1_1456 (.A(n_0_1_790), .ZN(A_imm[8]));
   AOI21_X1 i_0_1_1457 (.A(n_0_1_791), .B1(n_0_7), .B2(A_in), .ZN(n_0_1_790));
   NOR2_X1 i_0_1_1458 (.A1(n_0_1_845), .A2(A_in), .ZN(n_0_1_791));
   INV_X1 i_0_1_1459 (.A(n_0_1_792), .ZN(A_imm[9]));
   AOI21_X1 i_0_1_1460 (.A(n_0_1_793), .B1(n_0_8), .B2(A_in), .ZN(n_0_1_792));
   NOR2_X1 i_0_1_1461 (.A1(n_0_1_846), .A2(A_in), .ZN(n_0_1_793));
   INV_X1 i_0_1_1462 (.A(n_0_1_794), .ZN(A_imm[10]));
   AOI21_X1 i_0_1_1463 (.A(n_0_1_795), .B1(n_0_9), .B2(A_in), .ZN(n_0_1_794));
   NOR2_X1 i_0_1_1464 (.A1(n_0_1_847), .A2(A_in), .ZN(n_0_1_795));
   INV_X1 i_0_1_1465 (.A(n_0_1_796), .ZN(A_imm[11]));
   NOR2_X1 i_0_1_1467 (.A1(n_0_1_848), .A2(A_in), .ZN(n_0_1_797));
   INV_X1 i_0_1_1468 (.A(n_0_1_798), .ZN(A_imm[12]));
   AOI21_X1 i_0_1_1469 (.A(n_0_1_799), .B1(n_0_11), .B2(A_in), .ZN(n_0_1_798));
   NOR2_X1 i_0_1_1470 (.A1(n_0_1_849), .A2(A_in), .ZN(n_0_1_799));
   INV_X1 i_0_1_1471 (.A(n_0_1_800), .ZN(A_imm[13]));
   AOI21_X1 i_0_1_1472 (.A(n_0_1_801), .B1(n_0_12), .B2(A_in), .ZN(n_0_1_800));
   NOR2_X1 i_0_1_1473 (.A1(n_0_1_850), .A2(A_in), .ZN(n_0_1_801));
   INV_X1 i_0_1_1474 (.A(n_0_1_802), .ZN(A_imm[14]));
   NOR2_X1 i_0_1_1476 (.A1(n_0_1_851), .A2(A_in), .ZN(n_0_1_803));
   INV_X1 i_0_1_1477 (.A(n_0_1_804), .ZN(A_imm[15]));
   NOR2_X1 i_0_1_1479 (.A1(n_0_1_852), .A2(A_in), .ZN(n_0_1_805));
   INV_X1 i_0_1_1480 (.A(n_0_1_806), .ZN(A_imm[16]));
   NOR2_X1 i_0_1_1482 (.A1(n_0_1_853), .A2(A_in), .ZN(n_0_1_807));
   NOR2_X1 i_0_1_1485 (.A1(n_0_1_854), .A2(A_in), .ZN(n_0_1_809));
   INV_X1 i_0_1_1486 (.A(n_0_1_810), .ZN(A_imm[18]));
   NOR2_X1 i_0_1_1488 (.A1(n_0_1_855), .A2(A_in), .ZN(n_0_1_811));
   INV_X1 i_0_1_1489 (.A(n_0_1_812), .ZN(A_imm[19]));
   AOI21_X1 i_0_1_1490 (.A(n_0_1_813), .B1(n_0_18), .B2(A_in), .ZN(n_0_1_812));
   NOR2_X1 i_0_1_1491 (.A1(n_0_1_856), .A2(A_in), .ZN(n_0_1_813));
   INV_X1 i_0_1_1492 (.A(n_0_1_814), .ZN(A_imm[20]));
   AOI21_X1 i_0_1_1493 (.A(n_0_1_815), .B1(n_0_19), .B2(A_in), .ZN(n_0_1_814));
   NOR2_X1 i_0_1_1494 (.A1(n_0_1_857), .A2(A_in), .ZN(n_0_1_815));
   AOI21_X1 i_0_1_1496 (.A(n_0_1_817), .B1(n_0_20), .B2(A_in), .ZN(n_0_1_816));
   NOR2_X1 i_0_1_1497 (.A1(n_0_1_858), .A2(A_in), .ZN(n_0_1_817));
   INV_X1 i_0_1_1498 (.A(n_0_1_818), .ZN(A_imm[22]));
   NOR2_X1 i_0_1_1500 (.A1(n_0_1_859), .A2(A_in), .ZN(n_0_1_819));
   INV_X1 i_0_1_1501 (.A(n_0_1_820), .ZN(A_imm[23]));
   AOI21_X1 i_0_1_1502 (.A(n_0_1_821), .B1(n_0_22), .B2(A_in), .ZN(n_0_1_820));
   NOR2_X1 i_0_1_1503 (.A1(n_0_1_860), .A2(A_in), .ZN(n_0_1_821));
   INV_X1 i_0_1_1504 (.A(n_0_1_822), .ZN(A_imm[24]));
   AOI21_X1 i_0_1_1505 (.A(n_0_1_823), .B1(n_0_23), .B2(A_in), .ZN(n_0_1_822));
   NOR2_X1 i_0_1_1506 (.A1(n_0_1_861), .A2(A_in), .ZN(n_0_1_823));
   AOI21_X1 i_0_1_1508 (.A(n_0_1_825), .B1(n_0_24), .B2(A_in), .ZN(n_0_1_824));
   NOR2_X1 i_0_1_1509 (.A1(n_0_1_862), .A2(A_in), .ZN(n_0_1_825));
   NOR2_X1 i_0_1_1512 (.A1(n_0_1_863), .A2(A_in), .ZN(n_0_1_827));
   NOR2_X1 i_0_1_1515 (.A1(n_0_1_864), .A2(A_in), .ZN(n_0_1_829));
   INV_X1 i_0_1_1516 (.A(n_0_1_830), .ZN(A_imm[28]));
   NOR2_X1 i_0_1_1518 (.A1(n_0_1_865), .A2(A_in), .ZN(n_0_1_831));
   NOR2_X1 i_0_1_1521 (.A1(n_0_1_866), .A2(A_in), .ZN(n_0_1_833));
   NOR2_X1 i_0_1_1524 (.A1(n_0_1_867), .A2(A_in), .ZN(n_0_1_835));
   INV_X1 i_0_1_1525 (.A(n_0_1_836), .ZN(A_imm[31]));
   INV_X1 i_0_1_1529 (.A(n_0_153), .ZN(n_0_1_839));
   INV_X1 i_0_1_1530 (.A(n_0_152), .ZN(n_0_1_840));
   INV_X1 i_0_1_1531 (.A(n_0_151), .ZN(n_0_1_841));
   INV_X1 i_0_1_1532 (.A(n_0_150), .ZN(n_0_1_842));
   INV_X1 i_0_1_1533 (.A(n_0_149), .ZN(n_0_1_843));
   INV_X1 i_0_1_1534 (.A(n_0_148), .ZN(n_0_1_844));
   INV_X1 i_0_1_1535 (.A(n_0_147), .ZN(n_0_1_845));
   INV_X1 i_0_1_1536 (.A(n_0_146), .ZN(n_0_1_846));
   INV_X1 i_0_1_1537 (.A(n_0_145), .ZN(n_0_1_847));
   INV_X1 i_0_1_1538 (.A(n_0_144), .ZN(n_0_1_848));
   INV_X1 i_0_1_1539 (.A(n_0_143), .ZN(n_0_1_849));
   INV_X1 i_0_1_1540 (.A(n_0_142), .ZN(n_0_1_850));
   INV_X1 i_0_1_1541 (.A(n_0_141), .ZN(n_0_1_851));
   INV_X1 i_0_1_1542 (.A(n_0_140), .ZN(n_0_1_852));
   INV_X1 i_0_1_1543 (.A(n_0_139), .ZN(n_0_1_853));
   INV_X1 i_0_1_1544 (.A(n_0_138), .ZN(n_0_1_854));
   INV_X1 i_0_1_1545 (.A(n_0_137), .ZN(n_0_1_855));
   INV_X1 i_0_1_1546 (.A(n_0_136), .ZN(n_0_1_856));
   INV_X1 i_0_1_1547 (.A(n_0_135), .ZN(n_0_1_857));
   INV_X1 i_0_1_1548 (.A(n_0_134), .ZN(n_0_1_858));
   INV_X1 i_0_1_1549 (.A(n_0_133), .ZN(n_0_1_859));
   INV_X1 i_0_1_1550 (.A(n_0_132), .ZN(n_0_1_860));
   INV_X1 i_0_1_1551 (.A(n_0_131), .ZN(n_0_1_861));
   INV_X1 i_0_1_1552 (.A(n_0_130), .ZN(n_0_1_862));
   INV_X1 i_0_1_1553 (.A(n_0_129), .ZN(n_0_1_863));
   INV_X1 i_0_1_1554 (.A(n_0_128), .ZN(n_0_1_864));
   INV_X1 i_0_1_1555 (.A(n_0_127), .ZN(n_0_1_865));
   INV_X1 i_0_1_1556 (.A(n_0_126), .ZN(n_0_1_866));
   INV_X1 i_0_1_1557 (.A(n_0_125), .ZN(n_0_1_867));
   INV_X1 i_0_1_1558 (.A(n_0_157), .ZN(n_0_1_868));
   INV_X1 i_0_1_1 (.A(A_imm[5]), .ZN(n_0_1_784));
   INV_X1 i_0_1_2 (.A(A_imm[1]), .ZN(n_0_1_776));
   OAI22_X1 i_0_1_3 (.A1(n_0_1_767), .A2(n_0_1_0), .B1(n_0_1_907), .B2(n_0_1_1), 
      .ZN(n_0_188));
   INV_X1 i_0_1_4 (.A(n_0_62), .ZN(n_0_1_0));
   OAI22_X1 i_0_1_5 (.A1(n_0_1_767), .A2(n_0_1_2), .B1(n_0_1_903), .B2(n_0_1_1), 
      .ZN(n_0_189));
   NAND2_X1 i_0_1_6 (.A1(n_0_1_908), .A2(n_0_1_837), .ZN(n_0_1_1));
   INV_X1 i_0_1_7 (.A(n_0_63), .ZN(n_0_1_2));
   OAI21_X1 i_0_1_8 (.A(n_0_1_3), .B1(n_0_1_752), .B2(n_0_1_904), .ZN(n_0_190));
   NAND2_X1 i_0_1_9 (.A1(n_0_1_702), .A2(n_0_64), .ZN(n_0_1_3));
   OAI21_X1 i_0_1_10 (.A(n_0_1_4), .B1(n_0_1_752), .B2(n_0_1_905), .ZN(n_0_191));
   NAND2_X1 i_0_1_11 (.A1(n_0_1_702), .A2(n_0_65), .ZN(n_0_1_4));
   OAI21_X1 i_0_1_12 (.A(n_0_1_5), .B1(n_0_1_752), .B2(n_0_1_906), .ZN(n_0_192));
   NAND2_X1 i_0_1_13 (.A1(n_0_1_702), .A2(n_0_66), .ZN(n_0_1_5));
   OAI21_X1 i_0_1_14 (.A(n_0_1_6), .B1(n_0_1_752), .B2(n_0_1_898), .ZN(n_0_193));
   NAND2_X1 i_0_1_15 (.A1(n_0_1_702), .A2(n_0_67), .ZN(n_0_1_6));
   OAI21_X1 i_0_1_16 (.A(n_0_1_7), .B1(n_0_1_752), .B2(n_0_1_899), .ZN(n_0_194));
   NAND2_X1 i_0_1_17 (.A1(n_0_1_702), .A2(n_0_68), .ZN(n_0_1_7));
   OAI21_X1 i_0_1_18 (.A(n_0_1_8), .B1(n_0_1_752), .B2(n_0_1_900), .ZN(n_0_195));
   NAND2_X1 i_0_1_19 (.A1(n_0_1_702), .A2(n_0_69), .ZN(n_0_1_8));
   OAI21_X1 i_0_1_20 (.A(n_0_1_9), .B1(n_0_1_752), .B2(n_0_1_901), .ZN(n_0_196));
   NAND2_X1 i_0_1_21 (.A1(n_0_1_702), .A2(n_0_70), .ZN(n_0_1_9));
   OAI21_X1 i_0_1_22 (.A(n_0_1_10), .B1(n_0_1_752), .B2(n_0_1_872), .ZN(n_0_197));
   NAND2_X1 i_0_1_23 (.A1(n_0_1_702), .A2(n_0_71), .ZN(n_0_1_10));
   OAI21_X1 i_0_1_24 (.A(n_0_1_11), .B1(n_0_1_752), .B2(n_0_1_873), .ZN(n_0_198));
   NAND2_X1 i_0_1_25 (.A1(n_0_1_702), .A2(n_0_72), .ZN(n_0_1_11));
   OAI21_X1 i_0_1_26 (.A(n_0_1_12), .B1(n_0_1_752), .B2(n_0_1_874), .ZN(n_0_199));
   NAND2_X1 i_0_1_27 (.A1(n_0_1_702), .A2(n_0_73), .ZN(n_0_1_12));
   OAI21_X1 i_0_1_28 (.A(n_0_1_13), .B1(n_0_1_752), .B2(n_0_1_875), .ZN(n_0_200));
   NAND2_X1 i_0_1_29 (.A1(n_0_1_702), .A2(n_0_74), .ZN(n_0_1_13));
   OAI21_X1 i_0_1_30 (.A(n_0_1_14), .B1(n_0_1_752), .B2(n_0_1_884), .ZN(n_0_201));
   NAND2_X1 i_0_1_31 (.A1(n_0_1_702), .A2(n_0_75), .ZN(n_0_1_14));
   OAI21_X1 i_0_1_32 (.A(n_0_1_15), .B1(n_0_1_752), .B2(n_0_1_885), .ZN(n_0_202));
   NAND2_X1 i_0_1_33 (.A1(n_0_1_702), .A2(n_0_76), .ZN(n_0_1_15));
   OAI21_X1 i_0_1_34 (.A(n_0_1_16), .B1(n_0_1_752), .B2(n_0_1_17), .ZN(n_0_203));
   NAND2_X1 i_0_1_35 (.A1(n_0_1_702), .A2(n_0_77), .ZN(n_0_1_16));
   INV_X1 i_0_1_36 (.A(\aggregated_res[14] [16]), .ZN(n_0_1_17));
   OAI21_X1 i_0_1_37 (.A(n_0_1_18), .B1(n_0_1_752), .B2(n_0_1_19), .ZN(n_0_204));
   NAND2_X1 i_0_1_38 (.A1(n_0_1_702), .A2(n_0_78), .ZN(n_0_1_18));
   INV_X1 i_0_1_39 (.A(\aggregated_res[14] [17]), .ZN(n_0_1_19));
   OAI21_X1 i_0_1_40 (.A(n_0_1_20), .B1(n_0_1_752), .B2(n_0_1_21), .ZN(n_0_205));
   NAND2_X1 i_0_1_41 (.A1(n_0_1_702), .A2(n_0_79), .ZN(n_0_1_20));
   INV_X1 i_0_1_42 (.A(\aggregated_res[14] [18]), .ZN(n_0_1_21));
   OAI21_X1 i_0_1_43 (.A(n_0_1_22), .B1(n_0_1_752), .B2(n_0_1_23), .ZN(n_0_206));
   NAND2_X1 i_0_1_44 (.A1(n_0_1_702), .A2(n_0_80), .ZN(n_0_1_22));
   INV_X1 i_0_1_45 (.A(\aggregated_res[14] [19]), .ZN(n_0_1_23));
   OAI21_X1 i_0_1_46 (.A(n_0_1_24), .B1(n_0_1_752), .B2(n_0_1_25), .ZN(n_0_207));
   NAND2_X1 i_0_1_47 (.A1(n_0_1_702), .A2(n_0_81), .ZN(n_0_1_24));
   INV_X1 i_0_1_48 (.A(\aggregated_res[14] [20]), .ZN(n_0_1_25));
   OAI21_X1 i_0_1_49 (.A(n_0_1_26), .B1(n_0_1_752), .B2(n_0_1_27), .ZN(n_0_208));
   NAND2_X1 i_0_1_50 (.A1(n_0_1_702), .A2(n_0_82), .ZN(n_0_1_26));
   INV_X1 i_0_1_51 (.A(\aggregated_res[14] [21]), .ZN(n_0_1_27));
   OAI21_X1 i_0_1_52 (.A(n_0_1_28), .B1(n_0_1_752), .B2(n_0_1_29), .ZN(n_0_209));
   NAND2_X1 i_0_1_53 (.A1(n_0_1_702), .A2(n_0_83), .ZN(n_0_1_28));
   INV_X1 i_0_1_54 (.A(\aggregated_res[14] [22]), .ZN(n_0_1_29));
   OAI21_X1 i_0_1_55 (.A(n_0_1_30), .B1(n_0_1_752), .B2(n_0_1_31), .ZN(n_0_210));
   NAND2_X1 i_0_1_56 (.A1(n_0_1_702), .A2(n_0_84), .ZN(n_0_1_30));
   INV_X1 i_0_1_57 (.A(\aggregated_res[14] [23]), .ZN(n_0_1_31));
   OAI21_X1 i_0_1_58 (.A(n_0_1_32), .B1(n_0_1_752), .B2(n_0_1_33), .ZN(n_0_211));
   NAND2_X1 i_0_1_59 (.A1(n_0_1_702), .A2(n_0_85), .ZN(n_0_1_32));
   INV_X1 i_0_1_60 (.A(\aggregated_res[14] [24]), .ZN(n_0_1_33));
   OAI21_X1 i_0_1_61 (.A(n_0_1_34), .B1(n_0_1_752), .B2(n_0_1_35), .ZN(n_0_212));
   NAND2_X1 i_0_1_62 (.A1(n_0_1_702), .A2(n_0_86), .ZN(n_0_1_34));
   INV_X1 i_0_1_63 (.A(\aggregated_res[14] [25]), .ZN(n_0_1_35));
   OAI21_X1 i_0_1_64 (.A(n_0_1_36), .B1(n_0_1_752), .B2(n_0_1_37), .ZN(n_0_213));
   NAND2_X1 i_0_1_65 (.A1(n_0_1_702), .A2(n_0_87), .ZN(n_0_1_36));
   INV_X1 i_0_1_66 (.A(\aggregated_res[14] [26]), .ZN(n_0_1_37));
   OAI21_X1 i_0_1_67 (.A(n_0_1_38), .B1(n_0_1_752), .B2(n_0_1_39), .ZN(n_0_214));
   NAND2_X1 i_0_1_68 (.A1(n_0_1_702), .A2(n_0_88), .ZN(n_0_1_38));
   INV_X1 i_0_1_69 (.A(\aggregated_res[14] [27]), .ZN(n_0_1_39));
   OAI21_X1 i_0_1_70 (.A(n_0_1_40), .B1(n_0_1_752), .B2(n_0_1_41), .ZN(n_0_215));
   NAND2_X1 i_0_1_71 (.A1(n_0_1_702), .A2(n_0_89), .ZN(n_0_1_40));
   INV_X1 i_0_1_72 (.A(\aggregated_res[14] [28]), .ZN(n_0_1_41));
   OAI21_X1 i_0_1_73 (.A(n_0_1_42), .B1(n_0_1_752), .B2(n_0_1_43), .ZN(n_0_216));
   NAND2_X1 i_0_1_74 (.A1(n_0_1_702), .A2(n_0_90), .ZN(n_0_1_42));
   INV_X1 i_0_1_75 (.A(\aggregated_res[14] [29]), .ZN(n_0_1_43));
   OAI21_X1 i_0_1_76 (.A(n_0_1_44), .B1(n_0_1_752), .B2(n_0_1_45), .ZN(n_0_217));
   NAND2_X1 i_0_1_77 (.A1(n_0_1_702), .A2(n_0_91), .ZN(n_0_1_44));
   INV_X1 i_0_1_78 (.A(\aggregated_res[14] [30]), .ZN(n_0_1_45));
   OAI21_X1 i_0_1_79 (.A(n_0_1_46), .B1(n_0_1_752), .B2(n_0_1_886), .ZN(n_0_218));
   NAND2_X1 i_0_1_80 (.A1(n_0_1_702), .A2(n_0_92), .ZN(n_0_1_46));
   OAI21_X1 i_0_1_81 (.A(n_0_1_47), .B1(n_0_1_752), .B2(n_0_1_887), .ZN(n_0_219));
   NAND2_X1 i_0_1_82 (.A1(n_0_1_702), .A2(n_0_93), .ZN(n_0_1_47));
   OAI21_X1 i_0_1_83 (.A(n_0_1_48), .B1(n_0_1_752), .B2(n_0_1_49), .ZN(n_0_220));
   NAND2_X1 i_0_1_84 (.A1(n_0_1_702), .A2(n_0_94), .ZN(n_0_1_48));
   INV_X1 i_0_1_85 (.A(\aggregated_res[14] [33]), .ZN(n_0_1_49));
   OAI21_X1 i_0_1_86 (.A(n_0_1_50), .B1(n_0_1_752), .B2(n_0_1_51), .ZN(n_0_221));
   NAND2_X1 i_0_1_87 (.A1(n_0_1_702), .A2(n_0_95), .ZN(n_0_1_50));
   INV_X1 i_0_1_88 (.A(\aggregated_res[14] [34]), .ZN(n_0_1_51));
   OAI21_X1 i_0_1_89 (.A(n_0_1_52), .B1(n_0_1_752), .B2(n_0_1_53), .ZN(n_0_222));
   NAND2_X1 i_0_1_90 (.A1(n_0_1_702), .A2(n_0_96), .ZN(n_0_1_52));
   INV_X1 i_0_1_91 (.A(\aggregated_res[14] [35]), .ZN(n_0_1_53));
   OAI21_X1 i_0_1_92 (.A(n_0_1_54), .B1(n_0_1_752), .B2(n_0_1_55), .ZN(n_0_223));
   NAND2_X1 i_0_1_93 (.A1(n_0_1_702), .A2(n_0_97), .ZN(n_0_1_54));
   INV_X1 i_0_1_94 (.A(\aggregated_res[14] [36]), .ZN(n_0_1_55));
   OAI21_X1 i_0_1_95 (.A(n_0_1_56), .B1(n_0_1_752), .B2(n_0_1_57), .ZN(n_0_224));
   NAND2_X1 i_0_1_96 (.A1(n_0_1_702), .A2(n_0_98), .ZN(n_0_1_56));
   INV_X1 i_0_1_97 (.A(\aggregated_res[14] [37]), .ZN(n_0_1_57));
   OAI21_X1 i_0_1_98 (.A(n_0_1_58), .B1(n_0_1_752), .B2(n_0_1_59), .ZN(n_0_225));
   NAND2_X1 i_0_1_99 (.A1(n_0_1_702), .A2(n_0_99), .ZN(n_0_1_58));
   INV_X1 i_0_1_100 (.A(\aggregated_res[14] [38]), .ZN(n_0_1_59));
   OAI21_X1 i_0_1_101 (.A(n_0_1_60), .B1(n_0_1_752), .B2(n_0_1_61), .ZN(n_0_226));
   NAND2_X1 i_0_1_102 (.A1(n_0_1_702), .A2(n_0_100), .ZN(n_0_1_60));
   INV_X1 i_0_1_103 (.A(\aggregated_res[14] [39]), .ZN(n_0_1_61));
   OAI21_X1 i_0_1_104 (.A(n_0_1_62), .B1(n_0_1_752), .B2(n_0_1_63), .ZN(n_0_227));
   NAND2_X1 i_0_1_105 (.A1(n_0_1_702), .A2(n_0_101), .ZN(n_0_1_62));
   INV_X1 i_0_1_106 (.A(\aggregated_res[14] [40]), .ZN(n_0_1_63));
   OAI21_X1 i_0_1_107 (.A(n_0_1_64), .B1(n_0_1_752), .B2(n_0_1_65), .ZN(n_0_228));
   NAND2_X1 i_0_1_108 (.A1(n_0_1_702), .A2(n_0_102), .ZN(n_0_1_64));
   INV_X1 i_0_1_109 (.A(\aggregated_res[14] [41]), .ZN(n_0_1_65));
   OAI21_X1 i_0_1_110 (.A(n_0_1_66), .B1(n_0_1_752), .B2(n_0_1_67), .ZN(n_0_229));
   NAND2_X1 i_0_1_111 (.A1(n_0_1_702), .A2(n_0_103), .ZN(n_0_1_66));
   INV_X1 i_0_1_112 (.A(\aggregated_res[14] [42]), .ZN(n_0_1_67));
   OAI21_X1 i_0_1_113 (.A(n_0_1_68), .B1(n_0_1_752), .B2(n_0_1_69), .ZN(n_0_230));
   NAND2_X1 i_0_1_114 (.A1(n_0_1_702), .A2(n_0_104), .ZN(n_0_1_68));
   INV_X1 i_0_1_115 (.A(\aggregated_res[14] [43]), .ZN(n_0_1_69));
   OAI21_X1 i_0_1_116 (.A(n_0_1_70), .B1(n_0_1_752), .B2(n_0_1_71), .ZN(n_0_231));
   NAND2_X1 i_0_1_117 (.A1(n_0_1_702), .A2(n_0_105), .ZN(n_0_1_70));
   INV_X1 i_0_1_118 (.A(\aggregated_res[14] [44]), .ZN(n_0_1_71));
   OAI21_X1 i_0_1_119 (.A(n_0_1_72), .B1(n_0_1_752), .B2(n_0_1_73), .ZN(n_0_232));
   NAND2_X1 i_0_1_120 (.A1(n_0_1_702), .A2(n_0_106), .ZN(n_0_1_72));
   INV_X1 i_0_1_121 (.A(\aggregated_res[14] [45]), .ZN(n_0_1_73));
   OAI21_X1 i_0_1_122 (.A(n_0_1_78), .B1(n_0_1_752), .B2(n_0_1_83), .ZN(n_0_233));
   NAND2_X1 i_0_1_123 (.A1(n_0_1_702), .A2(n_0_107), .ZN(n_0_1_78));
   INV_X1 i_0_1_124 (.A(\aggregated_res[14] [46]), .ZN(n_0_1_83));
   OAI21_X1 i_0_1_125 (.A(n_0_1_84), .B1(n_0_1_752), .B2(n_0_1_889), .ZN(n_0_234));
   NAND2_X1 i_0_1_126 (.A1(n_0_1_702), .A2(n_0_108), .ZN(n_0_1_84));
   OAI21_X1 i_0_1_127 (.A(n_0_1_85), .B1(n_0_1_752), .B2(n_0_1_890), .ZN(n_0_235));
   NAND2_X1 i_0_1_128 (.A1(n_0_1_702), .A2(n_0_109), .ZN(n_0_1_85));
   OAI22_X1 i_0_1_129 (.A1(n_0_1_86), .A2(n_0_1_767), .B1(n_0_1_891), .B2(
      n_0_1_752), .ZN(n_0_236));
   INV_X1 i_0_1_130 (.A(n_0_110), .ZN(n_0_1_86));
   OAI22_X1 i_0_1_131 (.A1(n_0_1_87), .A2(n_0_1_767), .B1(n_0_1_892), .B2(
      n_0_1_752), .ZN(n_0_237));
   INV_X1 i_0_1_132 (.A(n_0_111), .ZN(n_0_1_87));
   NAND2_X1 i_0_1_133 (.A1(n_0_1_89), .A2(n_0_1_88), .ZN(n_0_238));
   NAND2_X1 i_0_1_134 (.A1(n_0_1_755), .A2(\aggregated_res[14] [51]), .ZN(
      n_0_1_88));
   NAND2_X1 i_0_1_135 (.A1(n_0_112), .A2(n_0_1_702), .ZN(n_0_1_89));
   OAI21_X1 i_0_1_136 (.A(n_0_1_554), .B1(n_0_1_555), .B2(n_0_1_767), .ZN(
      n_0_239));
   NAND2_X1 i_0_1_137 (.A1(n_0_1_755), .A2(\aggregated_res[14] [52]), .ZN(
      n_0_1_554));
   INV_X1 i_0_1_142 (.A(n_0_113), .ZN(n_0_1_555));
   OAI21_X1 i_0_1_147 (.A(n_0_1_589), .B1(n_0_1_597), .B2(n_0_1_767), .ZN(
      n_0_240));
   NAND2_X1 i_0_1_148 (.A1(n_0_1_755), .A2(\aggregated_res[14] [53]), .ZN(
      n_0_1_589));
   INV_X1 i_0_1_149 (.A(n_0_114), .ZN(n_0_1_597));
   OAI21_X1 i_0_1_150 (.A(n_0_1_636), .B1(n_0_1_640), .B2(n_0_1_767), .ZN(
      n_0_241));
   NAND2_X1 i_0_1_151 (.A1(n_0_1_755), .A2(\aggregated_res[14] [54]), .ZN(
      n_0_1_636));
   INV_X1 i_0_1_152 (.A(n_0_115), .ZN(n_0_1_640));
   OAI21_X1 i_0_1_153 (.A(n_0_1_679), .B1(n_0_1_752), .B2(n_0_1_878), .ZN(
      n_0_242));
   NAND2_X1 i_0_1_154 (.A1(n_0_116), .A2(n_0_1_702), .ZN(n_0_1_679));
   INV_X1 i_0_1_155 (.A(n_0_1_767), .ZN(n_0_1_702));
   OAI22_X1 i_0_1_156 (.A1(n_0_1_714), .A2(n_0_1_767), .B1(n_0_1_879), .B2(
      n_0_1_752), .ZN(n_0_243));
   INV_X1 i_0_1_157 (.A(n_0_117), .ZN(n_0_1_714));
   OAI22_X1 i_0_1_158 (.A1(n_0_1_718), .A2(n_0_1_767), .B1(n_0_1_880), .B2(
      n_0_1_752), .ZN(n_0_244));
   INV_X1 i_0_1_159 (.A(n_0_118), .ZN(n_0_1_718));
   OAI22_X1 i_0_1_160 (.A1(n_0_1_723), .A2(n_0_1_767), .B1(n_0_1_881), .B2(
      n_0_1_752), .ZN(n_0_245));
   INV_X1 i_0_1_161 (.A(n_0_119), .ZN(n_0_1_723));
   OAI21_X1 i_0_1_162 (.A(n_0_1_724), .B1(n_0_1_726), .B2(n_0_1_767), .ZN(
      n_0_246));
   NAND2_X1 i_0_1_163 (.A1(n_0_1_755), .A2(\aggregated_res[14] [59]), .ZN(
      n_0_1_724));
   INV_X1 i_0_1_164 (.A(n_0_120), .ZN(n_0_1_726));
   OAI22_X1 i_0_1_165 (.A1(n_0_1_727), .A2(n_0_1_767), .B1(n_0_1_838), .B2(
      n_0_1_752), .ZN(n_0_247));
   INV_X1 i_0_1_166 (.A(n_0_121), .ZN(n_0_1_727));
   OAI22_X1 i_0_1_167 (.A1(n_0_1_749), .A2(n_0_1_767), .B1(n_0_1_869), .B2(
      n_0_1_752), .ZN(n_0_248));
   INV_X1 i_0_1_168 (.A(n_0_122), .ZN(n_0_1_749));
   OAI22_X1 i_0_1_169 (.A1(n_0_1_753), .A2(n_0_1_767), .B1(n_0_1_870), .B2(
      n_0_1_752), .ZN(n_0_249));
   INV_X1 i_0_1_170 (.A(n_0_1_755), .ZN(n_0_1_752));
   INV_X1 i_0_1_171 (.A(n_0_123), .ZN(n_0_1_753));
   OAI21_X1 i_0_1_172 (.A(n_0_1_754), .B1(n_0_1_909), .B2(n_0_1_767), .ZN(
      n_0_250));
   NAND2_X1 i_0_1_173 (.A1(n_0_1_755), .A2(\aggregated_res[14] [63]), .ZN(
      n_0_1_754));
   NOR2_X1 i_0_1_174 (.A1(n_0_1_769), .A2(reset), .ZN(n_0_1_755));
   NAND2_X1 i_0_1_175 (.A1(n_0_1_769), .A2(n_0_1_837), .ZN(n_0_1_767));
   NOR2_X1 i_0_1_176 (.A1(n_0_1_773), .A2(n_0_1_908), .ZN(n_0_1_769));
   INV_X1 i_0_1_177 (.A(n_0_1_777), .ZN(n_0_1_773));
   NAND4_X1 i_0_1_178 (.A1(n_0_1_779), .A2(n_0_1_907), .A3(n_0_1_893), .A4(
      n_0_1_882), .ZN(n_0_1_777));
   NOR4_X1 i_0_1_179 (.A1(n_0_1_785), .A2(n_0_1_877), .A3(n_0_1_876), .A4(
      n_0_1_871), .ZN(n_0_1_779));
   NAND3_X1 i_0_1_180 (.A1(n_0_1_838), .A2(n_0_1_870), .A3(n_0_1_869), .ZN(
      n_0_1_785));
   INV_X1 i_0_1_181 (.A(\aggregated_res[14] [60]), .ZN(n_0_1_838));
   INV_X1 i_0_1_182 (.A(\aggregated_res[14] [61]), .ZN(n_0_1_869));
   INV_X1 i_0_1_183 (.A(\aggregated_res[14] [62]), .ZN(n_0_1_870));
   NAND4_X1 i_0_1_184 (.A1(n_0_1_875), .A2(n_0_1_874), .A3(n_0_1_873), .A4(
      n_0_1_872), .ZN(n_0_1_871));
   INV_X1 i_0_1_185 (.A(\aggregated_res[14] [10]), .ZN(n_0_1_872));
   INV_X1 i_0_1_186 (.A(\aggregated_res[14] [11]), .ZN(n_0_1_873));
   INV_X1 i_0_1_187 (.A(\aggregated_res[14] [12]), .ZN(n_0_1_874));
   INV_X1 i_0_1_188 (.A(\aggregated_res[14] [13]), .ZN(n_0_1_875));
   OR4_X1 i_0_1_189 (.A1(\aggregated_res[14] [54]), .A2(\aggregated_res[14] [53]), 
      .A3(\aggregated_res[14] [52]), .A4(\aggregated_res[14] [51]), .ZN(
      n_0_1_876));
   NAND4_X1 i_0_1_190 (.A1(n_0_1_880), .A2(n_0_1_881), .A3(n_0_1_879), .A4(
      n_0_1_878), .ZN(n_0_1_877));
   INV_X1 i_0_1_191 (.A(\aggregated_res[14] [55]), .ZN(n_0_1_878));
   INV_X1 i_0_1_192 (.A(\aggregated_res[14] [56]), .ZN(n_0_1_879));
   INV_X1 i_0_1_193 (.A(\aggregated_res[14] [57]), .ZN(n_0_1_880));
   INV_X1 i_0_1_194 (.A(\aggregated_res[14] [58]), .ZN(n_0_1_881));
   NOR3_X1 i_0_1_195 (.A1(n_0_1_888), .A2(\aggregated_res[14] [59]), .A3(
      n_0_1_883), .ZN(n_0_1_882));
   NAND4_X1 i_0_1_196 (.A1(n_0_1_887), .A2(n_0_1_886), .A3(n_0_1_885), .A4(
      n_0_1_884), .ZN(n_0_1_883));
   INV_X1 i_0_1_197 (.A(\aggregated_res[14] [14]), .ZN(n_0_1_884));
   INV_X1 i_0_1_198 (.A(\aggregated_res[14] [15]), .ZN(n_0_1_885));
   INV_X1 i_0_1_199 (.A(\aggregated_res[14] [31]), .ZN(n_0_1_886));
   INV_X1 i_0_1_200 (.A(\aggregated_res[14] [32]), .ZN(n_0_1_887));
   NAND4_X1 i_0_1_201 (.A1(n_0_1_891), .A2(n_0_1_890), .A3(n_0_1_892), .A4(
      n_0_1_889), .ZN(n_0_1_888));
   INV_X1 i_0_1_202 (.A(\aggregated_res[14] [47]), .ZN(n_0_1_889));
   INV_X1 i_0_1_203 (.A(\aggregated_res[14] [48]), .ZN(n_0_1_890));
   INV_X1 i_0_1_204 (.A(\aggregated_res[14] [49]), .ZN(n_0_1_891));
   INV_X1 i_0_1_205 (.A(\aggregated_res[14] [50]), .ZN(n_0_1_892));
   INV_X1 i_0_1_206 (.A(n_0_1_894), .ZN(n_0_1_893));
   OR4_X1 i_0_1_207 (.A1(n_0_1_902), .A2(n_0_1_896), .A3(n_0_1_897), .A4(
      n_0_1_895), .ZN(n_0_1_894));
   NAND4_X1 i_0_1_208 (.A1(n_0_1_80), .A2(n_0_1_77), .A3(n_0_1_74), .A4(n_0_1_81), 
      .ZN(n_0_1_895));
   NAND4_X1 i_0_1_209 (.A1(n_0_1_75), .A2(n_0_1_76), .A3(n_0_1_82), .A4(n_0_1_79), 
      .ZN(n_0_1_896));
   NAND4_X1 i_0_1_210 (.A1(n_0_1_901), .A2(n_0_1_900), .A3(n_0_1_899), .A4(
      n_0_1_898), .ZN(n_0_1_897));
   INV_X1 i_0_1_211 (.A(\aggregated_res[14] [6]), .ZN(n_0_1_898));
   INV_X1 i_0_1_212 (.A(\aggregated_res[14] [7]), .ZN(n_0_1_899));
   INV_X1 i_0_1_213 (.A(\aggregated_res[14] [8]), .ZN(n_0_1_900));
   INV_X1 i_0_1_214 (.A(\aggregated_res[14] [9]), .ZN(n_0_1_901));
   NAND4_X1 i_0_1_215 (.A1(n_0_1_906), .A2(n_0_1_905), .A3(n_0_1_904), .A4(
      n_0_1_903), .ZN(n_0_1_902));
   INV_X1 i_0_1_216 (.A(\aggregated_res[14] [2]), .ZN(n_0_1_903));
   INV_X1 i_0_1_217 (.A(\aggregated_res[14] [3]), .ZN(n_0_1_904));
   INV_X1 i_0_1_218 (.A(\aggregated_res[14] [4]), .ZN(n_0_1_905));
   INV_X1 i_0_1_219 (.A(\aggregated_res[14] [5]), .ZN(n_0_1_906));
   INV_X1 i_0_1_1044 (.A(n_0_813), .ZN(n_0_1_907));
   XNOR2_X1 i_0_1_1045 (.A(A_in), .B(B_in), .ZN(n_0_1_908));
   INV_X1 i_0_1_1046 (.A(n_0_124), .ZN(n_0_1_909));
   NAND2_X1 i_0_1_1047 (.A1(n_0_1_910), .A2(n_0_1_837), .ZN(n_0_283));
   NAND2_X1 i_0_1_1048 (.A1(enable), .A2(clk), .ZN(n_0_1_910));
   OAI211_X1 i_0_1_1049 (.A(n_0_1_912), .B(n_0_1_911), .C1(n_0_1_834), .C2(
      n_0_1_557), .ZN(n_0_677));
   NAND2_X1 i_0_1_1050 (.A1(A_imm[29]), .A2(n_0_1_558), .ZN(n_0_1_911));
   AOI22_X1 i_0_1_1051 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_559), .B1(
      A_imm_2s_complement[29]), .B2(n_0_1_556), .ZN(n_0_1_912));
   OAI211_X1 i_0_1_1104 (.A(n_0_1_913), .B(n_0_1_915), .C1(n_0_1_836), .C2(
      n_0_1_557), .ZN(n_0_678));
   AOI22_X1 i_0_1_1105 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_559), .B1(
      A_imm[30]), .B2(n_0_1_558), .ZN(n_0_1_913));
   INV_X1 i_0_1_1120 (.A(n_0_1_914), .ZN(n_0_1_559));
   NAND2_X1 i_0_1_1121 (.A1(n_0_1_560), .A2(n_0_1_566), .ZN(n_0_1_914));
   NOR2_X1 i_0_1_1124 (.A1(n_0_1_562), .A2(n_0_1_566), .ZN(n_0_1_558));
   NAND2_X1 i_0_1_1125 (.A1(n_0_1_560), .A2(n_0_1_565), .ZN(n_0_1_557));
   NAND2_X1 i_0_1_1126 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_556), .ZN(
      n_0_1_915));
   NOR3_X1 i_0_1_1127 (.A1(n_0_1_607), .A2(n_0_1_564), .A3(n_0_1_565), .ZN(
      n_0_1_556));
   OAI211_X1 i_0_1_1188 (.A(n_0_1_916), .B(n_0_1_917), .C1(n_0_1_818), .C2(
      n_0_1_600), .ZN(n_0_702));
   AOI22_X1 i_0_1_1189 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_602), .B1(
      A_imm[21]), .B2(n_0_1_601), .ZN(n_0_1_916));
   NAND2_X1 i_0_1_1196 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_599), .ZN(
      n_0_1_917));
   OAI211_X1 i_0_1_1197 (.A(n_0_1_919), .B(n_0_1_918), .C1(n_0_1_834), .C2(
      n_0_1_600), .ZN(n_0_710));
   NAND2_X1 i_0_1_1200 (.A1(A_imm[29]), .A2(n_0_1_601), .ZN(n_0_1_918));
   NOR2_X1 i_0_1_1201 (.A1(n_0_1_607), .A2(n_0_1_608), .ZN(n_0_1_601));
   NAND2_X1 i_0_1_1202 (.A1(n_0_1_606), .A2(n_0_1_603), .ZN(n_0_1_600));
   AOI22_X1 i_0_1_1203 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_602), .B1(
      A_imm_2s_complement[29]), .B2(n_0_1_599), .ZN(n_0_1_919));
   INV_X1 i_0_1_1264 (.A(n_0_1_920), .ZN(n_0_1_602));
   NAND2_X1 i_0_1_1265 (.A1(n_0_1_607), .A2(n_0_1_603), .ZN(n_0_1_920));
   INV_X1 i_0_1_1276 (.A(n_0_1_921), .ZN(n_0_1_599));
   OR3_X1 i_0_1_1277 (.A1(n_0_1_606), .A2(n_0_1_609), .A3(n_0_1_652), .ZN(
      n_0_1_921));
   OAI211_X1 i_0_1_1278 (.A(n_0_1_922), .B(n_0_1_923), .C1(n_0_1_826), .C2(
      n_0_1_643), .ZN(n_0_739));
   AOI22_X1 i_0_1_1279 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_645), .B1(
      A_imm[25]), .B2(n_0_1_644), .ZN(n_0_1_922));
   NAND2_X1 i_0_1_1300 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_642), .ZN(
      n_0_1_923));
   OAI211_X1 i_0_1_1301 (.A(n_0_1_925), .B(n_0_1_924), .C1(n_0_1_834), .C2(
      n_0_1_643), .ZN(n_0_743));
   NAND2_X1 i_0_1_1324 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_642), .ZN(
      n_0_1_924));
   NOR3_X1 i_0_1_1325 (.A1(n_0_1_693), .A2(n_0_1_650), .A3(n_0_1_651), .ZN(
      n_0_1_642));
   NAND2_X1 i_0_1_1332 (.A1(n_0_1_646), .A2(n_0_1_651), .ZN(n_0_1_643));
   AOI22_X1 i_0_1_1333 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_645), .B1(
      A_imm[29]), .B2(n_0_1_644), .ZN(n_0_1_925));
   INV_X1 i_0_1_1342 (.A(n_0_1_926), .ZN(n_0_1_645));
   NAND2_X1 i_0_1_1343 (.A1(n_0_1_646), .A2(n_0_1_652), .ZN(n_0_1_926));
   NOR2_X1 i_0_1_1344 (.A1(n_0_1_648), .A2(n_0_1_652), .ZN(n_0_1_644));
   OAI211_X1 i_0_1_1345 (.A(n_0_1_927), .B(n_0_1_929), .C1(n_0_1_826), .C2(
      n_0_1_686), .ZN(n_0_772));
   AOI22_X1 i_0_1_1348 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_688), .B1(
      A_imm[25]), .B2(n_0_1_687), .ZN(n_0_1_927));
   INV_X1 i_0_1_1349 (.A(n_0_1_928), .ZN(n_0_1_688));
   NAND2_X1 i_0_1_1350 (.A1(n_0_1_693), .A2(n_0_1_689), .ZN(n_0_1_928));
   NOR2_X1 i_0_1_1351 (.A1(n_0_1_693), .A2(n_0_1_694), .ZN(n_0_1_687));
   NAND2_X1 i_0_1_1352 (.A1(n_0_1_692), .A2(n_0_1_689), .ZN(n_0_1_686));
   NAND2_X1 i_0_1_1353 (.A1(A_imm_2s_complement[25]), .A2(n_0_1_685), .ZN(
      n_0_1_929));
   INV_X1 i_0_1_1354 (.A(n_0_1_930), .ZN(n_0_1_685));
   OR3_X1 i_0_1_1355 (.A1(n_0_1_692), .A2(n_0_1_695), .A3(n_0_1_736), .ZN(
      n_0_1_930));
   OAI211_X1 i_0_1_1364 (.A(n_0_1_931), .B(n_0_1_932), .C1(n_0_1_729), .C2(
      n_0_1_786), .ZN(n_0_785));
   AOI22_X1 i_0_1_1366 (.A1(A_imm_2s_complement[6]), .A2(n_0_1_731), .B1(
      A_imm[5]), .B2(n_0_1_730), .ZN(n_0_1_931));
   AOI21_X1 i_0_1_1386 (.A(n_0_1_787), .B1(n_0_5), .B2(A_in), .ZN(n_0_1_786));
   NAND2_X1 i_0_1_1387 (.A1(A_imm_2s_complement[5]), .A2(n_0_1_728), .ZN(
      n_0_1_932));
   OAI211_X1 i_0_1_1392 (.A(n_0_1_933), .B(n_0_1_934), .C1(n_0_1_729), .C2(
      n_0_1_810), .ZN(n_0_797));
   AOI22_X1 i_0_1_1393 (.A1(A_imm_2s_complement[18]), .A2(n_0_1_731), .B1(
      A_imm[17]), .B2(n_0_1_730), .ZN(n_0_1_933));
   AOI21_X1 i_0_1_1394 (.A(n_0_1_811), .B1(n_0_17), .B2(A_in), .ZN(n_0_1_810));
   NAND2_X1 i_0_1_1395 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_728), .ZN(
      n_0_1_934));
   OAI211_X1 i_0_1_1396 (.A(n_0_1_935), .B(n_0_1_936), .C1(n_0_1_729), .C2(
      n_0_1_818), .ZN(n_0_801));
   AOI22_X1 i_0_1_1397 (.A1(A_imm_2s_complement[22]), .A2(n_0_1_731), .B1(
      A_imm[21]), .B2(n_0_1_730), .ZN(n_0_1_935));
   AOI21_X1 i_0_1_1398 (.A(n_0_1_819), .B1(n_0_21), .B2(A_in), .ZN(n_0_1_818));
   NAND2_X1 i_0_1_1399 (.A1(A_imm_2s_complement[21]), .A2(n_0_1_728), .ZN(
      n_0_1_936));
   OAI211_X1 i_0_1_1422 (.A(n_0_1_937), .B(n_0_1_938), .C1(n_0_1_828), .C2(
      n_0_1_729), .ZN(n_0_806));
   AOI22_X1 i_0_1_1423 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_731), .B1(
      A_imm[26]), .B2(n_0_1_730), .ZN(n_0_1_937));
   NAND2_X1 i_0_1_1426 (.A1(A_imm_2s_complement[26]), .A2(n_0_1_728), .ZN(
      n_0_1_938));
   OAI211_X1 i_0_1_1427 (.A(n_0_1_939), .B(n_0_1_940), .C1(n_0_1_729), .C2(
      n_0_1_830), .ZN(n_0_807));
   AOI22_X1 i_0_1_1428 (.A1(A_imm_2s_complement[28]), .A2(n_0_1_731), .B1(
      A_imm[27]), .B2(n_0_1_730), .ZN(n_0_1_939));
   AOI21_X1 i_0_1_1429 (.A(n_0_1_831), .B1(n_0_27), .B2(A_in), .ZN(n_0_1_830));
   NAND2_X1 i_0_1_1430 (.A1(A_imm_2s_complement[27]), .A2(n_0_1_728), .ZN(
      n_0_1_940));
   OAI211_X1 i_0_1_1431 (.A(n_0_1_941), .B(n_0_1_942), .C1(n_0_1_834), .C2(
      n_0_1_729), .ZN(n_0_809));
   AOI22_X1 i_0_1_1432 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_731), .B1(
      A_imm[29]), .B2(n_0_1_730), .ZN(n_0_1_941));
   NAND2_X1 i_0_1_1434 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_728), .ZN(
      n_0_1_942));
   NAND4_X1 i_0_1_1435 (.A1(n_0_1_943), .A2(n_0_1_947), .A3(n_0_1_946), .A4(
      n_0_1_945), .ZN(n_0_810));
   NAND2_X1 i_0_1_1436 (.A1(A_imm_2s_complement[31]), .A2(n_0_1_731), .ZN(
      n_0_1_943));
   INV_X1 i_0_1_1437 (.A(n_0_1_944), .ZN(n_0_1_731));
   NAND2_X1 i_0_1_1438 (.A1(n_0_1_732), .A2(n_0_1_736), .ZN(n_0_1_944));
   OR2_X1 i_0_1_1439 (.A1(n_0_1_836), .A2(n_0_1_729), .ZN(n_0_1_945));
   NAND2_X1 i_0_1_1440 (.A1(n_0_1_732), .A2(n_0_1_735), .ZN(n_0_1_729));
   NAND2_X1 i_0_1_1447 (.A1(n_0_30), .A2(A_in), .ZN(n_0_1_836));
   NAND2_X1 i_0_1_1448 (.A1(A_imm[30]), .A2(n_0_1_730), .ZN(n_0_1_946));
   NOR2_X1 i_0_1_1449 (.A1(n_0_1_737), .A2(n_0_1_736), .ZN(n_0_1_730));
   NAND2_X1 i_0_1_1451 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_728), .ZN(
      n_0_1_947));
   INV_X1 i_0_1_1466 (.A(n_0_1_948), .ZN(n_0_1_728));
   OR3_X1 i_0_1_1475 (.A1(n_0_1_735), .A2(n_0_1_738), .A3(n_0_1_775), .ZN(
      n_0_1_948));
   NAND2_X1 i_0_1_1478 (.A1(n_0_1_739), .A2(n_0_1_949), .ZN(n_0_813));
   NAND2_X1 i_0_1_1481 (.A1(n_0_1_959), .A2(A_imm[1]), .ZN(n_0_1_949));
   OAI21_X1 i_0_1_1483 (.A(n_0_1_950), .B1(n_0_1_772), .B2(n_0_1_796), .ZN(
      n_0_823));
   AOI22_X1 i_0_1_1484 (.A1(A_imm_2s_complement[11]), .A2(n_0_1_770), .B1(
      A_imm_2s_complement[10]), .B2(n_0_1_771), .ZN(n_0_1_950));
   AOI21_X1 i_0_1_1487 (.A(n_0_1_797), .B1(n_0_10), .B2(A_in), .ZN(n_0_1_796));
   OAI21_X1 i_0_1_1495 (.A(n_0_1_951), .B1(n_0_1_772), .B2(n_0_1_802), .ZN(
      n_0_826));
   AOI22_X1 i_0_1_1499 (.A1(A_imm_2s_complement[14]), .A2(n_0_1_770), .B1(
      A_imm_2s_complement[13]), .B2(n_0_1_771), .ZN(n_0_1_951));
   AOI21_X1 i_0_1_1507 (.A(n_0_1_803), .B1(n_0_13), .B2(A_in), .ZN(n_0_1_802));
   OAI21_X1 i_0_1_1510 (.A(n_0_1_952), .B1(n_0_1_772), .B2(n_0_1_804), .ZN(
      n_0_827));
   AOI22_X1 i_0_1_1511 (.A1(A_imm_2s_complement[15]), .A2(n_0_1_770), .B1(
      A_imm_2s_complement[14]), .B2(n_0_1_771), .ZN(n_0_1_952));
   AOI21_X1 i_0_1_1513 (.A(n_0_1_805), .B1(n_0_14), .B2(A_in), .ZN(n_0_1_804));
   OAI21_X1 i_0_1_1514 (.A(n_0_1_953), .B1(n_0_1_772), .B2(n_0_1_806), .ZN(
      n_0_828));
   AOI22_X1 i_0_1_1517 (.A1(A_imm_2s_complement[16]), .A2(n_0_1_770), .B1(
      A_imm_2s_complement[15]), .B2(n_0_1_771), .ZN(n_0_1_953));
   AOI21_X1 i_0_1_1519 (.A(n_0_1_807), .B1(n_0_15), .B2(A_in), .ZN(n_0_1_806));
   OAI21_X1 i_0_1_1520 (.A(n_0_1_954), .B1(n_0_1_808), .B2(n_0_1_772), .ZN(
      n_0_829));
   AOI22_X1 i_0_1_1522 (.A1(A_imm_2s_complement[17]), .A2(n_0_1_770), .B1(
      A_imm_2s_complement[16]), .B2(n_0_1_771), .ZN(n_0_1_954));
   OAI21_X1 i_0_1_1523 (.A(n_0_1_955), .B1(n_0_1_832), .B2(n_0_1_772), .ZN(
      n_0_841));
   AOI22_X1 i_0_1_1526 (.A1(A_imm_2s_complement[29]), .A2(n_0_1_770), .B1(
      A_imm_2s_complement[28]), .B2(n_0_1_771), .ZN(n_0_1_955));
   INV_X1 i_0_1_1527 (.A(n_0_1_957), .ZN(n_0_1_770));
   OAI211_X1 i_0_1_1528 (.A(n_0_1_958), .B(n_0_1_956), .C1(n_0_1_964), .C2(
      n_0_1_957), .ZN(n_0_843));
   NAND2_X1 i_0_1_1559 (.A1(A_imm_2s_complement[30]), .A2(n_0_1_771), .ZN(
      n_0_1_956));
   NOR2_X1 i_0_1_1560 (.A1(n_0_1_774), .A2(n_0_186), .ZN(n_0_1_771));
   NAND2_X1 i_0_1_1561 (.A1(n_0_1_775), .A2(n_0_186), .ZN(n_0_1_957));
   OAI21_X1 i_0_1_1562 (.A(n_0_1_958), .B1(n_0_1_964), .B2(n_0_1_960), .ZN(
      n_0_844));
   NAND3_X1 i_0_1_1563 (.A1(n_0_30), .A2(A_in), .A3(n_0_1_959), .ZN(n_0_1_958));
   INV_X1 i_0_1_1564 (.A(n_0_1_772), .ZN(n_0_1_959));
   NAND2_X1 i_0_1_1565 (.A1(n_0_1_774), .A2(n_0_186), .ZN(n_0_1_772));
   INV_X1 i_0_1_1566 (.A(n_0_1_775), .ZN(n_0_1_960));
   OAI21_X1 i_0_1_1567 (.A(n_0_1_961), .B1(n_0_1_962), .B2(n_0_1_963), .ZN(
      n_0_1_775));
   NAND2_X1 i_0_1_1568 (.A1(n_0_1_963), .A2(n_0_185), .ZN(n_0_1_961));
   INV_X1 i_0_1_1569 (.A(n_0_31), .ZN(n_0_1_962));
   INV_X1 i_0_1_1570 (.A(B_in), .ZN(n_0_1_963));
   INV_X1 i_0_1_1571 (.A(A_imm_2s_complement[31]), .ZN(n_0_1_964));
   OAI21_X1 i_0_1_1572 (.A(n_0_1_965), .B1(n_0_1_966), .B2(n_0_1_969), .ZN(
      A_imm[1]));
   NAND2_X1 i_0_1_1573 (.A1(n_0_1_969), .A2(n_0_154), .ZN(n_0_1_965));
   INV_X1 i_0_1_1574 (.A(n_0_0), .ZN(n_0_1_966));
   INV_X1 i_0_1_1575 (.A(n_0_1_778), .ZN(A_imm[2]));
   AOI21_X1 i_0_1_1576 (.A(n_0_1_967), .B1(n_0_1), .B2(A_in), .ZN(n_0_1_778));
   NOR2_X1 i_0_1_1577 (.A1(A_in), .A2(n_0_1_839), .ZN(n_0_1_967));
   AOI21_X1 i_0_1_1578 (.A(n_0_1_968), .B1(n_0_1_969), .B2(n_0_1_842), .ZN(
      A_imm[5]));
   NOR2_X1 i_0_1_1579 (.A1(n_0_4), .A2(n_0_1_969), .ZN(n_0_1_968));
   INV_X1 i_0_1_1580 (.A(A_in), .ZN(n_0_1_969));
   INV_X1 i_0_1_1581 (.A(n_0_1_808), .ZN(A_imm[17]));
   AOI21_X1 i_0_1_1582 (.A(n_0_1_809), .B1(n_0_16), .B2(A_in), .ZN(n_0_1_808));
   INV_X1 i_0_1_1583 (.A(n_0_1_816), .ZN(A_imm[21]));
   INV_X1 i_0_1_1584 (.A(n_0_1_824), .ZN(A_imm[25]));
   INV_X1 i_0_1_1585 (.A(n_0_1_826), .ZN(A_imm[26]));
   AOI21_X1 i_0_1_1586 (.A(n_0_1_827), .B1(n_0_25), .B2(A_in), .ZN(n_0_1_826));
   INV_X1 i_0_1_1587 (.A(n_0_1_828), .ZN(A_imm[27]));
   AOI21_X1 i_0_1_1588 (.A(n_0_1_829), .B1(n_0_26), .B2(A_in), .ZN(n_0_1_828));
   INV_X1 i_0_1_1589 (.A(n_0_1_832), .ZN(A_imm[29]));
   AOI21_X1 i_0_1_1590 (.A(n_0_1_833), .B1(n_0_28), .B2(A_in), .ZN(n_0_1_832));
   INV_X1 i_0_1_1591 (.A(n_0_1_834), .ZN(A_imm[30]));
   AOI21_X1 i_0_1_1592 (.A(n_0_1_835), .B1(n_0_29), .B2(A_in), .ZN(n_0_1_834));
   INV_X1 i_0_1_1593 (.A(reset), .ZN(n_0_1_970));
   AND2_X1 i_0_1_1594 (.A1(B[0]), .A2(n_0_1_970), .ZN(n_0_251));
   AND2_X1 i_0_1_1595 (.A1(B[1]), .A2(n_0_1_970), .ZN(n_0_252));
   AND2_X1 i_0_1_1596 (.A1(B[2]), .A2(n_0_1_970), .ZN(n_0_253));
   AND2_X1 i_0_1_1597 (.A1(B[3]), .A2(n_0_1_970), .ZN(n_0_254));
   AND2_X1 i_0_1_1598 (.A1(B[4]), .A2(n_0_1_970), .ZN(n_0_255));
   AND2_X1 i_0_1_1599 (.A1(B[5]), .A2(n_0_1_970), .ZN(n_0_256));
   AND2_X1 i_0_1_1600 (.A1(B[6]), .A2(n_0_1_970), .ZN(n_0_257));
   AND2_X1 i_0_1_1601 (.A1(B[7]), .A2(n_0_1_970), .ZN(n_0_258));
   AND2_X1 i_0_1_1602 (.A1(B[8]), .A2(n_0_1_970), .ZN(n_0_259));
   AND2_X1 i_0_1_1603 (.A1(B[9]), .A2(n_0_1_970), .ZN(n_0_260));
   AND2_X1 i_0_1_1604 (.A1(B[10]), .A2(n_0_1_970), .ZN(n_0_261));
   AND2_X1 i_0_1_1605 (.A1(B[11]), .A2(n_0_1_970), .ZN(n_0_262));
   AND2_X1 i_0_1_1606 (.A1(B[12]), .A2(n_0_1_970), .ZN(n_0_263));
   AND2_X1 i_0_1_1607 (.A1(B[13]), .A2(n_0_1_970), .ZN(n_0_264));
   AND2_X1 i_0_1_1608 (.A1(B[14]), .A2(n_0_1_970), .ZN(n_0_265));
   AND2_X1 i_0_1_1609 (.A1(B[15]), .A2(n_0_1_970), .ZN(n_0_266));
   AND2_X1 i_0_1_1610 (.A1(B[16]), .A2(n_0_1_970), .ZN(n_0_267));
   AND2_X1 i_0_1_1611 (.A1(B[17]), .A2(n_0_1_970), .ZN(n_0_268));
   AND2_X1 i_0_1_1612 (.A1(B[18]), .A2(n_0_1_970), .ZN(n_0_269));
   AND2_X1 i_0_1_1613 (.A1(B[19]), .A2(n_0_1_970), .ZN(n_0_270));
   AND2_X1 i_0_1_1614 (.A1(B[20]), .A2(n_0_1_970), .ZN(n_0_271));
   AND2_X1 i_0_1_1615 (.A1(B[21]), .A2(n_0_1_970), .ZN(n_0_272));
   AND2_X1 i_0_1_1616 (.A1(B[22]), .A2(n_0_1_970), .ZN(n_0_273));
   AND2_X1 i_0_1_1617 (.A1(B[23]), .A2(n_0_1_970), .ZN(n_0_274));
   AND2_X1 i_0_1_1618 (.A1(B[24]), .A2(n_0_1_970), .ZN(n_0_275));
   AND2_X1 i_0_1_1619 (.A1(B[25]), .A2(n_0_1_970), .ZN(n_0_276));
   AND2_X1 i_0_1_1620 (.A1(B[26]), .A2(n_0_1_970), .ZN(n_0_277));
   AND2_X1 i_0_1_1621 (.A1(B[27]), .A2(n_0_1_970), .ZN(n_0_278));
   AND2_X1 i_0_1_1622 (.A1(B[28]), .A2(n_0_1_970), .ZN(n_0_279));
   AND2_X1 i_0_1_1623 (.A1(B[29]), .A2(n_0_1_970), .ZN(n_0_280));
   AND2_X1 i_0_1_1624 (.A1(B[30]), .A2(n_0_1_970), .ZN(n_0_281));
   AND2_X1 i_0_1_1625 (.A1(B[31]), .A2(n_0_1_970), .ZN(n_0_282));
   AND2_X1 i_0_1_1626 (.A1(A[0]), .A2(n_0_1_970), .ZN(n_0_284));
   AND2_X1 i_0_1_1627 (.A1(A[1]), .A2(n_0_1_970), .ZN(n_0_285));
   AND2_X1 i_0_1_1628 (.A1(A[2]), .A2(n_0_1_970), .ZN(n_0_286));
   AND2_X1 i_0_1_1629 (.A1(A[3]), .A2(n_0_1_970), .ZN(n_0_287));
   AND2_X1 i_0_1_1630 (.A1(A[4]), .A2(n_0_1_970), .ZN(n_0_288));
   AND2_X1 i_0_1_1631 (.A1(A[5]), .A2(n_0_1_970), .ZN(n_0_289));
   AND2_X1 i_0_1_1632 (.A1(A[6]), .A2(n_0_1_970), .ZN(n_0_290));
   AND2_X1 i_0_1_1633 (.A1(A[7]), .A2(n_0_1_970), .ZN(n_0_291));
   AND2_X1 i_0_1_1634 (.A1(A[8]), .A2(n_0_1_970), .ZN(n_0_292));
   AND2_X1 i_0_1_1635 (.A1(A[9]), .A2(n_0_1_970), .ZN(n_0_293));
   AND2_X1 i_0_1_1636 (.A1(A[10]), .A2(n_0_1_970), .ZN(n_0_294));
   AND2_X1 i_0_1_1637 (.A1(A[11]), .A2(n_0_1_970), .ZN(n_0_295));
   AND2_X1 i_0_1_1638 (.A1(A[12]), .A2(n_0_1_970), .ZN(n_0_296));
   AND2_X1 i_0_1_1639 (.A1(A[13]), .A2(n_0_1_970), .ZN(n_0_297));
   AND2_X1 i_0_1_1640 (.A1(A[14]), .A2(n_0_1_970), .ZN(n_0_298));
   AND2_X1 i_0_1_1641 (.A1(A[15]), .A2(n_0_1_970), .ZN(n_0_299));
   AND2_X1 i_0_1_1642 (.A1(A[16]), .A2(n_0_1_970), .ZN(n_0_300));
   AND2_X1 i_0_1_1643 (.A1(A[17]), .A2(n_0_1_970), .ZN(n_0_301));
   AND2_X1 i_0_1_1644 (.A1(A[18]), .A2(n_0_1_970), .ZN(n_0_302));
   AND2_X1 i_0_1_1645 (.A1(A[19]), .A2(n_0_1_970), .ZN(n_0_303));
   AND2_X1 i_0_1_1646 (.A1(A[20]), .A2(n_0_1_970), .ZN(n_0_304));
   AND2_X1 i_0_1_1647 (.A1(A[21]), .A2(n_0_1_970), .ZN(n_0_305));
   AND2_X1 i_0_1_1648 (.A1(A[22]), .A2(n_0_1_970), .ZN(n_0_306));
   AND2_X1 i_0_1_1649 (.A1(A[23]), .A2(n_0_1_970), .ZN(n_0_307));
   AND2_X1 i_0_1_1650 (.A1(A[24]), .A2(n_0_1_970), .ZN(n_0_308));
   AND2_X1 i_0_1_1651 (.A1(A[25]), .A2(n_0_1_970), .ZN(n_0_309));
   AND2_X1 i_0_1_1652 (.A1(A[26]), .A2(n_0_1_970), .ZN(n_0_310));
   AND2_X1 i_0_1_1653 (.A1(A[27]), .A2(n_0_1_970), .ZN(n_0_311));
   AND2_X1 i_0_1_1654 (.A1(A[28]), .A2(n_0_1_970), .ZN(n_0_312));
   AND2_X1 i_0_1_1655 (.A1(A[29]), .A2(n_0_1_970), .ZN(n_0_313));
   AND2_X1 i_0_1_1656 (.A1(A[30]), .A2(n_0_1_970), .ZN(n_0_314));
   AND2_X1 i_0_1_1657 (.A1(A[31]), .A2(n_0_1_970), .ZN(n_0_315));
   NAND2_X1 i_0_1_1658 (.A1(clk), .A2(n_0_1_970), .ZN(n_0_316));
   OR2_X1 i_0_1_1659 (.A1(A_in), .A2(Res[63]), .ZN(OVF));
   BUF_X1 i_0_1_1660 (.A(n_0_1_970), .Z(n_0_1_837));
endmodule
