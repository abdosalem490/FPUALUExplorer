
// 	Thu Dec 22 21:36:19 2022
//	vlsi
//	192.168.126.129

module datapath__0_68 (\aggregated_res[14] , p_0);

output [63:0] p_0;
input [63:0] \aggregated_res[14] ;
wire slo_n488;
wire spw_n829;
wire slo__xsl_n217;
wire slo__sro_n346;
wire slo__xsl_n166;
wire n_13;
wire n_10;
wire n_11;
wire n_8;
wire n_9;
wire n_5;
wire n_7;
wire n_3;
wire n_4;
wire n_6;
wire n_2;
wire n_32;
wire n_39;
wire n_15;
wire n_17;
wire n_47;
wire n_41;
wire n_45;
wire n_46;
wire n_53;
wire n_12;
wire n_43;
wire n_66;
wire n_58;
wire n_63;
wire n_65;
wire n_72;
wire n_68;
wire n_93;
wire n_77;
wire n_87;
wire n_81;
wire n_89;
wire n_86;
wire n_23;
wire n_92;
wire n_21;
wire n_22;
wire n_19;
wire n_20;
wire n_31;
wire n_18;
wire n_29;
wire n_30;
wire n_27;
wire n_28;
wire n_25;
wire slo__sro_n319;
wire n_78;
wire n_24;
wire n_80;
wire n_37;
wire n_98;
wire n_35;
wire n_36;
wire n_97;
wire n_34;
wire n_112;
wire n_107;
wire n_140;
wire n_130;
wire n_128;
wire n_83;
wire n_152;
wire n_151;
wire n_115;
wire n_180;
wire n_146;
wire n_177;
wire n_178;
wire n_176;
wire n_153;
wire n_181;
wire n_172;
wire n_169;
wire sgo__sro_n48;
wire n_0;
wire n_1;
wire n_14;
wire n_16;
wire n_33;
wire n_38;
wire n_40;
wire n_42;
wire n_44;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_60;
wire n_59;
wire n_61;
wire n_62;
wire n_67;
wire n_64;
wire n_69;
wire n_70;
wire n_71;
wire n_73;
wire n_74;
wire slo__mro_n131;
wire n_76;
wire n_79;
wire n_82;
wire n_84;
wire n_85;
wire n_88;
wire n_90;
wire n_91;
wire n_94;
wire n_95;
wire n_96;
wire n_105;
wire n_102;
wire n_104;
wire n_100;
wire n_99;
wire n_103;
wire n_106;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_113;
wire n_114;
wire n_116;
wire n_119;
wire n_118;
wire n_117;
wire n_121;
wire n_120;
wire n_122;
wire n_123;
wire slo__sro_n144;
wire n_125;
wire n_126;
wire n_127;
wire n_129;
wire n_131;
wire n_132;
wire n_134;
wire n_133;
wire n_135;
wire sgo__sro_n12;
wire n_137;
wire n_139;
wire n_138;
wire n_143;
wire n_142;
wire n_141;
wire n_144;
wire n_145;
wire n_149;
wire n_150;
wire n_147;
wire n_148;
wire n_155;
wire n_154;
wire n_157;
wire n_158;
wire n_164;
wire n_162;
wire n_159;
wire n_165;
wire n_163;
wire n_160;
wire n_161;
wire sgo__sro_n13;
wire n_168;
wire n_171;
wire n_170;
wire n_173;
wire n_174;
wire n_175;
wire n_179;
wire sgo__sro_n14;
wire sgo__sro_n49;
wire sgo__sro_n50;
wire sgo__sro_n51;
wire slo__sro_n145;
wire sgo__sro_n38;
wire sgo__sro_n39;
wire sgo__sro_n116;
wire slo__sro_n199;
wire slo__sro_n200;
wire slo__sro_n201;
wire slo__xsl_n218;
wire slo__sro_n276;
wire slo__sro_n277;
wire slo__sro_n278;
wire slo__sro_n320;
wire slo__sro_n321;
wire slo__sro_n322;
wire slo__sro_n347;
wire slo__n357;
wire slo__n427;


INV_X1 i_244 (.ZN (n_181), .A (\aggregated_res[14] [62] ));
INV_X1 i_243 (.ZN (n_180), .A (\aggregated_res[14] [61] ));
AND2_X1 i_242 (.ZN (n_179), .A1 (\aggregated_res[14] [63] ), .A2 (n_181));
NAND4_X1 i_241 (.ZN (n_178), .A1 (n_155), .A2 (n_180), .A3 (n_177), .A4 (n_179));
NOR2_X4 i_240 (.ZN (n_177), .A1 (n_170), .A2 (\aggregated_res[14] [60] ));
INV_X1 slo__sro_c305 (.ZN (slo__sro_n278), .A (\aggregated_res[14] [51] ));
NOR2_X1 i_238 (.ZN (n_175), .A1 (\aggregated_res[14] [61] ), .A2 (n_176));
INV_X1 slo__xsl_c266 (.ZN (slo__xsl_n218), .A (n_162));
NOR2_X1 i_236 (.ZN (n_174), .A1 (\aggregated_res[14] [60] ), .A2 (\aggregated_res[14] [59] ));
NAND3_X2 i_235 (.ZN (n_173), .A1 (n_164), .A2 (slo__xsl_n217), .A3 (n_174));
INV_X2 i_234 (.ZN (n_172), .A (n_173));
NOR2_X4 i_233 (.ZN (n_171), .A1 (n_161), .A2 (\aggregated_res[14] [59] ));
INV_X2 i_232 (.ZN (n_170), .A (n_171));
NAND2_X2 i_231 (.ZN (n_169), .A1 (n_155), .A2 (n_171));
NAND2_X1 i_230 (.ZN (n_168), .A1 (n_160), .A2 (\aggregated_res[14] [59] ));
NAND2_X1 i_229 (.ZN (p_0[59]), .A1 (n_169), .A2 (n_168));
NOR2_X2 sgo__sro_c15 (.ZN (sgo__sro_n14), .A1 (\aggregated_res[14] [32] ), .A2 (\aggregated_res[14] [34] ));
OR2_X2 i_227 (.ZN (n_165), .A1 (n_125), .A2 (n_132));
NOR2_X4 i_226 (.ZN (n_164), .A1 (n_165), .A2 (n_148));
NOR2_X1 slo__c374 (.ZN (slo__n357), .A1 (n_107), .A2 (n_116));
NOR2_X4 i_224 (.ZN (n_162), .A1 (n_163), .A2 (\aggregated_res[14] [58] ));
INV_X1 i_223 (.ZN (n_161), .A (n_162));
NAND2_X1 i_222 (.ZN (n_160), .A1 (n_164), .A2 (slo__xsl_n217));
OR3_X2 i_221 (.ZN (n_159), .A1 (n_165), .A2 (n_163), .A3 (n_148));
AOI22_X2 i_220 (.ZN (p_0[58]), .A1 (n_164), .A2 (slo__xsl_n217), .B1 (\aggregated_res[14] [58] ), .B2 (n_159));
NOR2_X1 i_219 (.ZN (n_158), .A1 (\aggregated_res[14] [56] ), .A2 (n_145));
AOI21_X1 i_218 (.ZN (n_157), .A (slo_n488), .B1 (n_155), .B2 (n_154));
AOI21_X1 i_217 (.ZN (p_0[57]), .A (n_157), .B1 (slo_n488), .B2 (n_158));
INV_X1 slo__c159 (.ZN (n_122), .A (slo__sro_n319));
INV_X4 i_215 (.ZN (n_155), .A (n_145));
INV_X1 i_214 (.ZN (n_154), .A (\aggregated_res[14] [56] ));
OAI22_X1 i_213 (.ZN (p_0[56]), .A1 (n_155), .A2 (\aggregated_res[14] [56] ), .B1 (n_145), .B2 (n_154));
INV_X1 i_212 (.ZN (n_150), .A (n_116));
INV_X1 i_211 (.ZN (n_149), .A (\aggregated_res[14] [55] ));
NAND4_X4 i_210 (.ZN (n_148), .A1 (n_149), .A2 (n_142), .A3 (n_143), .A4 (n_141));
INV_X2 i_209 (.ZN (n_147), .A (n_148));
AND3_X4 i_208 (.ZN (n_146), .A1 (n_134), .A2 (n_133), .A3 (n_147));
NAND3_X4 i_207 (.ZN (n_145), .A1 (n_146), .A2 (n_106), .A3 (n_150));
NOR2_X4 slo__c424 (.ZN (slo__n427), .A1 (n_90), .A2 (\aggregated_res[14] [31] ));
INV_X1 i_205 (.ZN (p_0[55]), .A (n_144));
INV_X1 i_204 (.ZN (n_143), .A (\aggregated_res[14] [54] ));
INV_X1 i_203 (.ZN (n_142), .A (\aggregated_res[14] [53] ));
INV_X1 i_202 (.ZN (n_141), .A (\aggregated_res[14] [52] ));
INV_X2 i_201 (.ZN (n_140), .A (n_137));
NOR4_X2 i_200 (.ZN (n_139), .A1 (n_130), .A2 (\aggregated_res[14] [52] ), .A3 (\aggregated_res[14] [53] ), .A4 (\aggregated_res[14] [54] ));
AOI21_X1 i_199 (.ZN (n_138), .A (n_143), .B1 (n_142), .B2 (n_140));
NOR2_X1 i_198 (.ZN (p_0[54]), .A1 (n_139), .A2 (n_138));
INV_X1 slo__sro_c249 (.ZN (slo__sro_n201), .A (\aggregated_res[14] [61] ));
OR4_X2 i_196 (.ZN (n_137), .A1 (n_135), .A2 (n_132), .A3 (\aggregated_res[14] [52] ), .A4 (n_117));
INV_X1 slo__xsl_c211 (.ZN (slo__xsl_n166), .A (n_27));
NAND4_X1 i_194 (.ZN (n_135), .A1 (n_99), .A2 (n_108), .A3 (n_94), .A4 (n_119));
INV_X1 i_193 (.ZN (n_134), .A (\aggregated_res[14] [49] ));
NOR2_X1 slo__sro_c339 (.ZN (slo__sro_n321), .A1 (\aggregated_res[14] [38] ), .A2 (\aggregated_res[14] [39] ));
NAND2_X1 i_191 (.ZN (n_132), .A1 (n_134), .A2 (n_133));
INV_X1 i_190 (.ZN (n_131), .A (n_132));
NAND2_X2 i_189 (.ZN (n_130), .A1 (slo__n357), .A2 (n_131));
OAI21_X1 i_188 (.ZN (n_129), .A (\aggregated_res[14] [51] ), .B1 (\aggregated_res[14] [50] ), .B2 (n_126));
AND2_X1 i_187 (.ZN (p_0[51]), .A1 (n_130), .A2 (n_129));
XOR2_X1 i_186 (.Z (p_0[50]), .A (n_126), .B (\aggregated_res[14] [50] ));
NAND2_X1 i_185 (.ZN (n_128), .A1 (n_126), .A2 (n_127));
NAND2_X1 i_184 (.ZN (n_127), .A1 (n_120), .A2 (\aggregated_res[14] [49] ));
OR3_X1 i_183 (.ZN (n_126), .A1 (n_125), .A2 (\aggregated_res[14] [48] ), .A3 (\aggregated_res[14] [49] ));
NAND4_X2 i_182 (.ZN (n_125), .A1 (sgo__sro_n48), .A2 (n_109), .A3 (n_118), .A4 (n_103));
NOR2_X4 slo__sro_c184 (.ZN (slo__sro_n145), .A1 (\aggregated_res[14] [24] ), .A2 (\aggregated_res[14] [22] ));
NAND2_X2 i_180 (.ZN (n_123), .A1 (slo__n427), .A2 (sgo__sro_n12));
INV_X1 slo__mro_c169 (.ZN (slo__mro_n131), .A (\aggregated_res[14] [53] ));
INV_X1 i_178 (.ZN (n_121), .A (spw_n829));
NAND2_X1 i_177 (.ZN (n_120), .A1 (n_121), .A2 (n_115));
AOI22_X1 i_176 (.ZN (p_0[48]), .A1 (n_121), .A2 (n_115), .B1 (spw_n829), .B2 (n_114));
INV_X1 i_175 (.ZN (n_119), .A (\aggregated_res[14] [45] ));
NOR2_X1 i_174 (.ZN (n_118), .A1 (\aggregated_res[14] [47] ), .A2 (\aggregated_res[14] [46] ));
INV_X1 i_173 (.ZN (n_117), .A (n_118));
NAND2_X1 i_172 (.ZN (n_116), .A1 (n_119), .A2 (n_118));
NOR2_X1 i_171 (.ZN (n_115), .A1 (n_107), .A2 (n_116));
INV_X1 i_170 (.ZN (n_114), .A (n_115));
AOI21_X1 i_169 (.ZN (p_0[47]), .A (n_115), .B1 (\aggregated_res[14] [47] ), .B2 (n_111));
INV_X1 i_168 (.ZN (n_113), .A (\aggregated_res[14] [46] ));
NOR2_X1 i_167 (.ZN (n_112), .A1 (\aggregated_res[14] [45] ), .A2 (n_107));
NAND2_X1 i_166 (.ZN (n_111), .A1 (n_113), .A2 (n_112));
OAI21_X1 i_165 (.ZN (n_110), .A (n_111), .B1 (n_113), .B2 (n_112));
INV_X1 i_164 (.ZN (p_0[46]), .A (n_110));
INV_X1 i_163 (.ZN (n_109), .A (\aggregated_res[14] [44] ));
AND2_X2 i_162 (.ZN (n_108), .A1 (n_109), .A2 (n_103));
NAND3_X4 i_161 (.ZN (n_107), .A1 (n_99), .A2 (n_108), .A3 (n_94));
INV_X2 i_160 (.ZN (n_106), .A (n_107));
AOI21_X1 i_159 (.ZN (p_0[44]), .A (n_106), .B1 (\aggregated_res[14] [44] ), .B2 (n_96));
INV_X1 i_158 (.ZN (n_105), .A (\aggregated_res[14] [43] ));
INV_X1 i_157 (.ZN (n_104), .A (\aggregated_res[14] [36] ));
NOR3_X2 i_156 (.ZN (n_103), .A1 (\aggregated_res[14] [41] ), .A2 (\aggregated_res[14] [40] ), .A3 (\aggregated_res[14] [42] ));
INV_X1 i_155 (.ZN (n_102), .A (n_103));
INV_X2 sgo__sro_c66 (.ZN (sgo__sro_n51), .A (n_123));
NOR3_X1 i_153 (.ZN (n_100), .A1 (\aggregated_res[14] [37] ), .A2 (\aggregated_res[14] [38] ), .A3 (\aggregated_res[14] [39] ));
AND2_X4 sgo__sro_c143 (.ZN (sgo__sro_n116), .A1 (n_146), .A2 (n_150));
NAND4_X1 i_151 (.ZN (n_98), .A1 (n_104), .A2 (n_100), .A3 (sgo__sro_n12), .A4 (n_94));
NOR2_X1 i_150 (.ZN (n_97), .A1 (n_102), .A2 (n_98));
NAND2_X1 i_149 (.ZN (n_96), .A1 (n_105), .A2 (n_97));
OAI21_X1 i_148 (.ZN (n_95), .A (n_96), .B1 (n_105), .B2 (n_97));
INV_X1 i_147 (.ZN (p_0[43]), .A (n_95));
NOR2_X4 i_146 (.ZN (n_94), .A1 (n_90), .A2 (\aggregated_res[14] [31] ));
INV_X1 i_145 (.ZN (n_92), .A (slo__n427));
AOI21_X1 i_144 (.ZN (p_0[31]), .A (n_94), .B1 (n_90), .B2 (\aggregated_res[14] [31] ));
NOR2_X2 i_143 (.ZN (n_91), .A1 (\aggregated_res[14] [30] ), .A2 (\aggregated_res[14] [28] ));
NAND3_X4 i_142 (.ZN (n_90), .A1 (n_82), .A2 (n_88), .A3 (n_91));
INV_X1 i_141 (.ZN (n_89), .A (n_90));
INV_X4 i_140 (.ZN (n_88), .A (\aggregated_res[14] [29] ));
NOR2_X1 i_139 (.ZN (n_87), .A1 (n_81), .A2 (\aggregated_res[14] [28] ));
NAND2_X1 i_138 (.ZN (n_86), .A1 (n_88), .A2 (n_87));
OAI21_X1 i_137 (.ZN (n_85), .A (n_86), .B1 (n_88), .B2 (n_87));
INV_X1 i_136 (.ZN (p_0[29]), .A (n_85));
INV_X1 i_135 (.ZN (n_84), .A (\aggregated_res[14] [26] ));
NAND3_X4 i_134 (.ZN (n_83), .A1 (n_74), .A2 (n_79), .A3 (n_84));
NOR2_X4 i_133 (.ZN (n_82), .A1 (n_83), .A2 (\aggregated_res[14] [27] ));
INV_X1 i_132 (.ZN (n_81), .A (n_82));
AOI21_X1 i_131 (.ZN (p_0[27]), .A (n_82), .B1 (\aggregated_res[14] [27] ), .B2 (n_83));
INV_X2 i_130 (.ZN (n_79), .A (\aggregated_res[14] [25] ));
NAND2_X1 i_129 (.ZN (n_77), .A1 (n_79), .A2 (n_74));
OAI21_X1 i_128 (.ZN (n_76), .A (n_77), .B1 (n_79), .B2 (n_74));
INV_X1 i_127 (.ZN (p_0[25]), .A (n_76));
XNOR2_X2 slo__mro_c170 (.ZN (p_0[53]), .A (n_137), .B (slo__mro_n131));
OR2_X2 slo__xsl_c214 (.ZN (n_27), .A1 (\aggregated_res[14] [37] ), .A2 (n_28));
AOI21_X1 i_124 (.ZN (p_0[24]), .A (n_74), .B1 (\aggregated_res[14] [24] ), .B2 (n_71));
INV_X1 i_123 (.ZN (n_73), .A (\aggregated_res[14] [23] ));
NOR2_X1 i_122 (.ZN (n_72), .A1 (n_68), .A2 (\aggregated_res[14] [22] ));
NAND2_X1 i_121 (.ZN (n_71), .A1 (n_73), .A2 (n_72));
OAI21_X1 i_120 (.ZN (n_70), .A (n_71), .B1 (n_73), .B2 (n_72));
INV_X1 i_119 (.ZN (p_0[23]), .A (n_70));
NOR3_X4 i_118 (.ZN (n_69), .A1 (\aggregated_res[14] [21] ), .A2 (n_58), .A3 (\aggregated_res[14] [18] ));
NAND2_X2 i_117 (.ZN (n_68), .A1 (n_64), .A2 (n_69));
AOI22_X1 i_116 (.ZN (p_0[21]), .A1 (n_64), .A2 (n_69), .B1 (\aggregated_res[14] [21] ), .B2 (n_62));
INV_X1 i_115 (.ZN (n_67), .A (\aggregated_res[14] [20] ));
NOR2_X1 i_114 (.ZN (n_66), .A1 (n_58), .A2 (\aggregated_res[14] [18] ));
INV_X1 i_113 (.ZN (n_65), .A (n_66));
NOR2_X4 i_112 (.ZN (n_64), .A1 (\aggregated_res[14] [20] ), .A2 (\aggregated_res[14] [19] ));
NOR2_X1 i_111 (.ZN (n_63), .A1 (\aggregated_res[14] [19] ), .A2 (n_65));
NAND2_X1 i_110 (.ZN (n_62), .A1 (n_67), .A2 (n_63));
OAI21_X1 i_109 (.ZN (n_61), .A (n_62), .B1 (n_67), .B2 (n_63));
INV_X1 i_108 (.ZN (p_0[20]), .A (n_61));
INV_X1 i_107 (.ZN (n_60), .A (\aggregated_res[14] [17] ));
NOR2_X1 i_106 (.ZN (n_59), .A1 (n_54), .A2 (n_41));
NAND3_X2 i_105 (.ZN (n_58), .A1 (n_60), .A2 (n_59), .A3 (n_56));
OAI21_X1 i_104 (.ZN (n_57), .A (n_58), .B1 (n_60), .B2 (n_51));
INV_X1 i_103 (.ZN (p_0[17]), .A (n_57));
INV_X1 i_102 (.ZN (n_56), .A (\aggregated_res[14] [16] ));
INV_X1 i_101 (.ZN (n_55), .A (\aggregated_res[14] [15] ));
NAND4_X1 i_100 (.ZN (n_54), .A1 (n_55), .A2 (n_50), .A3 (n_49), .A4 (n_48));
NOR2_X1 i_99 (.ZN (n_53), .A1 (n_41), .A2 (n_54));
INV_X1 i_98 (.ZN (n_52), .A (n_53));
NOR2_X1 i_97 (.ZN (n_51), .A1 (\aggregated_res[14] [16] ), .A2 (n_52));
AOI21_X1 i_96 (.ZN (p_0[16]), .A (n_51), .B1 (\aggregated_res[14] [16] ), .B2 (n_52));
INV_X1 i_95 (.ZN (n_50), .A (\aggregated_res[14] [14] ));
INV_X1 i_94 (.ZN (n_49), .A (\aggregated_res[14] [13] ));
INV_X1 i_93 (.ZN (n_48), .A (\aggregated_res[14] [12] ));
NOR2_X1 i_92 (.ZN (n_47), .A1 (\aggregated_res[14] [12] ), .A2 (n_41));
INV_X1 i_91 (.ZN (n_46), .A (n_47));
NOR2_X1 i_90 (.ZN (n_45), .A1 (\aggregated_res[14] [13] ), .A2 (n_46));
INV_X1 i_89 (.ZN (n_44), .A (n_45));
NOR2_X1 i_88 (.ZN (n_43), .A1 (\aggregated_res[14] [14] ), .A2 (n_44));
AOI21_X1 i_87 (.ZN (p_0[14]), .A (n_43), .B1 (\aggregated_res[14] [14] ), .B2 (n_44));
INV_X1 i_86 (.ZN (n_42), .A (\aggregated_res[14] [11] ));
NAND4_X1 i_85 (.ZN (n_41), .A1 (n_0), .A2 (n_38), .A3 (n_33), .A4 (n_42));
OAI21_X1 i_84 (.ZN (n_40), .A (n_41), .B1 (n_42), .B2 (n_14));
INV_X1 i_83 (.ZN (p_0[11]), .A (n_40));
INV_X1 i_81 (.ZN (n_39), .A (n_0));
INV_X1 i_80 (.ZN (n_38), .A (\aggregated_res[14] [10] ));
NOR2_X1 i_79 (.ZN (n_33), .A1 (\aggregated_res[14] [9] ), .A2 (\aggregated_res[14] [8] ));
NOR2_X1 i_78 (.ZN (n_32), .A1 (n_39), .A2 (\aggregated_res[14] [8] ));
INV_X1 i_77 (.ZN (n_17), .A (n_32));
NAND2_X1 i_76 (.ZN (n_16), .A1 (n_0), .A2 (n_33));
INV_X1 i_75 (.ZN (n_15), .A (n_16));
NOR2_X1 i_74 (.ZN (n_14), .A1 (\aggregated_res[14] [10] ), .A2 (n_16));
AOI21_X1 i_73 (.ZN (p_0[10]), .A (n_14), .B1 (\aggregated_res[14] [10] ), .B2 (n_16));
NOR2_X1 i_72 (.ZN (n_13), .A1 (\aggregated_res[14] [1] ), .A2 (\aggregated_res[14] [0] ));
INV_X1 i_71 (.ZN (n_11), .A (n_13));
NOR2_X1 i_70 (.ZN (n_10), .A1 (\aggregated_res[14] [2] ), .A2 (n_11));
INV_X1 i_69 (.ZN (n_9), .A (n_10));
NOR2_X1 i_68 (.ZN (n_8), .A1 (\aggregated_res[14] [3] ), .A2 (n_9));
INV_X1 i_67 (.ZN (n_7), .A (n_8));
NOR4_X1 i_66 (.ZN (n_6), .A1 (\aggregated_res[14] [6] ), .A2 (\aggregated_res[14] [5] )
    , .A3 (\aggregated_res[14] [4] ), .A4 (n_7));
INV_X1 i_65 (.ZN (n_1), .A (n_6));
NOR2_X1 i_64 (.ZN (n_0), .A1 (\aggregated_res[14] [7] ), .A2 (n_1));
AOI21_X1 i_63 (.ZN (p_0[7]), .A (n_0), .B1 (\aggregated_res[14] [7] ), .B2 (n_1));
INV_X1 i_62 (.ZN (n_80), .A (sgo__sro_n12));
AOI21_X1 i_61 (.ZN (p_0[60]), .A (n_172), .B1 (n_169), .B2 (\aggregated_res[14] [60] ));
NAND2_X1 i_60 (.ZN (n_153), .A1 (n_181), .A2 (n_180));
NOR2_X4 i_59 (.ZN (n_152), .A1 (n_176), .A2 (n_153));
OAI21_X1 i_58 (.ZN (p_0[63]), .A (n_178), .B1 (n_152), .B2 (\aggregated_res[14] [63] ));
NAND4_X1 i_57 (.ZN (n_151), .A1 (n_115), .A2 (n_180), .A3 (n_146), .A4 (n_177));
AOI21_X1 i_56 (.ZN (p_0[62]), .A (n_152), .B1 (n_151), .B2 (\aggregated_res[14] [62] ));
INV_X1 i_55 (.ZN (n_93), .A (n_83));
INV_X1 slo__sro_c361 (.ZN (slo__sro_n347), .A (\aggregated_res[14] [57] ));
INV_X1 i_53 (.ZN (p_0[49]), .A (n_128));
INV_X1 i_52 (.ZN (n_78), .A (n_98));
AOI21_X1 i_48 (.ZN (p_0[52]), .A (n_140), .B1 (\aggregated_res[14] [52] ), .B2 (n_130));
AOI21_X1 i_82 (.ZN (p_0[45]), .A (n_112), .B1 (\aggregated_res[14] [45] ), .B2 (n_107));
NOR2_X1 i_47 (.ZN (n_37), .A1 (\aggregated_res[14] [40] ), .A2 (n_98));
INV_X1 i_46 (.ZN (n_36), .A (n_37));
NOR2_X1 i_44 (.ZN (n_35), .A1 (\aggregated_res[14] [41] ), .A2 (n_36));
INV_X1 i_43 (.ZN (n_34), .A (n_35));
AOI21_X1 i_42 (.ZN (p_0[42]), .A (n_97), .B1 (\aggregated_res[14] [42] ), .B2 (n_34));
AOI21_X1 i_41 (.ZN (p_0[41]), .A (n_35), .B1 (\aggregated_res[14] [41] ), .B2 (n_36));
AOI21_X1 i_40 (.ZN (p_0[40]), .A (n_37), .B1 (\aggregated_res[14] [40] ), .B2 (n_98));
NOR2_X2 i_38 (.ZN (n_31), .A1 (n_92), .A2 (n_80));
INV_X1 i_37 (.ZN (n_30), .A (n_31));
NOR2_X2 i_35 (.ZN (n_29), .A1 (\aggregated_res[14] [36] ), .A2 (n_30));
INV_X1 i_34 (.ZN (n_28), .A (n_29));
INV_X1 slo__sro_c250 (.ZN (slo__sro_n200), .A (n_173));
INV_X1 slo__sro_c338 (.ZN (slo__sro_n322), .A (\aggregated_res[14] [43] ));
NOR2_X2 i_31 (.ZN (n_25), .A1 (\aggregated_res[14] [38] ), .A2 (n_27));
INV_X1 i_30 (.ZN (n_24), .A (n_25));
AOI21_X1 i_29 (.ZN (p_0[39]), .A (n_78), .B1 (\aggregated_res[14] [39] ), .B2 (n_24));
AOI21_X1 i_28 (.ZN (p_0[38]), .A (n_25), .B1 (\aggregated_res[14] [38] ), .B2 (n_27));
AOI21_X1 i_27 (.ZN (p_0[37]), .A (slo__xsl_n166), .B1 (\aggregated_res[14] [37] ), .B2 (n_28));
AOI21_X1 i_26 (.ZN (p_0[36]), .A (n_29), .B1 (\aggregated_res[14] [36] ), .B2 (n_30));
NOR2_X1 i_25 (.ZN (n_23), .A1 (\aggregated_res[14] [32] ), .A2 (n_92));
INV_X1 i_22 (.ZN (n_22), .A (n_23));
NOR2_X1 i_21 (.ZN (n_21), .A1 (\aggregated_res[14] [33] ), .A2 (n_22));
INV_X1 i_20 (.ZN (n_20), .A (n_21));
NOR2_X1 i_19 (.ZN (n_19), .A1 (\aggregated_res[14] [34] ), .A2 (n_20));
INV_X1 i_18 (.ZN (n_18), .A (n_19));
AOI21_X1 i_17 (.ZN (p_0[35]), .A (n_31), .B1 (\aggregated_res[14] [35] ), .B2 (n_18));
AOI21_X1 i_51 (.ZN (p_0[34]), .A (n_19), .B1 (\aggregated_res[14] [34] ), .B2 (n_20));
AOI21_X1 i_50 (.ZN (p_0[33]), .A (n_21), .B1 (\aggregated_res[14] [33] ), .B2 (n_22));
AOI21_X1 i_49 (.ZN (p_0[32]), .A (n_23), .B1 (\aggregated_res[14] [32] ), .B2 (n_92));
AOI21_X1 i_16 (.ZN (p_0[30]), .A (n_89), .B1 (\aggregated_res[14] [30] ), .B2 (n_86));
AOI21_X1 i_45 (.ZN (p_0[28]), .A (n_87), .B1 (\aggregated_res[14] [28] ), .B2 (n_81));
AOI21_X1 i_15 (.ZN (p_0[26]), .A (n_93), .B1 (\aggregated_res[14] [26] ), .B2 (n_77));
AOI21_X1 i_39 (.ZN (p_0[22]), .A (n_72), .B1 (\aggregated_res[14] [22] ), .B2 (n_68));
AOI21_X1 i_36 (.ZN (p_0[19]), .A (n_63), .B1 (\aggregated_res[14] [19] ), .B2 (n_65));
AOI21_X1 i_14 (.ZN (p_0[18]), .A (n_66), .B1 (\aggregated_res[14] [18] ), .B2 (n_58));
INV_X1 i_13 (.ZN (n_12), .A (n_43));
AOI21_X1 i_12 (.ZN (p_0[15]), .A (n_53), .B1 (\aggregated_res[14] [15] ), .B2 (n_12));
AOI21_X1 i_24 (.ZN (p_0[13]), .A (n_45), .B1 (\aggregated_res[14] [13] ), .B2 (n_46));
AOI21_X1 i_23 (.ZN (p_0[12]), .A (n_47), .B1 (\aggregated_res[14] [12] ), .B2 (n_41));
AOI21_X1 i_11 (.ZN (p_0[9]), .A (n_15), .B1 (\aggregated_res[14] [9] ), .B2 (n_17));
AOI21_X1 i_10 (.ZN (p_0[8]), .A (n_32), .B1 (\aggregated_res[14] [8] ), .B2 (n_39));
NOR2_X1 i_9 (.ZN (n_5), .A1 (\aggregated_res[14] [4] ), .A2 (n_7));
INV_X1 i_8 (.ZN (n_4), .A (n_5));
NOR2_X1 i_7 (.ZN (n_3), .A1 (\aggregated_res[14] [5] ), .A2 (n_4));
INV_X1 i_6 (.ZN (n_2), .A (n_3));
AOI21_X1 i_5 (.ZN (p_0[6]), .A (n_6), .B1 (\aggregated_res[14] [6] ), .B2 (n_2));
AOI21_X1 i_4 (.ZN (p_0[5]), .A (n_3), .B1 (\aggregated_res[14] [5] ), .B2 (n_4));
AOI21_X1 i_3 (.ZN (p_0[4]), .A (n_5), .B1 (\aggregated_res[14] [4] ), .B2 (n_7));
AOI21_X1 i_2 (.ZN (p_0[3]), .A (n_8), .B1 (\aggregated_res[14] [3] ), .B2 (n_9));
AOI21_X1 i_1 (.ZN (p_0[2]), .A (n_10), .B1 (\aggregated_res[14] [2] ), .B2 (n_11));
AOI21_X1 i_0 (.ZN (p_0[1]), .A (n_13), .B1 (\aggregated_res[14] [1] ), .B2 (\aggregated_res[14] [0] ));
NOR2_X2 sgo__sro_c16 (.ZN (sgo__sro_n13), .A1 (\aggregated_res[14] [33] ), .A2 (\aggregated_res[14] [35] ));
AND2_X4 sgo__sro_c17 (.ZN (sgo__sro_n12), .A1 (sgo__sro_n13), .A2 (sgo__sro_n14));
NOR2_X1 sgo__sro_c67 (.ZN (sgo__sro_n50), .A1 (\aggregated_res[14] [36] ), .A2 (\aggregated_res[14] [37] ));
NAND2_X2 sgo__sro_c68 (.ZN (sgo__sro_n49), .A1 (sgo__sro_n51), .A2 (sgo__sro_n50));
NOR2_X2 sgo__sro_c69 (.ZN (sgo__sro_n48), .A1 (n_122), .A2 (sgo__sro_n49));
NOR2_X2 slo__sro_c185 (.ZN (slo__sro_n144), .A1 (n_68), .A2 (\aggregated_res[14] [23] ));
AND2_X4 slo__sro_c186 (.ZN (n_74), .A1 (slo__sro_n145), .A2 (slo__sro_n144));
NOR2_X1 slo__sro_c251 (.ZN (slo__sro_n199), .A1 (slo__sro_n200), .A2 (slo__sro_n201));
NOR2_X1 slo__sro_c252 (.ZN (p_0[61]), .A1 (n_175), .A2 (slo__sro_n199));
INV_X1 slo__xsl_c267 (.ZN (slo__xsl_n217), .A (slo__xsl_n218));
NAND3_X2 sgo__sro_c49 (.ZN (sgo__sro_n39), .A1 (sgo__sro_n12), .A2 (n_104), .A3 (n_105));
INV_X1 sgo__sro_c50 (.ZN (sgo__sro_n38), .A (sgo__sro_n39));
AND2_X2 sgo__sro_c51 (.ZN (n_99), .A1 (sgo__sro_n38), .A2 (n_100));
NAND3_X4 sgo__sro_c144 (.ZN (n_176), .A1 (n_177), .A2 (n_106), .A3 (sgo__sro_n116));
INV_X1 slo__sro_c306 (.ZN (slo__sro_n277), .A (\aggregated_res[14] [50] ));
NAND2_X1 slo__sro_c307 (.ZN (slo__sro_n276), .A1 (slo__sro_n278), .A2 (slo__sro_n277));
NOR2_X1 slo__sro_c308 (.ZN (n_133), .A1 (\aggregated_res[14] [48] ), .A2 (slo__sro_n276));
NAND2_X1 slo__sro_c340 (.ZN (slo__sro_n320), .A1 (slo__sro_n321), .A2 (slo__sro_n322));
NOR2_X1 slo__sro_c341 (.ZN (slo__sro_n319), .A1 (\aggregated_res[14] [45] ), .A2 (slo__sro_n320));
INV_X1 slo__sro_c362 (.ZN (slo__sro_n346), .A (\aggregated_res[14] [56] ));
NAND2_X2 slo__sro_c363 (.ZN (n_163), .A1 (slo__sro_n346), .A2 (slo__sro_n347));
OAI21_X1 slo__sro_c379 (.ZN (n_144), .A (n_145), .B1 (n_139), .B2 (n_149));
CLKBUF_X1 slo___L1_c1_c461 (.Z (slo_n488), .A (\aggregated_res[14] [57] ));
CLKBUF_X1 spw__L1_c1_c829 (.Z (spw_n829), .A (\aggregated_res[14] [48] ));

endmodule //datapath__0_68

module datapath__0_67 (p_0, p_1, p_2, p_3, p_4, p_5, p_6, p_7, p_8, p_9, p_10, p_11, 
    p_12, p_13, p_14, p_15, \aggregated_res[14] );

output [63:0] \aggregated_res[14] ;
input [63:0] p_0;
input [63:0] p_10;
input [63:0] p_11;
input [63:0] p_12;
input [63:0] p_13;
input [63:0] p_14;
input [63:0] p_15;
input [63:0] p_1;
input [63:0] p_2;
input [63:0] p_3;
input [63:0] p_4;
input [63:0] p_5;
input [63:0] p_6;
input [63:0] p_7;
input [63:0] p_8;
input [63:0] p_9;
wire slo__sro_n1181;
wire slo__xsl_n395;
wire slo___n509;
wire slo__sro_n1107;
wire slo__sro_n460;
wire slo__n651;
wire CLOCK_slo__sro_n2895;
wire n_1175;
wire n_1315;
wire n_16;
wire n_912;
wire n_97;
wire n_913;
wire n_96;
wire n_81;
wire n_914;
wire n_99;
wire n_38;
wire n_77;
wire n_915;
wire n_49;
wire n_25;
wire n_73;
wire n_922;
wire n_69;
wire n_918;
wire n_105;
wire n_31;
wire n_29;
wire n_71;
wire n_23;
wire n_27;
wire n_273;
wire n_926;
wire n_271;
wire n_145;
wire n_185;
wire n_417;
wire n_932;
wire n_525;
wire n_418;
wire n_947;
wire n_941;
wire n_453;
wire n_1137;
wire n_943;
wire n_543;
wire n_447;
wire n_455;
wire n_953;
wire n_950;
wire n_951;
wire n_948;
wire n_659;
wire n_649;
wire n_955;
wire slo__n539;
wire n_657;
wire n_655;
wire n_1121;
wire n_952;
wire n_653;
wire n_636;
wire n_511;
wire n_507;
wire n_661;
wire n_555;
wire slo__sro_n704;
wire n_961;
wire n_958;
wire n_959;
wire n_956;
wire n_752;
wire n_1131;
wire n_1160;
wire n_983;
wire n_984;
wire n_981;
wire n_944;
wire n_1000;
wire n_896;
wire n_938;
wire sgo__sro_n18;
wire n_992;
wire n_991;
wire n_988;
wire n_1094;
wire n_1097;
wire n_1072;
wire n_1018;
wire n_1078;
wire n_1007;
wire n_1218;
wire n_1003;
wire n_1002;
wire n_1184;
wire n_1208;
wire n_1219;
wire n_1216;
wire n_1221;
wire n_1217;
wire n_1047;
wire n_1030;
wire n_1029;
wire n_1026;
wire n_1393;
wire n_1394;
wire n_1250;
wire n_1293;
wire n_1384;
wire n_1039;
wire n_1369;
wire n_1040;
wire n_1370;
wire n_651;
wire n_1267;
wire n_1207;
wire n_1237;
wire n_1235;
wire n_1309;
wire n_1241;
wire n_1281;
wire n_1292;
wire n_1238;
wire n_1283;
wire n_451;
wire n_519;
wire n_927;
wire n_1400;
wire n_537;
wire n_931;
wire n_930;
wire n_533;
wire n_539;
wire n_449;
wire n_535;
wire n_517;
wire n_407;
wire n_459;
wire n_267;
wire n_994;
wire n_275;
wire n_263;
wire n_387;
wire n_363;
wire n_1117;
wire n_1347;
wire n_1090;
wire n_1365;
wire n_1044;
wire n_17;
wire n_19;
wire n_21;
wire n_1059;
wire n_1362;
wire n_1075;
wire n_1367;
wire n_1169;
wire n_1173;
wire n_1067;
wire n_1073;
wire n_1071;
wire n_1391;
wire n_1091;
wire sgo__n166;
wire n_1392;
wire n_1076;
wire n_1074;
wire n_1328;
wire n_1081;
wire n_1080;
wire n_1327;
wire n_1395;
wire n_1396;
wire n_1098;
wire n_1100;
wire n_1099;
wire n_1353;
wire n_1107;
wire n_1101;
wire n_1352;
wire n_1344;
wire n_1350;
wire n_1371;
wire n_1111;
wire n_1110;
wire n_1114;
wire n_1124;
wire n_1118;
wire n_1113;
wire n_1120;
wire n_1368;
wire n_0;
wire n_1348;
wire n_1377;
wire n_1355;
wire n_1378;
wire n_1379;
wire slo__n638;
wire n_1127;
wire n_1126;
wire n_1331;
wire n_1374;
wire n_1130;
wire n_1145;
wire n_1269;
wire n_1;
wire n_7;
wire n_6;
wire n_1342;
wire CLOCK_slo__xsl_n2867;
wire n_739;
wire n_1340;
wire n_733;
wire n_1341;
wire n_614;
wire n_616;
wire n_553;
wire n_590;
wire n_665;
wire n_592;
wire n_727;
wire slo__sro_n902;
wire n_729;
wire n_1361;
wire n_1056;
wire n_1077;
wire slo__sro_n366;
wire n_1095;
wire n_1096;
wire sgo__sro_n17;
wire n_1033;
wire n_1070;
wire n_1174;
wire n_1398;
wire n_1346;
wire sgo__sro_n101;
wire n_1386;
wire n_9;
wire n_1373;
wire n_2;
wire n_3;
wire n_1376;
wire n_1389;
wire n_5;
wire n_1287;
wire n_1306;
wire n_1245;
wire n_8;
wire n_1274;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_51;
wire slo__sro_n1193;
wire n_55;
wire n_53;
wire n_58;
wire n_57;
wire n_65;
wire n_59;
wire n_63;
wire n_61;
wire n_103;
wire n_67;
wire n_101;
wire n_75;
wire n_79;
wire n_83;
wire n_107;
wire n_20;
wire n_109;
wire n_18;
wire n_22;
wire n_122;
wire n_111;
wire n_126;
wire n_124;
wire n_142;
wire n_24;
wire n_30;
wire n_147;
wire n_26;
wire n_149;
wire n_28;
wire n_157;
wire n_151;
wire n_153;
wire n_155;
wire n_181;
wire n_159;
wire n_178;
wire n_161;
wire n_183;
wire n_179;
wire n_35;
wire n_34;
wire n_37;
wire n_36;
wire n_33;
wire n_32;
wire n_39;
wire n_187;
wire n_48;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_45;
wire n_44;
wire n_47;
wire n_46;
wire n_189;
wire n_54;
wire n_191;
wire n_52;
wire n_193;
wire n_50;
wire n_195;
wire n_56;
wire n_198;
wire n_197;
wire n_262;
wire n_199;
wire n_241;
wire n_265;
wire n_279;
wire n_277;
wire n_269;
wire n_281;
wire n_64;
wire n_283;
wire n_66;
wire n_285;
wire n_62;
wire n_286;
wire n_60;
wire n_287;
wire n_68;
wire n_310;
wire n_70;
wire n_367;
wire n_365;
wire n_369;
wire n_76;
wire n_371;
wire n_78;
wire n_373;
wire n_74;
wire n_375;
wire n_72;
wire n_377;
wire n_80;
wire n_379;
wire n_82;
wire n_381;
wire n_391;
wire n_385;
wire n_389;
wire n_390;
wire n_393;
wire n_102;
wire n_395;
wire n_100;
wire n_397;
wire n_98;
wire n_399;
wire n_106;
wire n_91;
wire n_90;
wire n_95;
wire n_94;
wire n_89;
wire n_88;
wire n_87;
wire n_86;
wire n_85;
wire n_84;
wire n_401;
wire n_104;
wire n_93;
wire n_92;
wire n_403;
wire n_108;
wire n_405;
wire n_411;
wire n_409;
wire n_415;
wire n_413;
wire n_421;
wire sgo__sro_n75;
wire n_419;
wire n_131;
wire n_130;
wire n_129;
wire n_128;
wire n_117;
wire n_116;
wire n_115;
wire n_114;
wire n_135;
wire n_134;
wire n_139;
wire n_138;
wire n_121;
wire n_120;
wire n_125;
wire n_425;
wire n_113;
wire n_112;
wire n_119;
wire n_118;
wire n_133;
wire n_132;
wire n_137;
wire n_136;
wire n_123;
wire n_427;
wire n_141;
wire n_140;
wire n_143;
wire n_429;
wire n_431;
wire n_144;
wire n_433;
wire n_152;
wire n_435;
wire n_156;
wire n_437;
wire n_150;
wire n_439;
wire n_148;
wire n_441;
wire n_146;
wire n_443;
wire n_154;
wire n_445;
wire slo__sro_n1778;
wire n_160;
wire n_163;
wire n_162;
wire n_171;
wire n_170;
wire slo__sro_n802;
wire n_174;
wire n_169;
wire n_168;
wire n_167;
wire n_166;
wire n_165;
wire n_164;
wire n_173;
wire n_172;
wire n_177;
wire n_176;
wire n_457;
wire n_127;
wire n_461;
wire n_182;
wire n_463;
wire n_180;
wire n_465;
wire n_192;
wire n_467;
wire n_186;
wire n_469;
wire n_184;
wire n_471;
wire n_190;
wire n_472;
wire n_188;
wire n_473;
wire slo__sro_n742;
wire n_498;
wire n_196;
wire n_503;
wire n_501;
wire n_509;
wire n_505;
wire n_513;
wire n_531;
wire n_515;
wire sgo__sro_n9;
wire n_541;
wire n_549;
wire n_547;
wire n_521;
wire n_529;
wire n_227;
wire n_225;
wire n_251;
wire n_250;
wire n_226;
wire n_224;
wire n_222;
wire n_233;
wire n_232;
wire n_220;
wire slo__sro_n1830;
wire n_228;
wire n_235;
wire n_234;
wire slo__sro_n1816;
wire n_213;
wire n_211;
wire n_215;
wire n_237;
wire n_236;
wire n_239;
wire n_248;
wire n_246;
wire n_244;
wire n_255;
wire n_254;
wire n_242;
wire slo__sro_n764;
wire n_257;
wire n_256;
wire n_261;
wire n_260;
wire n_206;
wire n_210;
wire n_204;
wire n_202;
wire n_200;
wire n_212;
wire n_217;
wire n_216;
wire n_240;
wire n_209;
wire n_208;
wire n_214;
wire n_219;
wire slo__sro_n726;
wire n_243;
wire n_203;
wire n_201;
wire n_223;
wire n_221;
wire n_207;
wire n_205;
wire slo__sro_n790;
wire n_557;
wire n_268;
wire n_559;
wire n_266;
wire n_561;
wire n_264;
wire n_563;
wire n_278;
wire n_249;
wire n_565;
wire n_272;
wire n_567;
wire n_270;
wire n_569;
wire n_276;
wire n_571;
wire n_282;
wire n_247;
wire n_245;
wire n_572;
wire n_274;
wire n_573;
wire n_280;
wire n_588;
wire n_284;
wire n_594;
wire n_641;
wire n_647;
wire n_643;
wire n_314;
wire n_312;
wire n_322;
wire n_329;
wire n_328;
wire n_340;
wire n_338;
wire n_325;
wire n_355;
wire n_354;
wire n_346;
wire n_344;
wire n_342;
wire n_353;
wire n_352;
wire n_359;
wire n_358;
wire n_300;
wire n_307;
wire n_306;
wire n_303;
wire n_301;
wire n_324;
wire n_331;
wire n_330;
wire n_302;
wire n_304;
wire n_309;
wire n_308;
wire n_335;
wire n_334;
wire n_350;
wire n_348;
wire n_327;
wire n_357;
wire n_356;
wire n_305;
wire n_326;
wire n_333;
wire n_361;
wire n_663;
wire slo__sro_n716;
wire n_288;
wire n_298;
wire n_320;
wire n_318;
wire n_316;
wire n_337;
wire n_336;
wire n_296;
wire n_294;
wire n_292;
wire n_290;
wire n_667;
wire n_368;
wire n_669;
wire n_366;
wire n_671;
wire n_364;
wire n_673;
wire n_380;
wire n_321;
wire n_319;
wire n_317;
wire n_349;
wire n_675;
wire n_372;
wire n_677;
wire n_370;
wire n_679;
wire n_378;
wire n_315;
wire n_313;
wire n_295;
wire n_293;
wire n_291;
wire n_323;
wire n_351;
wire n_343;
wire n_341;
wire n_339;
wire n_681;
wire n_376;
wire n_347;
wire n_345;
wire n_683;
wire n_374;
wire n_685;
wire n_382;
wire n_687;
wire n_386;
wire n_289;
wire n_299;
wire n_297;
wire n_689;
wire n_384;
wire slo__sro_n927;
wire n_711;
wire n_693;
wire n_717;
wire n_712;
wire n_715;
wire n_721;
wire n_738;
wire n_719;
wire n_735;
wire n_723;
wire n_725;
wire n_767;
wire slo__n419;
wire n_771;
wire n_398;
wire n_773;
wire n_396;
wire n_775;
wire n_394;
wire n_776;
wire n_408;
wire n_777;
wire n_414;
wire n_779;
wire n_781;
wire n_406;
wire n_783;
wire n_412;
wire n_785;
wire n_392;
wire n_786;
wire n_404;
wire n_787;
wire n_402;
wire n_789;
wire n_410;
wire n_791;
wire n_416;
wire n_795;
wire n_793;
wire n_797;
wire n_799;
wire n_801;
wire slo__sro_n1021;
wire n_805;
wire n_807;
wire n_430;
wire n_809;
wire n_422;
wire n_811;
wire n_420;
wire n_910;
wire n_812;
wire n_434;
wire n_813;
wire n_438;
wire n_814;
wire n_426;
wire n_818;
wire n_424;
wire n_907;
wire n_822;
wire n_432;
wire n_828;
wire n_428;
wire n_829;
wire n_436;
wire n_831;
wire n_440;
wire n_832;
wire slo__sro_n1207;
wire n_833;
wire n_444;
wire n_835;
wire n_846;
wire n_856;
wire n_854;
wire n_839;
wire n_836;
wire n_844;
wire n_841;
wire n_851;
wire n_859;
wire n_452;
wire n_905;
wire n_861;
wire n_458;
wire n_864;
wire n_450;
wire n_866;
wire n_448;
wire n_871;
wire n_446;
wire n_874;
wire n_460;
wire n_876;
wire n_466;
wire n_877;
wire n_456;
wire n_903;
wire n_879;
wire n_462;
wire n_881;
wire n_454;
wire n_884;
wire n_464;
wire n_886;
wire n_468;
wire n_891;
wire n_470;
wire n_909;
wire n_917;
wire n_916;
wire n_901;
wire n_899;
wire n_906;
wire n_904;
wire n_911;
wire n_908;
wire n_493;
wire n_492;
wire n_496;
wire n_481;
wire n_480;
wire n_479;
wire n_478;
wire n_487;
wire n_486;
wire n_485;
wire n_484;
wire n_483;
wire n_482;
wire n_491;
wire n_490;
wire n_919;
wire n_500;
wire n_898;
wire n_920;
wire n_514;
wire n_921;
wire n_518;
wire n_477;
wire n_476;
wire n_475;
wire n_474;
wire n_900;
wire n_489;
wire n_488;
wire n_495;
wire n_494;
wire n_923;
wire n_506;
wire n_924;
wire n_504;
wire n_925;
wire n_502;
wire n_928;
wire n_512;
wire n_902;
wire n_929;
wire n_510;
wire n_933;
wire n_508;
wire n_934;
wire n_516;
wire slo__sro_n1267;
wire n_936;
wire slo__sro_n1277;
wire n_937;
wire n_524;
wire n_939;
wire n_962;
wire n_942;
wire n_940;
wire n_957;
wire n_963;
wire n_960;
wire n_954;
wire n_945;
wire n_946;
wire n_964;
wire n_530;
wire n_965;
wire n_528;
wire n_966;
wire n_526;
wire n_967;
wire n_538;
wire n_968;
wire n_534;
wire n_895;
wire n_969;
wire n_540;
wire n_970;
wire n_544;
wire n_971;
wire n_532;
wire n_972;
wire n_536;
wire n_973;
wire n_542;
wire n_974;
wire n_546;
wire n_976;
wire n_980;
wire n_977;
wire n_978;
wire n_979;
wire n_1001;
wire n_982;
wire n_985;
wire n_986;
wire n_997;
wire n_990;
wire n_987;
wire n_999;
wire n_989;
wire CLOCK_sgo__sro_n2704;
wire n_995;
wire n_996;
wire n_1397;
wire n_998;
wire n_1004;
wire n_556;
wire n_1005;
wire n_560;
wire n_1006;
wire n_566;
wire n_1008;
wire n_554;
wire n_1009;
wire n_552;
wire n_1010;
wire n_550;
wire n_1011;
wire n_562;
wire n_897;
wire n_1012;
wire n_893;
wire n_1014;
wire n_564;
wire n_1015;
wire n_568;
wire slo__sro_n1494;
wire n_1017;
wire n_1019;
wire n_1025;
wire n_1023;
wire n_1027;
wire n_1024;
wire n_1021;
wire n_1020;
wire n_1022;
wire n_579;
wire n_578;
wire n_577;
wire n_576;
wire n_603;
wire n_602;
wire n_623;
wire n_622;
wire n_889;
wire n_627;
wire n_626;
wire slo__sro_n1367;
wire n_575;
wire n_574;
wire n_581;
wire n_580;
wire n_892;
wire n_605;
wire slo__sro_n1130;
wire n_888;
wire n_621;
wire n_620;
wire n_619;
wire n_618;
wire n_885;
wire n_629;
wire n_628;
wire n_633;
wire n_632;
wire n_585;
wire n_584;
wire n_589;
wire n_1028;
wire n_611;
wire n_610;
wire n_601;
wire n_600;
wire n_599;
wire n_598;
wire n_597;
wire n_596;
wire n_624;
wire n_607;
wire n_606;
wire n_631;
wire n_630;
wire n_890;
wire n_587;
wire slo__sro_n1393;
wire n_613;
wire n_612;
wire slo__sro_n1150;
wire n_591;
wire n_1031;
wire slo__sro_n1355;
wire n_637;
wire n_1034;
wire n_644;
wire n_1035;
wire n_650;
wire n_1036;
wire n_642;
wire n_887;
wire n_1037;
wire n_646;
wire n_1038;
wire n_640;
wire n_1041;
wire n_638;
wire n_883;
wire n_1042;
wire n_648;
wire n_1043;
wire n_652;
wire n_654;
wire n_1046;
wire n_656;
wire n_1060;
wire n_1064;
wire n_1062;
wire n_1052;
wire n_1048;
wire n_1051;
wire n_1049;
wire n_1055;
wire n_1061;
wire n_1050;
wire n_1066;
wire n_1053;
wire n_1054;
wire n_1065;
wire n_1063;
wire n_1058;
wire n_1057;
wire n_593;
wire n_1068;
wire n_1069;
wire n_595;
wire n_1079;
wire n_658;
wire n_1082;
wire n_664;
wire n_880;
wire n_1084;
wire n_668;
wire n_1085;
wire n_662;
wire n_1086;
wire n_660;
wire n_1087;
wire n_666;
wire n_1088;
wire n_670;
wire n_1089;
wire slo__sro_n1106;
wire n_1092;
wire n_674;
wire n_1093;
wire n_1102;
wire n_1103;
wire n_1104;
wire n_1106;
wire n_1108;
wire n_1109;
wire sgo__sro_n14;
wire n_1116;
wire n_1119;
wire n_1122;
wire n_1123;
wire n_1128;
wire n_1129;
wire n_1132;
wire n_1133;
wire n_1134;
wire n_1135;
wire n_1138;
wire n_680;
wire n_1139;
wire n_678;
wire n_1140;
wire n_684;
wire n_1141;
wire n_676;
wire n_882;
wire n_1142;
wire n_682;
wire n_878;
wire slo__sro_n832;
wire n_1144;
wire n_688;
wire n_1146;
wire n_690;
wire n_1147;
wire sgo__sro_n54;
wire n_1152;
wire n_1155;
wire n_1154;
wire n_1153;
wire n_1148;
wire n_1150;
wire n_1149;
wire n_1151;
wire n_1156;
wire n_695;
wire n_694;
wire n_875;
wire n_703;
wire n_702;
wire n_699;
wire n_698;
wire n_697;
wire n_696;
wire n_701;
wire n_700;
wire n_705;
wire n_704;
wire n_707;
wire slo__sro_n1700;
wire n_709;
wire n_708;
wire n_1157;
wire n_710;
wire n_1158;
wire n_714;
wire n_873;
wire n_1159;
wire n_718;
wire n_1176;
wire n_1161;
wire n_716;
wire n_720;
wire n_1163;
wire n_722;
wire n_1164;
wire n_724;
wire n_1188;
wire n_1197;
wire n_1196;
wire n_1165;
wire n_1168;
wire n_1166;
wire n_1167;
wire n_1171;
wire n_1170;
wire n_1172;
wire n_713;
wire n_1177;
wire n_730;
wire n_870;
wire n_1178;
wire n_734;
wire n_1179;
wire n_728;
wire n_1180;
wire n_726;
wire n_1181;
wire n_732;
wire n_1182;
wire n_736;
wire n_1183;
wire n_1185;
wire n_1189;
wire n_1186;
wire n_1187;
wire n_1192;
wire n_1199;
wire n_1195;
wire n_1191;
wire slo__sro_n587;
wire n_1193;
wire n_1198;
wire n_743;
wire n_742;
wire n_757;
wire n_756;
wire n_755;
wire n_754;
wire n_865;
wire n_761;
wire n_760;
wire n_741;
wire n_740;
wire n_872;
wire n_745;
wire n_744;
wire n_869;
wire n_759;
wire n_758;
wire n_747;
wire n_746;
wire n_868;
wire n_749;
wire slo__sro_n1732;
wire n_763;
wire n_762;
wire n_751;
wire n_750;
wire n_1200;
wire n_764;
wire n_1201;
wire n_768;
wire n_867;
wire n_1202;
wire n_770;
wire n_1203;
wire n_766;
wire n_863;
wire CLOCK_sgo__sro_n2645;
wire n_1205;
wire n_774;
wire slo__sro_n1854;
wire n_753;
wire n_1224;
wire n_1231;
wire n_1227;
wire n_1212;
wire n_1209;
wire n_1211;
wire n_1229;
wire n_1226;
wire n_1228;
wire n_1210;
wire n_1230;
wire n_1215;
wire n_1213;
wire n_1214;
wire n_1220;
wire n_1223;
wire n_1225;
wire n_1222;
wire n_1232;
wire n_778;
wire n_860;
wire n_1233;
wire n_782;
wire n_1234;
wire n_780;
wire n_1236;
wire n_784;
wire n_1239;
wire n_1240;
wire n_1242;
wire n_1243;
wire n_1244;
wire n_1248;
wire n_1246;
wire n_1252;
wire n_1253;
wire n_1256;
wire n_1247;
wire n_1249;
wire n_1251;
wire n_1258;
wire n_1254;
wire n_1257;
wire n_1255;
wire sgo__sro_n16;
wire n_1259;
wire n_1261;
wire n_788;
wire n_858;
wire n_1262;
wire n_792;
wire n_862;
wire n_1263;
wire n_790;
wire n_1264;
wire n_794;
wire n_1265;
wire n_796;
wire n_1276;
wire n_1270;
wire n_1277;
wire n_1275;
wire n_1271;
wire n_1266;
wire n_1268;
wire n_1272;
wire n_1273;
wire n_1278;
wire n_798;
wire n_1279;
wire n_800;
wire n_855;
wire n_1280;
wire n_802;
wire n_804;
wire n_1282;
wire n_1285;
wire n_1284;
wire n_1286;
wire n_1288;
wire n_1289;
wire n_806;
wire n_857;
wire n_1290;
wire n_808;
wire n_853;
wire n_1291;
wire n_810;
wire n_1311;
wire n_1307;
wire n_1312;
wire n_1310;
wire n_1294;
wire n_1299;
wire n_1304;
wire n_1302;
wire n_1301;
wire n_1297;
wire n_1305;
wire n_1295;
wire n_1296;
wire n_1298;
wire n_1300;
wire n_1313;
wire n_1308;
wire n_1303;
wire n_852;
wire n_821;
wire n_820;
wire n_849;
wire n_827;
wire n_826;
wire n_815;
wire n_1314;
wire n_848;
wire n_823;
wire n_1316;
wire n_845;
wire n_1318;
wire n_1317;
wire n_847;
wire n_843;
wire n_1319;
wire n_830;
wire n_1321;
wire n_1320;
wire n_1332;
wire n_1343;
wire n_1336;
wire n_1326;
wire n_1322;
wire n_1325;
wire n_1337;
wire n_1335;
wire n_1323;
wire n_1334;
wire n_1333;
wire n_1324;
wire n_1338;
wire n_1330;
wire n_1329;
wire n_840;
wire n_834;
wire n_1345;
wire n_1349;
wire n_842;
wire n_838;
wire n_837;
wire n_1351;
wire n_1360;
wire n_1364;
wire n_1354;
wire n_1356;
wire n_1357;
wire n_1358;
wire n_1366;
wire n_1359;
wire n_1372;
wire sgo__sro_n8;
wire n_1375;
wire n_1380;
wire n_1381;
wire n_1383;
wire n_850;
wire n_817;
wire n_816;
wire n_825;
wire n_824;
wire n_819;
wire n_1385;
wire n_1387;
wire n_1390;
wire n_1388;
wire n_1399;
wire sgo__sro_n55;
wire sgo__sro_n84;
wire sgo__sro_n87;
wire sgo__sro_n32;
wire sgo__sro_n33;
wire sgo__sro_n34;
wire sgo__n97;
wire sgo__sro_n102;
wire sgo__sro_n105;
wire sgo__n107;
wire sgo__sro_n137;
wire sgo__sro_n138;
wire sgo__n115;
wire sgo__sro_n187;
wire sgo__n199;
wire sgo__sro_n149;
wire sgo__sro_n150;
wire sgo__sro_n151;
wire sgo__n168;
wire sgo__n185;
wire sgo__sro_n191;
wire sgo__n228;
wire sgo__sro_n255;
wire sgo__sro_n293;
wire sgo__n265;
wire sgo__sro_n309;
wire sgo__sro_n310;
wire sgo__sro_n311;
wire slo__sro_n332;
wire slo__sro_n333;
wire slo__n416;
wire slo__n432;
wire slo__sro_n442;
wire slo__sro_n464;
wire slo__sro_n465;
wire slo__sro_n466;
wire slo__sro_n467;
wire slo__sro_n468;
wire slo__sro_n499;
wire slo__n521;
wire slo__sro_n535;
wire slo__sro_n544;
wire slo__sro_n545;
wire slo__sro_n546;
wire slo__n557;
wire slo__sro_n567;
wire slo__sro_n568;
wire slo__sro_n588;
wire slo__sro_n589;
wire CLOCK_slo__n2890;
wire slo__sro_n604;
wire slo__sro_n692;
wire slo__sro_n693;
wire slo__sro_n694;
wire slo__sro_n695;
wire slo__sro_n705;
wire slo__sro_n706;
wire slo__sro_n707;
wire slo__sro_n708;
wire slo__sro_n717;
wire slo__sro_n718;
wire slo__sro_n719;
wire slo__sro_n727;
wire slo__sro_n728;
wire slo__sro_n729;
wire slo__sro_n730;
wire slo__sro_n743;
wire slo__sro_n744;
wire slo__sro_n745;
wire slo__sro_n750;
wire slo__sro_n751;
wire slo__sro_n752;
wire slo__sro_n753;
wire slo__sro_n754;
wire slo__sro_n755;
wire slo__sro_n765;
wire slo__sro_n766;
wire slo__sro_n767;
wire CLOCK_sgo__sro_n2584;
wire slo__sro_n776;
wire slo__sro_n777;
wire slo__sro_n778;
wire slo__sro_n779;
wire slo__sro_n780;
wire slo__sro_n791;
wire slo__sro_n792;
wire slo__sro_n793;
wire slo__sro_n803;
wire slo__sro_n804;
wire slo__sro_n814;
wire slo__sro_n815;
wire slo__sro_n816;
wire slo__sro_n817;
wire slo__sro_n818;
wire slo__sro_n819;
wire slo__sro_n820;
wire slo__sro_n833;
wire slo__sro_n834;
wire slo__sro_n835;
wire slo__sro_n840;
wire slo__sro_n841;
wire slo__sro_n842;
wire slo__sro_n846;
wire slo__sro_n847;
wire slo__sro_n848;
wire slo__sro_n849;
wire slo__sro_n854;
wire slo__sro_n855;
wire slo__sro_n856;
wire slo__sro_n901;
wire slo__xsl_n869;
wire slo__sro_n903;
wire slo__sro_n907;
wire slo__sro_n908;
wire slo__sro_n909;
wire slo__sro_n910;
wire slo__sro_n915;
wire slo__sro_n916;
wire slo__sro_n917;
wire slo__sro_n918;
wire slo__sro_n919;
wire slo__sro_n928;
wire slo__sro_n929;
wire slo__sro_n930;
wire slo__sro_n931;
wire slo__sro_n939;
wire slo__sro_n940;
wire slo__sro_n941;
wire slo__sro_n942;
wire slo__sro_n943;
wire slo__sro_n944;
wire slo__sro_n951;
wire slo__sro_n952;
wire slo__sro_n953;
wire slo__sro_n954;
wire slo__sro_n959;
wire slo__sro_n960;
wire slo__sro_n961;
wire slo__sro_n965;
wire slo__sro_n966;
wire slo__sro_n967;
wire slo__sro_n968;
wire slo__sro_n1020;
wire slo__xsl_n988;
wire slo__sro_n1022;
wire slo__sro_n1023;
wire slo__sro_n1024;
wire slo__sro_n1025;
wire slo__sro_n1032;
wire slo__sro_n1033;
wire slo__sro_n1034;
wire slo__sro_n1040;
wire slo__sro_n1041;
wire slo__sro_n1042;
wire slo__sro_n1043;
wire slo__sro_n1044;
wire slo__sro_n1045;
wire slo__sro_n1046;
wire slo__xsl_n1063;
wire slo__xsl_n1064;
wire slo__sro_n1091;
wire slo__sro_n1108;
wire slo__sro_n1118;
wire slo__sro_n1119;
wire slo__sro_n1120;
wire slo__sro_n1121;
wire slo__sro_n1122;
wire slo__sro_n1131;
wire slo__sro_n1132;
wire slo__sro_n1133;
wire slo__sro_n1134;
wire slo__sro_n1135;
wire slo__sro_n1151;
wire slo__sro_n1152;
wire slo__sro_n1153;
wire slo__sro_n1154;
wire slo__sro_n1155;
wire slo__sro_n1166;
wire slo__sro_n1182;
wire slo__sro_n1183;
wire slo__sro_n1184;
wire slo__sro_n1185;
wire slo__sro_n1194;
wire slo__sro_n1195;
wire slo__sro_n1196;
wire slo__sro_n1208;
wire slo__sro_n1209;
wire slo__sro_n1210;
wire slo__sro_n1211;
wire slo__sro_n1212;
wire slo__sro_n1241;
wire slo__sro_n1242;
wire slo__sro_n1243;
wire slo__sro_n1244;
wire slo__sro_n1253;
wire slo__sro_n1254;
wire slo__sro_n1255;
wire slo__sro_n1256;
wire slo__sro_n1257;
wire slo__sro_n1258;
wire slo__sro_n1268;
wire slo__sro_n1270;
wire slo__sro_n1278;
wire slo__sro_n1279;
wire slo__sro_n1280;
wire slo__sro_n1281;
wire slo__sro_n1282;
wire slo__sro_n1289;
wire slo__sro_n1290;
wire slo__sro_n1291;
wire slo__sro_n1292;
wire slo__sro_n1297;
wire slo__sro_n1298;
wire slo__sro_n1299;
wire slo__sro_n1300;
wire slo__sro_n1331;
wire slo__sro_n1332;
wire slo__sro_n1333;
wire slo__sro_n1334;
wire slo__sro_n1339;
wire slo__sro_n1340;
wire slo__sro_n1341;
wire slo__sro_n1342;
wire slo__sro_n1343;
wire slo__sro_n1356;
wire slo__sro_n1357;
wire slo__sro_n1358;
wire slo__sro_n1359;
wire slo__sro_n1368;
wire slo__sro_n1369;
wire slo__sro_n1370;
wire slo__sro_n1371;
wire slo__sro_n1372;
wire slo__sro_n1379;
wire slo__sro_n1380;
wire slo__sro_n1381;
wire slo__sro_n1382;
wire slo__sro_n1383;
wire CLOCK_sgo__sro_n2583;
wire slo__sro_n1394;
wire slo__sro_n1395;
wire slo__sro_n1396;
wire slo__sro_n1401;
wire slo__sro_n1402;
wire slo__sro_n1403;
wire slo__sro_n1404;
wire slo__sro_n1405;
wire slo__sro_n1439;
wire slo__sro_n1440;
wire slo__sro_n1441;
wire slo__sro_n1442;
wire slo__sro_n1474;
wire slo__sro_n1475;
wire slo__sro_n1476;
wire slo__sro_n1477;
wire slo__sro_n1478;
wire slo__sro_n1479;
wire slo__sro_n1480;
wire slo__sro_n1481;
wire slo__sro_n1495;
wire slo__sro_n1496;
wire slo__sro_n1497;
wire CLOCK_sgo__sro_n2608;
wire slo__sro_n1519;
wire slo__sro_n1520;
wire slo__sro_n1521;
wire slo__sro_n1522;
wire slo__sro_n1537;
wire slo__sro_n1538;
wire slo__sro_n1539;
wire slo__sro_n1540;
wire slo__sro_n1547;
wire slo__sro_n1548;
wire slo__sro_n1549;
wire slo__sro_n1550;
wire slo__sro_n1569;
wire slo__sro_n1570;
wire slo__sro_n1571;
wire slo__sro_n1572;
wire slo__n1579;
wire slo__sro_n1587;
wire slo__sro_n1588;
wire slo__sro_n1589;
wire slo__sro_n1593;
wire slo__sro_n1594;
wire slo__sro_n1595;
wire slo__sro_n1599;
wire slo__sro_n1600;
wire slo__sro_n1601;
wire slo__sro_n1605;
wire slo__sro_n1606;
wire slo__sro_n1607;
wire slo__sro_n1611;
wire slo__sro_n1612;
wire slo__sro_n1613;
wire slo__sro_n1614;
wire slo__sro_n1615;
wire slo__sro_n1621;
wire slo__sro_n1622;
wire slo__sro_n1623;
wire slo__sro_n1624;
wire slo__n1633;
wire slo__sro_n1644;
wire slo__sro_n1645;
wire slo__sro_n1646;
wire slo__sro_n1650;
wire slo__sro_n1651;
wire slo__sro_n1652;
wire slo__sro_n1653;
wire slo__sro_n1654;
wire slo__sro_n1655;
wire slo__sro_n1662;
wire slo__sro_n1663;
wire slo__sro_n1664;
wire slo__sro_n1665;
wire slo__n1685;
wire slo__sro_n1688;
wire slo__sro_n1689;
wire slo__sro_n1690;
wire slo__sro_n1691;
wire slo__sro_n1692;
wire slo__sro_n1701;
wire slo__sro_n1702;
wire slo__sro_n1703;
wire slo__sro_n1704;
wire slo__sro_n1705;
wire slo__sro_n1714;
wire slo__sro_n1715;
wire slo__sro_n1716;
wire slo__sro_n1717;
wire slo__sro_n1718;
wire CLOCK_sgo__n2634;
wire slo__sro_n1733;
wire slo__sro_n1734;
wire slo__sro_n1735;
wire slo__sro_n1736;
wire slo__sro_n1737;
wire slo__sro_n1746;
wire slo__sro_n1747;
wire slo__sro_n1748;
wire slo__sro_n1749;
wire slo__sro_n1756;
wire slo__sro_n1757;
wire slo__sro_n1758;
wire slo__sro_n1759;
wire slo__sro_n1760;
wire slo__sro_n1761;
wire slo__sro_n1762;
wire slo__sro_n1779;
wire slo__sro_n1780;
wire slo__sro_n1781;
wire slo__sro_n1798;
wire slo__sro_n1799;
wire slo__sro_n1800;
wire slo__sro_n1801;
wire slo__sro_n1802;
wire slo__sro_n1803;
wire slo__sro_n1804;
wire slo__sro_n1805;
wire slo__sro_n1817;
wire slo__sro_n1818;
wire slo__sro_n1819;
wire slo__sro_n1820;
wire slo__sro_n1821;
wire slo__sro_n1831;
wire slo__sro_n1832;
wire slo__sro_n1833;
wire slo__sro_n1834;
wire slo__sro_n1835;
wire slo__n1848;
wire slo__sro_n1855;
wire slo__sro_n1856;
wire slo__sro_n1857;
wire slo__sro_n1858;
wire slo__sro_n1859;
wire slo__sro_n1868;
wire slo__sro_n1869;
wire slo__sro_n1870;
wire slo__sro_n1871;
wire slo__sro_n1872;
wire slo__sro_n1873;
wire CLOCK_sgo__n2761;
wire CLOCK_sgo__n2632;
wire opt_ipo_n1905;
wire CLOCK_sgo__sro_n2705;
wire CLOCK_sgo__sro_n2706;
wire CLOCK_slo__xsl_n2800;
wire CLOCK_slo__xsl_n2801;
wire CLOCK_slo__mro_n2819;
wire CLOCK_slo__mro_n2828;
wire opt_ipo_n1924;
wire CLOCK_slo__mro_n2829;
wire CLOCK_slo__sro_n2896;
wire CLOCK_slo__sro_n2897;
wire CLOCK_slo__sro_n2898;
wire opt_ipo_n1940;
wire opt_ipo_n2336;
wire opt_ipo_n2338;
wire opt_ipo_n1948;
wire spw__n3514;
wire opt_ipo_n1965;
wire opt_ipo_n1967;
wire opt_ipo_n2021;
wire opt_ipo_n2091;
wire opt_ipo_n2116;
wire opt_ipo_n2117;
wire opt_ipo_n2150;
wire opt_ipo_n2152;
wire opt_ipo_n2153;
wire opt_ipo_n2154;
wire CLOCK_spw__n3015;
wire opt_ipo_n2168;


NAND2_X1 i_1043 (.ZN (n_1400), .A1 (n_549), .A2 (n_547));
AOI21_X4 i_1042 (.ZN (n_1399), .A (n_519), .B1 (n_549), .B2 (n_547));
NAND4_X2 i_1041 (.ZN (n_1397), .A1 (n_1399), .A2 (n_453), .A3 (n_541), .A4 (n_533));
NAND2_X1 i_1040 (.ZN (n_1396), .A1 (n_1317), .A2 (n_825));
NAND2_X1 i_1039 (.ZN (n_1395), .A1 (n_824), .A2 (n_819));
INV_X1 i_1038 (.ZN (n_1394), .A (n_1395));
NOR2_X1 i_1037 (.ZN (n_1393), .A1 (n_824), .A2 (n_819));
INV_X1 i_1036 (.ZN (n_1392), .A (n_1393));
NOR2_X1 i_1035 (.ZN (n_1391), .A1 (n_1317), .A2 (n_825));
OAI221_X1 i_1034 (.ZN (n_1390), .A (n_1392), .B1 (n_1317), .B2 (n_825), .C1 (n_1318), .C2 (n_1320));
INV_X1 i_1033 (.ZN (n_1389), .A (n_1390));
AOI21_X1 i_1032 (.ZN (n_1388), .A (n_1394), .B1 (n_1384), .B2 (n_1293));
OAI221_X1 i_1031 (.ZN (n_1387), .A (n_1329), .B1 (n_1330), .B2 (n_1396), .C1 (n_1390), .C2 (n_1388));
INV_X1 i_1030 (.ZN (n_1386), .A (n_1387));
XOR2_X1 i_1029 (.Z (n_1385), .A (p_10[54]), .B (p_11[54]));
XOR2_X1 i_1028 (.Z (n_850), .A (n_1334), .B (n_1385));
FA_X1 i_1027 (.CO (n_819), .S (n_1384), .A (n_1290), .B (n_1291), .CI (n_816));
HA_X1 i_1026 (.CO (n_825), .S (n_824), .A (n_817), .B (n_1316));
FA_X1 i_1025 (.CO (n_817), .S (n_816), .A (n_1307), .B (n_1314), .CI (n_850));
INV_X1 i_1024 (.ZN (n_1383), .A (n_1358));
OAI21_X2 sgo__sro_c8 (.ZN (sgo__sro_n9), .A (n_1108), .B1 (n_1022), .B2 (n_978));
OAI22_X1 i_1022 (.ZN (n_1381), .A1 (p_14[60]), .A2 (n_1366), .B1 (n_1383), .B2 (n_1359));
NOR2_X1 i_1021 (.ZN (n_1380), .A1 (p_14[61]), .A2 (n_1381));
INV_X1 i_1020 (.ZN (n_1379), .A (n_1380));
NAND2_X1 i_1019 (.ZN (n_1378), .A1 (p_14[61]), .A2 (n_1381));
NOR2_X1 i_1018 (.ZN (n_1377), .A1 (n_1372), .A2 (n_1354));
NAND2_X1 i_1017 (.ZN (n_1376), .A1 (n_1378), .A2 (n_1377));
AOI21_X1 i_1016 (.ZN (n_1375), .A (n_1376), .B1 (n_1347), .B2 (n_1371));
AOI211_X1 i_1015 (.ZN (n_1374), .A (n_1375), .B (n_1380), .C1 (n_1355), .C2 (n_1378));
OAI21_X1 i_1014 (.ZN (n_1373), .A (n_1374), .B1 (p_14[62]), .B2 (n_1283));
NOR2_X1 i_1013 (.ZN (n_1372), .A1 (n_1344), .A2 (n_1350));
NAND2_X1 i_1012 (.ZN (n_1371), .A1 (n_1344), .A2 (n_1350));
AOI21_X1 i_1011 (.ZN (n_1370), .A (n_1372), .B1 (n_1344), .B2 (n_1350));
INV_X1 i_1010 (.ZN (n_1369), .A (n_1370));
NOR2_X1 i_1009 (.ZN (n_1368), .A1 (n_1355), .A2 (n_1369));
INV_X1 i_1008 (.ZN (n_1366), .A (p_13[60]));
INV_X1 i_1007 (.ZN (n_1364), .A (p_13[58]));
NOR2_X1 i_1006 (.ZN (n_1360), .A1 (p_13[59]), .A2 (p_14[59]));
INV_X1 i_1005 (.ZN (n_1359), .A (n_1360));
NAND2_X1 i_1004 (.ZN (n_1358), .A1 (n_1366), .A2 (p_14[60]));
OAI21_X1 i_1003 (.ZN (n_1357), .A (n_1358), .B1 (n_1366), .B2 (p_14[60]));
XOR2_X1 i_1002 (.Z (n_1356), .A (n_1360), .B (n_1357));
AND2_X1 i_1001 (.ZN (n_1355), .A1 (n_837), .A2 (n_1356));
NOR2_X1 i_1000 (.ZN (n_1354), .A1 (n_837), .A2 (n_1356));
NOR2_X1 i_999 (.ZN (n_1353), .A1 (n_1355), .A2 (n_1354));
INV_X1 i_998 (.ZN (n_1352), .A (n_1353));
OAI222_X1 i_997 (.ZN (n_842), .A1 (p_12[58]), .A2 (n_1349), .B1 (n_1364), .B2 (p_12[58])
    , .C1 (n_1364), .C2 (n_1349));
AOI21_X1 i_996 (.ZN (n_1351), .A (n_1360), .B1 (p_13[59]), .B2 (p_14[59]));
INV_X1 i_995 (.ZN (n_838), .A (n_1351));
HA_X1 i_994 (.CO (n_837), .S (n_1350), .A (n_842), .B (n_838));
INV_X1 i_993 (.ZN (n_1349), .A (p_14[58]));
OR2_X1 i_992 (.ZN (n_1348), .A1 (n_1321), .A2 (n_834));
NAND2_X2 i_991 (.ZN (n_1347), .A1 (n_1321), .A2 (n_834));
AND2_X1 i_990 (.ZN (n_1346), .A1 (n_1348), .A2 (n_1347));
XOR2_X1 i_989 (.Z (n_1345), .A (p_12[58]), .B (p_13[58]));
XNOR2_X1 i_988 (.ZN (n_840), .A (p_14[58]), .B (n_1345));
FA_X1 i_987 (.CO (n_1344), .S (n_834), .A (n_1332), .B (n_840), .CI (n_1319));
INV_X1 i_986 (.ZN (n_1343), .A (p_13[57]));
INV_X1 i_985 (.ZN (n_1338), .A (p_11[56]));
INV_X1 i_984 (.ZN (n_1337), .A (p_11[55]));
INV_X1 i_983 (.ZN (n_1336), .A (p_12[57]));
INV_X1 i_982 (.ZN (n_1335), .A (p_12[55]));
INV_X1 i_981 (.ZN (n_1334), .A (p_12[54]));
INV_X1 i_980 (.ZN (n_1333), .A (p_10[54]));
NAND2_X1 i_979 (.ZN (n_1332), .A1 (n_1343), .A2 (n_1336));
NOR2_X1 i_978 (.ZN (n_1330), .A1 (n_1318), .A2 (n_1320));
NAND2_X1 i_977 (.ZN (n_1329), .A1 (n_1318), .A2 (n_1320));
AOI21_X1 i_976 (.ZN (n_1328), .A (n_1330), .B1 (n_1318), .B2 (n_1320));
INV_X1 i_975 (.ZN (n_1327), .A (n_1328));
NAND2_X1 i_974 (.ZN (n_1326), .A1 (n_1338), .A2 (p_12[56]));
OR2_X1 i_973 (.ZN (n_1325), .A1 (n_1338), .A2 (p_12[56]));
NAND2_X1 i_972 (.ZN (n_1324), .A1 (n_1326), .A2 (n_1325));
XNOR2_X1 i_971 (.ZN (n_845), .A (p_13[56]), .B (n_1324));
NAND2_X1 i_970 (.ZN (n_849), .A1 (n_1337), .A2 (n_1335));
OAI21_X1 i_969 (.ZN (n_1323), .A (p_11[54]), .B1 (p_12[54]), .B2 (n_1333));
OAI21_X1 i_968 (.ZN (n_852), .A (n_1323), .B1 (n_1334), .B2 (p_10[54]));
OAI21_X1 i_967 (.ZN (n_848), .A (n_849), .B1 (n_1337), .B2 (n_1335));
NAND2_X1 i_966 (.ZN (n_1322), .A1 (p_13[56]), .A2 (n_1325));
NAND2_X1 i_965 (.ZN (n_847), .A1 (n_1326), .A2 (n_1322));
OAI21_X1 i_964 (.ZN (n_843), .A (n_1332), .B1 (n_1343), .B2 (n_1336));
HA_X1 i_963 (.CO (n_1321), .S (n_1320), .A (n_827), .B (n_830));
FA_X1 i_962 (.CO (n_1319), .S (n_830), .A (p_14[57]), .B (n_847), .CI (n_843));
FA_X1 i_961 (.CO (n_1318), .S (n_1317), .A (n_845), .B (n_826), .CI (n_823));
FA_X1 i_960 (.CO (n_823), .S (n_1316), .A (n_815), .B (n_820), .CI (n_848));
FA_X1 i_959 (.CO (n_815), .S (n_1314), .A (p_13[54]), .B (p_14[54]), .CI (n_1289));
FA_X1 i_958 (.CO (n_827), .S (n_826), .A (p_14[56]), .B (n_849), .CI (n_821));
FA_X1 i_957 (.CO (n_821), .S (n_820), .A (p_13[55]), .B (p_14[55]), .CI (n_852));
INV_X1 i_956 (.ZN (n_1313), .A (n_1248));
INV_X1 i_955 (.ZN (n_1312), .A (p_10[53]));
INV_X1 i_954 (.ZN (n_1311), .A (p_10[52]));
INV_X1 i_953 (.ZN (n_1310), .A (p_11[53]));
INV_X1 i_952 (.ZN (n_1309), .A (n_1286));
INV_X1 i_951 (.ZN (n_1308), .A (n_1287));
NAND2_X1 i_950 (.ZN (n_1307), .A1 (n_1312), .A2 (n_1310));
NOR2_X1 i_949 (.ZN (n_1306), .A1 (n_1292), .A2 (n_1281));
AOI21_X1 i_948 (.ZN (n_1305), .A (n_1306), .B1 (n_1292), .B2 (n_1281));
INV_X1 i_947 (.ZN (n_1304), .A (n_1305));
AOI21_X1 i_946 (.ZN (n_1303), .A (n_1269), .B1 (n_1268), .B2 (n_1274));
OAI21_X1 i_945 (.ZN (n_1302), .A (n_1309), .B1 (n_1308), .B2 (n_1303));
NAND3_X1 i_944 (.ZN (n_1301), .A1 (n_1246), .A2 (n_1253), .A3 (n_1252));
OAI211_X1 i_943 (.ZN (n_1300), .A (n_1305), .B (n_1273), .C1 (n_1301), .C2 (n_1313));
NOR3_X1 i_942 (.ZN (n_1299), .A1 (n_1300), .A2 (n_1269), .A3 (n_1286));
AND2_X1 i_941 (.ZN (n_1298), .A1 (n_1268), .A2 (n_1243));
NAND3_X1 i_940 (.ZN (n_1297), .A1 (n_1248), .A2 (n_1287), .A3 (n_1298));
OAI21_X1 i_939 (.ZN (n_1296), .A (n_1287), .B1 (n_1269), .B2 (n_1298));
INV_X1 i_938 (.ZN (n_1295), .A (n_1296));
OAI33_X1 i_937 (.ZN (n_1294), .A1 (n_1301), .A2 (n_1297), .A3 (n_1305), .B1 (n_1286)
    , .B2 (n_1304), .B3 (n_1295));
OAI21_X1 slo__sro_c1634 (.ZN (slo__sro_n1107), .A (slo__sro_n1341), .B1 (slo__sro_n1130), .B2 (n_632));
OAI21_X1 i_935 (.ZN (n_853), .A (n_1307), .B1 (n_1312), .B2 (n_1310));
OAI222_X1 i_934 (.ZN (n_857), .A1 (p_9[52]), .A2 (n_1288), .B1 (n_1311), .B2 (p_9[52])
    , .C1 (n_1311), .C2 (n_1288));
HA_X1 i_933 (.CO (n_1293), .S (n_1292), .A (n_1280), .B (n_810));
FA_X1 i_932 (.CO (n_1291), .S (n_810), .A (n_853), .B (n_1279), .CI (n_808));
FA_X1 i_931 (.CO (n_1290), .S (n_808), .A (n_1278), .B (n_857), .CI (n_806));
FA_X1 i_930 (.CO (n_1289), .S (n_806), .A (p_12[53]), .B (p_13[53]), .CI (p_14[53]));
INV_X1 i_929 (.ZN (n_1288), .A (p_11[52]));
NAND2_X1 i_928 (.ZN (n_1287), .A1 (n_1265), .A2 (n_804));
NOR2_X1 i_927 (.ZN (n_1286), .A1 (n_1265), .A2 (n_804));
OAI21_X1 i_926 (.ZN (n_1285), .A (n_1287), .B1 (n_1265), .B2 (n_804));
AOI21_X2 i_925 (.ZN (n_1284), .A (n_1269), .B1 (n_1271), .B2 (n_1268));
XNOR2_X2 i_924 (.ZN (\aggregated_res[14] [52] ), .A (n_1284), .B (n_1285));
XOR2_X1 i_923 (.Z (n_1282), .A (p_9[52]), .B (p_10[52]));
XNOR2_X1 i_922 (.ZN (n_855), .A (p_11[52]), .B (n_1282));
FA_X1 i_921 (.CO (n_1281), .S (n_804), .A (n_1262), .B (n_802), .CI (n_1264));
FA_X1 i_920 (.CO (n_1280), .S (n_802), .A (n_798), .B (n_855), .CI (n_800));
FA_X1 i_919 (.CO (n_1279), .S (n_800), .A (n_1261), .B (n_1270), .CI (n_1263));
FA_X1 i_918 (.CO (n_1278), .S (n_798), .A (p_12[52]), .B (p_13[52]), .CI (p_14[52]));
INV_X1 i_917 (.ZN (n_1277), .A (p_9[51]));
INV_X1 i_916 (.ZN (n_1276), .A (p_9[50]));
INV_X1 i_915 (.ZN (n_1275), .A (p_10[51]));
NOR2_X1 i_914 (.ZN (n_1274), .A1 (n_1237), .A2 (n_1207));
INV_X1 i_913 (.ZN (n_1273), .A (n_1274));
AOI21_X2 i_912 (.ZN (n_1272), .A (n_1274), .B1 (n_1244), .B2 (n_1243));
INV_X4 i_911 (.ZN (n_1271), .A (n_1272));
NAND2_X1 i_910 (.ZN (n_1270), .A1 (n_1277), .A2 (n_1275));
NOR2_X2 i_909 (.ZN (n_1269), .A1 (n_1239), .A2 (n_796));
NAND2_X1 i_908 (.ZN (n_1268), .A1 (n_1239), .A2 (n_796));
INV_X1 i_907 (.ZN (n_1267), .A (n_1268));
NOR2_X1 i_906 (.ZN (n_1266), .A1 (n_1269), .A2 (n_1267));
XNOR2_X2 i_905 (.ZN (\aggregated_res[14] [51] ), .A (n_1271), .B (n_1266));
OAI21_X1 i_904 (.ZN (n_858), .A (n_1270), .B1 (n_1277), .B2 (n_1275));
OAI222_X1 i_903 (.ZN (n_862), .A1 (p_8[50]), .A2 (n_1259), .B1 (n_1276), .B2 (p_8[50])
    , .C1 (n_1276), .C2 (n_1259));
HA_X1 i_902 (.CO (n_1265), .S (n_796), .A (n_792), .B (n_794));
FA_X1 i_901 (.CO (n_1264), .S (n_794), .A (n_790), .B (n_1233), .CI (n_1236));
FA_X1 i_900 (.CO (n_1263), .S (n_790), .A (p_14[51]), .B (n_1232), .CI (n_862));
FA_X1 i_899 (.CO (n_1262), .S (n_792), .A (n_1234), .B (n_788), .CI (n_858));
FA_X1 i_898 (.CO (n_1261), .S (n_788), .A (p_11[51]), .B (p_12[51]), .CI (p_13[51]));
AND2_X2 sgo__sro_c79 (.ZN (sgo__sro_n55), .A1 (n_1102), .A2 (n_1057));
INV_X1 i_896 (.ZN (n_1259), .A (p_10[50]));
NOR3_X4 i_895 (.ZN (n_1258), .A1 (n_1223), .A2 (n_1220), .A3 (n_1216));
OAI21_X2 i_894 (.ZN (n_1257), .A (n_1258), .B1 (n_1164), .B2 (n_1183));
INV_X1 i_893 (.ZN (n_1256), .A (n_1257));
NOR2_X1 i_892 (.ZN (n_1255), .A1 (n_1078), .A2 (n_1018));
OAI21_X2 sgo__sro_c80 (.ZN (sgo__sro_n54), .A (sgo__sro_n55), .B1 (n_1104), .B2 (n_1103));
NAND3_X2 i_890 (.ZN (n_1253), .A1 (n_985), .A2 (n_1119), .A3 (n_1254));
NAND2_X1 i_889 (.ZN (n_1252), .A1 (n_1116), .A2 (slo__n521));
OAI21_X1 i_888 (.ZN (n_1251), .A (n_1258), .B1 (n_1225), .B2 (n_1219));
OAI21_X2 i_887 (.ZN (n_1249), .A (n_1251), .B1 (n_1223), .B2 (n_1222));
AOI21_X4 i_886 (.ZN (n_1248), .A (n_1249), .B1 (sgo__n228), .B2 (n_1200));
NOR2_X2 i_885 (.ZN (n_1247), .A1 (n_1106), .A2 (opt_ipo_n2168));
OAI21_X2 i_884 (.ZN (n_1246), .A (n_1256), .B1 (n_1191), .B2 (n_1247));
NAND4_X4 i_883 (.ZN (n_1245), .A1 (n_1246), .A2 (n_1248), .A3 (n_1252), .A4 (n_1253));
INV_X1 i_882 (.ZN (n_1244), .A (n_1245));
NAND2_X1 i_881 (.ZN (n_1243), .A1 (n_1237), .A2 (n_1207));
OAI21_X1 i_880 (.ZN (n_1242), .A (n_1243), .B1 (n_1237), .B2 (n_1207));
XNOR2_X2 i_879 (.ZN (\aggregated_res[14] [50] ), .A (slo___n509), .B (n_1242));
XOR2_X1 i_878 (.Z (n_1240), .A (p_8[50]), .B (p_9[50]));
XNOR2_X1 i_877 (.ZN (n_860), .A (p_10[50]), .B (n_1240));
FA_X1 i_876 (.CO (n_1239), .S (n_1237), .A (n_782), .B (n_784), .CI (n_1205));
FA_X1 i_875 (.CO (n_1236), .S (n_784), .A (n_780), .B (n_1202), .CI (slo__sro_n1870));
FA_X1 i_874 (.CO (n_1234), .S (n_780), .A (p_14[50]), .B (n_1203), .CI (n_1224));
FA_X1 i_873 (.CO (n_1233), .S (n_782), .A (n_1201), .B (n_778), .CI (n_860));
FA_X1 i_872 (.CO (n_1232), .S (n_778), .A (p_11[50]), .B (p_12[50]), .CI (p_13[50]));
INV_X1 i_871 (.ZN (n_1231), .A (p_9[49]));
INV_X1 i_870 (.ZN (n_1230), .A (p_7[48]));
INV_X1 i_869 (.ZN (n_1229), .A (p_7[47]));
INV_X1 i_868 (.ZN (n_1228), .A (p_7[46]));
INV_X1 i_867 (.ZN (n_1227), .A (p_8[49]));
INV_X1 i_866 (.ZN (n_1226), .A (p_8[47]));
INV_X1 i_865 (.ZN (n_1225), .A (n_1187));
NAND2_X1 i_864 (.ZN (n_1224), .A1 (n_1231), .A2 (n_1227));
NOR2_X2 i_863 (.ZN (n_1223), .A1 (sgo__n228), .A2 (n_1200));
NAND2_X1 i_862 (.ZN (n_1222), .A1 (n_764), .A2 (n_753));
INV_X1 i_861 (.ZN (n_1221), .A (n_1222));
NOR2_X1 i_860 (.ZN (n_1220), .A1 (n_1184), .A2 (n_1208));
AND2_X1 i_859 (.ZN (n_1219), .A1 (n_1208), .A2 (n_1184));
NOR2_X1 i_858 (.ZN (n_1218), .A1 (n_1220), .A2 (n_1219));
OAI21_X1 sgo__sro_c253 (.ZN (sgo__sro_n138), .A (n_729), .B1 (n_727), .B2 (slo__xsl_n869));
NOR2_X2 i_856 (.ZN (n_1216), .A1 (n_764), .A2 (n_753));
AOI21_X1 i_855 (.ZN (n_1215), .A (n_1223), .B1 (n_1200), .B2 (sgo__n228));
INV_X1 sgo__sro_c553 (.ZN (sgo__sro_n293), .A (n_217));
NAND2_X2 sgo__sro_c584 (.ZN (sgo__sro_n309), .A1 (sgo__sro_n311), .A2 (sgo__sro_n310));
NAND2_X2 slo__sro_c769 (.ZN (slo__sro_n460), .A1 (n_1245), .A2 (n_8));
NAND2_X1 i_851 (.ZN (n_1212), .A1 (n_1230), .A2 (p_8[48]));
OR2_X1 i_850 (.ZN (n_1211), .A1 (n_1230), .A2 (p_8[48]));
NAND2_X1 i_849 (.ZN (n_1210), .A1 (n_1212), .A2 (n_1211));
XNOR2_X1 i_848 (.ZN (n_865), .A (p_9[48]), .B (n_1210));
NAND2_X1 i_847 (.ZN (n_869), .A1 (n_1229), .A2 (n_1226));
OAI222_X1 i_846 (.ZN (n_872), .A1 (p_6[46]), .A2 (n_1198), .B1 (n_1228), .B2 (p_6[46])
    , .C1 (n_1228), .C2 (n_1198));
OAI21_X1 i_845 (.ZN (n_868), .A (n_869), .B1 (n_1229), .B2 (n_1226));
NAND2_X1 i_844 (.ZN (n_1209), .A1 (p_9[48]), .A2 (n_1211));
NAND2_X1 i_843 (.ZN (n_867), .A1 (n_1212), .A2 (n_1209));
OAI21_X1 i_842 (.ZN (n_863), .A (n_1224), .B1 (n_1231), .B2 (n_1227));
HA_X1 i_841 (.CO (n_753), .S (slo__n1685), .A (n_1182), .B (n_750));
HA_X1 i_840 (.CO (n_1207), .S (slo__n1848), .A (n_763), .B (n_774));
INV_X1 slo__sro_c2718 (.ZN (slo__sro_n1873), .A (n_759));
OAI21_X4 CLOCK_sgo__sro_c3512 (.ZN (n_519), .A (CLOCK_sgo__sro_n2608), .B1 (n_521), .B2 (slo__sro_n587));
FA_X1 i_837 (.CO (n_1203), .S (n_766), .A (p_10[49]), .B (p_11[49]), .CI (p_12[49]));
FA_X1 i_836 (.CO (n_1202), .S (n_770), .A (n_867), .B (n_757), .CI (n_768));
FA_X1 i_835 (.CO (n_1201), .S (n_768), .A (p_13[49]), .B (p_14[49]), .CI (n_755));
FA_X1 i_834 (.CO (n_1200), .S (n_764), .A (n_760), .B (n_762), .CI (n_751));
XNOR2_X2 CLOCK_sgo__sro_c3465 (.ZN (CLOCK_sgo__sro_n2583), .A (n_470), .B (CLOCK_sgo__sro_n2584));
NAND2_X1 slo__sro_c2222 (.ZN (slo__sro_n1540), .A1 (n_496), .A2 (n_494));
INV_X1 slo__sro_c2538 (.ZN (slo__sro_n1737), .A (n_463));
FA_X1 i_830 (.CO (n_747), .S (n_746), .A (n_1177), .B (n_742), .CI (n_740));
FA_X1 i_829 (.CO (n_759), .S (n_758), .A (n_741), .B (n_869), .CI (n_745));
FA_X1 i_828 (.CO (n_745), .S (n_744), .A (n_1179), .B (n_1180), .CI (n_872));
FA_X1 i_827 (.CO (n_741), .S (n_740), .A (p_9[47]), .B (p_10[47]), .CI (p_11[47]));
FA_X1 i_826 (.CO (n_761), .S (n_760), .A (n_756), .B (n_754), .CI (n_865));
FA_X1 i_825 (.CO (n_755), .S (n_754), .A (p_10[48]), .B (p_11[48]), .CI (p_12[48]));
FA_X1 i_824 (.CO (n_757), .S (n_756), .A (p_13[48]), .B (p_14[48]), .CI (n_743));
FA_X1 i_823 (.CO (n_743), .S (n_742), .A (p_12[47]), .B (p_13[47]), .CI (p_14[47]));
INV_X2 i_822 (.ZN (n_1199), .A (n_1129));
INV_X1 i_821 (.ZN (n_1198), .A (p_8[46]));
INV_X1 i_820 (.ZN (n_1197), .A (p_6[45]));
INV_X1 i_819 (.ZN (n_1196), .A (p_7[45]));
NAND3_X4 i_818 (.ZN (n_1195), .A1 (n_1171), .A2 (n_1150), .A3 (n_1169));
NOR2_X4 CLOCK_slo__c3939 (.ZN (CLOCK_slo__n2890), .A1 (slo__sro_n704), .A2 (n_337));
OAI21_X1 i_816 (.ZN (n_1193), .A (n_1170), .B1 (n_1172), .B2 (n_1173));
NOR2_X2 i_815 (.ZN (n_1192), .A1 (slo__sro_n567), .A2 (n_1193));
INV_X1 i_814 (.ZN (n_1191), .A (n_1192));
XNOR2_X1 sgo__sro_c349 (.ZN (n_1017), .A (slo__sro_n1474), .B (sgo__sro_n187));
OAI21_X4 i_812 (.ZN (n_1189), .A (slo__xsl_n1063), .B1 (n_1199), .B2 (opt_ipo_n2168));
NAND2_X2 i_811 (.ZN (n_1188), .A1 (n_1197), .A2 (n_1196));
NAND2_X1 i_810 (.ZN (n_1187), .A1 (n_1183), .A2 (n_1164));
OAI21_X1 i_809 (.ZN (n_1186), .A (n_1187), .B1 (n_1183), .B2 (n_1164));
XNOR2_X1 i_808 (.ZN (\aggregated_res[14] [46] ), .A (n_1189), .B (n_1186));
XOR2_X1 i_807 (.Z (n_1185), .A (p_6[46]), .B (p_7[46]));
XNOR2_X1 i_806 (.ZN (n_870), .A (p_8[46]), .B (n_1185));
FA_X1 i_805 (.CO (n_1184), .S (n_1183), .A (n_734), .B (n_1163), .CI (n_736));
FA_X1 i_804 (.CO (n_1182), .S (n_736), .A (n_1159), .B (n_732), .CI (slo__sro_n1402));
FA_X1 i_803 (.CO (n_1181), .S (n_732), .A (n_1158), .B (n_728), .CI (n_726));
FA_X1 i_802 (.CO (n_1180), .S (n_726), .A (p_9[46]), .B (p_10[46]), .CI (p_11[46]));
FA_X1 i_801 (.CO (n_1179), .S (n_728), .A (p_12[46]), .B (p_13[46]), .CI (p_14[46]));
FA_X1 i_800 (.CO (n_1178), .S (n_734), .A (n_870), .B (n_730), .CI (n_1161));
FA_X1 i_799 (.CO (n_1177), .S (n_730), .A (n_713), .B (n_1157), .CI (n_1188));
FA_X1 i_798 (.CO (n_713), .S (n_1176), .A (p_11[45]), .B (p_12[45]), .CI (p_13[45]));
INV_X1 i_797 (.ZN (n_1175), .A (p_7[44]));
OAI21_X2 i_796 (.ZN (n_1174), .A (n_1149), .B1 (slo__n416), .B2 (n_1151));
NAND2_X1 i_795 (.ZN (n_1173), .A1 (n_1147), .A2 (n_708));
NOR2_X1 i_794 (.ZN (n_1172), .A1 (n_709), .A2 (n_724));
INV_X2 i_793 (.ZN (n_1171), .A (n_1172));
NAND2_X1 i_792 (.ZN (n_1170), .A1 (n_709), .A2 (n_724));
OR2_X2 i_791 (.ZN (n_1169), .A1 (n_708), .A2 (n_1147));
NAND2_X1 i_790 (.ZN (n_1168), .A1 (n_1171), .A2 (n_1170));
NAND2_X1 i_789 (.ZN (n_1167), .A1 (n_1174), .A2 (n_1169));
NAND2_X2 i_788 (.ZN (n_1166), .A1 (n_1167), .A2 (n_1173));
XNOR2_X2 i_787 (.ZN (\aggregated_res[14] [45] ), .A (n_1166), .B (n_1168));
XOR2_X1 i_786 (.Z (n_1165), .A (p_5[44]), .B (p_6[44]));
XNOR2_X1 i_785 (.ZN (n_875), .A (p_7[44]), .B (n_1165));
OAI21_X1 i_784 (.ZN (n_873), .A (n_1188), .B1 (n_1197), .B2 (n_1196));
HA_X1 i_783 (.CO (n_1164), .S (n_724), .A (n_707), .B (n_722));
FA_X1 i_782 (.CO (n_1163), .S (n_722), .A (n_718), .B (n_705), .CI (n_720));
INV_X1 slo__sro_c2073 (.ZN (slo__sro_n1442), .A (n_309));
NAND2_X1 slo__sro_c1942 (.ZN (slo__sro_n1343), .A1 (n_612), .A2 (n_610));
FA_X1 i_779 (.CO (n_1159), .S (n_718), .A (n_710), .B (n_873), .CI (n_714));
FA_X1 i_778 (.CO (n_1158), .S (n_714), .A (p_14[45]), .B (n_697), .CI (n_695));
FA_X1 i_777 (.CO (n_1157), .S (n_710), .A (p_8[45]), .B (p_9[45]), .CI (p_10[45]));
NAND2_X1 slo__sro_c1170 (.ZN (slo__sro_n820), .A1 (n_676), .A2 (n_878));
INV_X1 slo__sro_c2492 (.ZN (slo__sro_n1705), .A (n_1178));
FA_X1 i_774 (.CO (n_705), .S (n_704), .A (n_698), .B (n_1140), .CI (n_700));
FA_X1 i_773 (.CO (n_701), .S (n_700), .A (n_1152), .B (n_1138), .CI (n_696));
FA_X1 i_772 (.CO (n_697), .S (n_696), .A (p_11[44]), .B (p_12[44]), .CI (p_13[44]));
FA_X1 i_771 (.CO (n_699), .S (n_698), .A (p_14[44]), .B (n_1139), .CI (n_1141));
FA_X1 i_770 (.CO (n_703), .S (n_702), .A (n_694), .B (n_875), .CI (n_1142));
FA_X1 i_769 (.CO (n_695), .S (n_694), .A (p_8[44]), .B (p_9[44]), .CI (p_10[44]));
INV_X1 i_768 (.ZN (n_1156), .A (n_1134));
INV_X1 i_767 (.ZN (n_1155), .A (p_5[43]));
INV_X1 i_766 (.ZN (n_1154), .A (p_6[43]));
AOI21_X1 i_765 (.ZN (n_1153), .A (n_1156), .B1 (n_1129), .B2 (n_1133));
NAND2_X1 i_764 (.ZN (n_1152), .A1 (n_1155), .A2 (n_1154));
NOR2_X1 i_763 (.ZN (n_1151), .A1 (n_1092), .A2 (sgo__sro_n16));
INV_X1 i_762 (.ZN (n_1150), .A (slo__n557));
NAND2_X1 i_761 (.ZN (n_1149), .A1 (n_1092), .A2 (sgo__sro_n16));
NAND2_X1 i_760 (.ZN (n_1148), .A1 (n_1150), .A2 (n_1149));
XOR2_X2 i_759 (.Z (\aggregated_res[14] [43] ), .A (n_1153), .B (n_1148));
OAI21_X1 i_758 (.ZN (n_878), .A (n_1152), .B1 (n_1155), .B2 (n_1154));
AOI21_X1 i_757 (.ZN (n_882), .A (n_17), .B1 (p_4[42]), .B2 (n_19));
NAND2_X4 sgo__sro_c135 (.ZN (n_997), .A1 (opt_ipo_n2021), .A2 (n_998));
NAND2_X1 slo__sro_c1217 (.ZN (slo__sro_n849), .A1 (n_20), .A2 (n_51));
NAND2_X1 slo__sro_c1313 (.ZN (slo__sro_n903), .A1 (n_416), .A2 (n_414));
INV_X1 slo__sro_c1191 (.ZN (slo__sro_n835), .A (n_1082));
NAND2_X1 slo__sro_c1205 (.ZN (slo__sro_n842), .A1 (n_688), .A2 (n_684));
FA_X1 i_751 (.CO (n_1141), .S (n_676), .A (p_7[43]), .B (p_8[43]), .CI (p_9[43]));
FA_X1 i_750 (.CO (n_1140), .S (n_684), .A (n_1085), .B (n_680), .CI (n_678));
FA_X1 i_749 (.CO (n_1139), .S (n_678), .A (p_10[43]), .B (p_11[43]), .CI (p_12[43]));
FA_X1 i_748 (.CO (n_1138), .S (n_680), .A (p_13[43]), .B (p_14[43]), .CI (n_1086));
NAND2_X1 slo__sro_c1017 (.ZN (slo__sro_n695), .A1 (n_260), .A2 (slo__sro_n1798));
XNOR2_X1 i_746 (.ZN (\aggregated_res[14] [42] ), .A (n_1129), .B (n_1135));
NAND2_X1 i_745 (.ZN (n_1135), .A1 (n_1133), .A2 (n_1134));
NAND2_X1 i_744 (.ZN (n_1134), .A1 (n_1046), .A2 (n_674));
INV_X1 i_743 (.ZN (n_1133), .A (n_1132));
NOR2_X1 i_742 (.ZN (n_1132), .A1 (n_1046), .A2 (n_674));
OAI21_X4 i_741 (.ZN (n_1129), .A (n_1106), .B1 (n_1123), .B2 (n_1128));
OAI21_X2 i_740 (.ZN (n_1128), .A (n_1122), .B1 (n_1078), .B2 (n_1018));
AOI21_X4 i_739 (.ZN (n_1123), .A (n_1116), .B1 (n_985), .B2 (n_1119));
INV_X1 i_738 (.ZN (n_1122), .A (n_1104));
AOI21_X2 sgo__sro_c475 (.ZN (n_1214), .A (sgo__sro_n255), .B1 (n_1217), .B2 (n_1218));
OR2_X1 sgo__sro_c112 (.ZN (sgo__sro_n75), .A1 (n_793), .A2 (n_711));
NAND2_X4 sgo__sro_c255 (.ZN (n_723), .A1 (n_725), .A2 (sgo__sro_n137));
OAI21_X2 sgo__sro_c113 (.ZN (n_839), .A (sgo__sro_n75), .B1 (n_799), .B2 (n_801));
AND2_X2 i_733 (.ZN (n_1109), .A1 (n_946), .A2 (n_1000));
NAND2_X1 i_732 (.ZN (n_1108), .A1 (n_1017), .A2 (slo__sro_n466));
INV_X2 i_731 (.ZN (n_1106), .A (sgo__sro_n54));
NAND2_X2 CLOCK_sgo__sro_c3686 (.ZN (CLOCK_sgo__sro_n2704), .A1 (CLOCK_sgo__sro_n2706), .A2 (CLOCK_sgo__sro_n2705));
NAND3_X4 i_729 (.ZN (n_1104), .A1 (n_1095), .A2 (n_1075), .A3 (n_1058));
AOI21_X1 i_728 (.ZN (n_1103), .A (n_1097), .B1 (n_1078), .B2 (n_1018));
NAND3_X1 i_727 (.ZN (n_1102), .A1 (n_1033), .A2 (n_1070), .A3 (n_1058));
INV_X1 i_726 (.ZN (n_1097), .A (n_1096));
NAND2_X1 i_725 (.ZN (n_1096), .A1 (n_1069), .A2 (n_595));
INV_X1 i_724 (.ZN (n_1095), .A (n_1094));
NOR2_X1 i_723 (.ZN (n_1094), .A1 (n_595), .A2 (n_1069));
XOR2_X1 i_722 (.Z (n_880), .A (n_1093), .B (p_4[42]));
XNOR2_X1 i_721 (.ZN (n_1093), .A (p_6[42]), .B (p_5[42]));
INV_X1 slo__sro_c1535 (.ZN (slo__sro_n1046), .A (n_668));
NAND2_X1 slo__sro_c1633 (.ZN (slo__sro_n1108), .A1 (slo__sro_n1130), .A2 (n_632));
NAND2_X1 slo__sro_c1521 (.ZN (slo__sro_n1034), .A1 (slo__sro_n1040), .A2 (n_1043));
FA_X1 i_717 (.CO (n_1087), .S (n_666), .A (n_1034), .B (n_662), .CI (n_660));
FA_X1 i_716 (.CO (n_1086), .S (n_660), .A (p_10[42]), .B (p_11[42]), .CI (p_12[42]));
FA_X1 i_715 (.CO (n_1085), .S (n_662), .A (p_13[42]), .B (p_14[42]), .CI (n_1036));
FA_X1 i_714 (.CO (n_1084), .S (n_668), .A (n_658), .B (n_880), .CI (n_664));
FA_X1 i_713 (.CO (n_1082), .S (n_664), .A (n_1038), .B (n_1041), .CI (n_1060));
FA_X1 i_712 (.CO (n_1079), .S (n_658), .A (p_7[42]), .B (p_8[42]), .CI (p_9[42]));
INV_X1 slo__sro_c1409 (.ZN (slo__sro_n968), .A (n_1015));
NOR2_X4 i_710 (.ZN (n_1077), .A1 (n_1033), .A2 (n_1070));
INV_X4 i_709 (.ZN (n_1075), .A (n_1077));
NOR2_X2 CLOCK_sgo__c3790 (.ZN (CLOCK_sgo__n2761), .A1 (n_982), .A2 (n_1022));
INV_X1 slo__sro_c1503 (.ZN (slo__sro_n1025), .A (n_1042));
INV_X1 i_706 (.ZN (n_1066), .A (p_3[40]));
INV_X1 i_705 (.ZN (n_1065), .A (p_3[39]));
INV_X1 i_704 (.ZN (n_1064), .A (p_4[41]));
INV_X1 i_703 (.ZN (n_1063), .A (p_4[39]));
INV_X1 i_702 (.ZN (n_1062), .A (p_5[41]));
INV_X1 i_701 (.ZN (n_1061), .A (p_2[38]));
NAND2_X1 i_700 (.ZN (n_1060), .A1 (n_1064), .A2 (n_1062));
NAND2_X1 slo__sro_c2407 (.ZN (slo__sro_n1646), .A1 (n_514), .A2 (n_487));
NAND2_X1 i_698 (.ZN (n_1057), .A1 (n_637), .A2 (n_656));
NAND2_X1 i_697 (.ZN (n_1056), .A1 (n_1058), .A2 (n_1057));
NAND2_X1 i_696 (.ZN (n_889), .A1 (n_1065), .A2 (n_1063));
OAI21_X1 i_695 (.ZN (n_888), .A (n_889), .B1 (n_1065), .B2 (n_1063));
NAND2_X1 i_694 (.ZN (n_1055), .A1 (p_3[38]), .A2 (n_1061));
INV_X1 i_693 (.ZN (n_1054), .A (n_1055));
OAI22_X1 i_692 (.ZN (n_1053), .A1 (p_3[38]), .A2 (n_1061), .B1 (n_1054), .B2 (p_4[38]));
INV_X1 i_691 (.ZN (n_892), .A (n_1053));
NAND2_X1 i_690 (.ZN (n_1052), .A1 (n_1066), .A2 (p_5[40]));
OR2_X1 i_689 (.ZN (n_1051), .A1 (n_1066), .A2 (p_5[40]));
NAND2_X1 i_688 (.ZN (n_1050), .A1 (n_1052), .A2 (n_1051));
XNOR2_X1 i_687 (.ZN (n_885), .A (p_4[40]), .B (n_1050));
OAI21_X1 i_686 (.ZN (n_1049), .A (n_1055), .B1 (p_3[38]), .B2 (n_1061));
XNOR2_X1 i_684 (.ZN (n_890), .A (p_4[38]), .B (n_1049));
NAND2_X1 i_683 (.ZN (n_1048), .A1 (p_4[40]), .A2 (n_1051));
NAND2_X1 i_682 (.ZN (n_887), .A1 (n_1052), .A2 (n_1048));
OAI21_X1 i_681 (.ZN (n_883), .A (n_1060), .B1 (n_1064), .B2 (n_1062));
HA_X1 i_680 (.CO (n_1046), .S (n_656), .A (slo__sro_n1132), .B (n_654));
NOR2_X2 slo__c2384 (.ZN (slo__n1633), .A1 (n_637), .A2 (n_656));
INV_X1 slo__sro_c2354 (.ZN (slo__sro_n1615), .A (n_597));
FA_X1 i_677 (.CO (n_1042), .S (n_648), .A (n_640), .B (n_638), .CI (n_883));
FA_X1 i_676 (.CO (n_1041), .S (n_638), .A (p_6[41]), .B (p_7[41]), .CI (p_8[41]));
FA_X1 i_675 (.CO (n_1038), .S (n_640), .A (p_9[41]), .B (p_10[41]), .CI (p_11[41]));
FA_X1 i_673 (.CO (n_1037), .S (n_646), .A (n_887), .B (slo__sro_n1612), .CI (n_642));
FA_X1 i_672 (.CO (n_1036), .S (n_642), .A (p_12[41]), .B (p_13[41]), .CI (p_14[41]));
FA_X1 i_671 (.CO (n_1035), .S (n_650), .A (n_644), .B (n_629), .CI (n_627));
FA_X1 i_670 (.CO (n_1034), .S (n_644), .A (n_623), .B (n_621), .CI (n_619));
NAND2_X1 slo__sro_c1654 (.ZN (slo__sro_n1122), .A1 (n_892), .A2 (n_575));
NAND2_X1 slo__sro_c1958 (.ZN (slo__sro_n1359), .A1 (n_1012), .A2 (n_1010));
INV_X1 CLOCK_sgo__sro_c3463 (.ZN (CLOCK_sgo__sro_n2584), .A (n_832));
INV_X1 slo__sro_c1693 (.ZN (slo__sro_n1155), .A (slo__sro_n1357));
FA_X1 i_665 (.CO (n_613), .S (n_612), .A (n_587), .B (n_606), .CI (slo__sro_n1150));
NAND2_X1 slo__sro_c2004 (.ZN (slo__sro_n1396), .A1 (n_965), .A2 (n_897));
FA_X1 i_663 (.CO (n_631), .S (n_630), .A (n_605), .B (n_624), .CI (n_607));
FA_X1 i_662 (.CO (n_607), .S (n_606), .A (n_600), .B (n_598), .CI (n_596));
NAND2_X1 slo__sro_c2368 (.ZN (slo__sro_n1624), .A1 (n_652), .A2 (n_650));
FA_X1 i_660 (.CO (n_597), .S (n_596), .A (p_5[39]), .B (p_6[39]), .CI (p_7[39]));
FA_X1 i_659 (.CO (n_599), .S (n_598), .A (p_8[39]), .B (p_9[39]), .CI (p_10[39]));
FA_X1 i_658 (.CO (n_601), .S (n_600), .A (p_11[39]), .B (p_12[39]), .CI (p_13[39]));
FA_X1 i_657 (.CO (n_611), .S (n_610), .A (n_602), .B (n_585), .CI (n_589));
FA_X1 i_656 (.CO (n_589), .S (n_1028), .A (n_580), .B (n_1011), .CI (n_1005));
FA_X1 i_655 (.CO (n_585), .S (n_584), .A (n_1004), .B (n_578), .CI (n_576));
FA_X1 i_654 (.CO (n_633), .S (n_632), .A (n_626), .B (slo__sro_n1152), .CI (n_628));
FA_X1 i_653 (.CO (n_629), .S (n_628), .A (n_620), .B (n_618), .CI (n_885));
FA_X1 i_652 (.CO (n_619), .S (n_618), .A (p_6[40]), .B (p_7[40]), .CI (p_8[40]));
FA_X1 i_651 (.CO (n_621), .S (n_620), .A (p_9[40]), .B (p_10[40]), .CI (p_11[40]));
AND2_X2 slo__sro_c1707 (.ZN (slo__sro_n1166), .A1 (n_1040), .A2 (n_1370));
INV_X1 slo__sro_c1668 (.ZN (slo__sro_n1135), .A (n_611));
FA_X1 i_648 (.CO (n_581), .S (n_580), .A (p_14[38]), .B (n_1008), .CI (n_1009));
FA_X1 i_647 (.CO (n_575), .S (n_574), .A (p_5[38]), .B (p_6[38]), .CI (p_7[38]));
INV_X1 slo__sro_c1970 (.ZN (slo__sro_n1372), .A (n_1014));
FA_X1 i_645 (.CO (n_627), .S (n_626), .A (n_889), .B (n_603), .CI (n_622));
FA_X1 i_644 (.CO (n_623), .S (n_622), .A (p_12[40]), .B (p_13[40]), .CI (p_14[40]));
FA_X1 i_643 (.CO (n_603), .S (n_602), .A (p_14[39]), .B (n_579), .CI (n_577));
FA_X1 i_642 (.CO (n_577), .S (n_576), .A (p_8[38]), .B (p_9[38]), .CI (p_10[38]));
FA_X1 i_641 (.CO (n_579), .S (n_578), .A (p_11[38]), .B (p_12[38]), .CI (p_13[38]));
INV_X1 i_640 (.ZN (n_1027), .A (p_2[37]));
INV_X1 i_639 (.ZN (n_1025), .A (p_2[36]));
INV_X1 i_638 (.ZN (n_1024), .A (p_3[37]));
NAND2_X1 i_637 (.ZN (n_1023), .A1 (n_1027), .A2 (n_1024));
NOR2_X4 i_636 (.ZN (n_1022), .A1 (slo__sro_n466), .A2 (n_1017));
AOI21_X2 i_635 (.ZN (n_1021), .A (n_979), .B1 (n_980), .B2 (n_978));
AOI21_X1 i_634 (.ZN (n_1020), .A (n_1022), .B1 (n_1017), .B2 (slo__sro_n466));
XOR2_X2 i_633 (.Z (\aggregated_res[14] [37] ), .A (n_1021), .B (n_1020));
OAI21_X1 i_632 (.ZN (n_893), .A (n_1023), .B1 (n_1027), .B2 (n_1024));
AOI21_X1 i_631 (.ZN (n_1019), .A (p_3[36]), .B1 (p_2[36]), .B2 (n_21));
AOI21_X1 i_630 (.ZN (n_897), .A (n_1019), .B1 (n_1025), .B2 (p_1[36]));
NOR2_X2 sgo__c378 (.ZN (sgo__n199), .A1 (opt_ipo_n1967), .A2 (n_636));
INV_X1 slo__sro_c2152 (.ZN (slo__sro_n1497), .A (n_973));
FA_X1 i_626 (.CO (n_1014), .S (n_564), .A (n_893), .B (slo__sro_n1393), .CI (n_967));
INV_X1 slo__sro_c2016 (.ZN (slo__sro_n1405), .A (n_703));
FA_X1 i_624 (.CO (n_1011), .S (n_562), .A (n_554), .B (n_552), .CI (n_550));
FA_X1 i_623 (.CO (n_1010), .S (n_550), .A (p_4[37]), .B (p_5[37]), .CI (p_6[37]));
FA_X1 i_622 (.CO (n_1009), .S (n_552), .A (p_7[37]), .B (p_8[37]), .CI (p_9[37]));
FA_X1 i_621 (.CO (n_1008), .S (n_554), .A (p_10[37]), .B (p_11[37]), .CI (p_12[37]));
FA_X1 i_620 (.CO (n_1006), .S (n_566), .A (n_972), .B (n_560), .CI (n_969));
FA_X1 i_619 (.CO (n_1005), .S (n_560), .A (n_968), .B (n_971), .CI (n_556));
FA_X1 i_618 (.CO (n_1004), .S (n_556), .A (p_13[37]), .B (p_14[37]), .CI (n_964));
INV_X1 i_617 (.ZN (n_1001), .A (n_954));
NAND2_X2 i_616 (.ZN (n_1000), .A1 (n_938), .A2 (n_896));
OAI21_X2 i_615 (.ZN (n_999), .A (n_844), .B1 (n_711), .B2 (n_793));
INV_X1 i_614 (.ZN (n_998), .A (n_999));
NOR2_X1 sgo__sro_c171 (.ZN (sgo__sro_n102), .A1 (n_1183), .A2 (n_1164));
OR2_X1 sgo__sro_c474 (.ZN (sgo__sro_n255), .A1 (n_1220), .A2 (n_1216));
OAI21_X4 i_611 (.ZN (n_995), .A (opt_ipo_n2338), .B1 (n_996), .B2 (opt_ipo_n1965));
NOR2_X4 i_609 (.ZN (n_990), .A1 (opt_ipo_n1905), .A2 (n_723));
AOI21_X4 i_608 (.ZN (n_989), .A (n_801), .B1 (opt_ipo_n1924), .B2 (n_663));
OAI21_X2 i_607 (.ZN (n_987), .A (n_841), .B1 (n_989), .B2 (n_999));
OAI21_X4 i_606 (.ZN (n_986), .A (n_987), .B1 (CLOCK_sgo__sro_n2583), .B2 (n_833));
OAI211_X4 i_605 (.ZN (n_985), .A (n_908), .B (n_986), .C1 (n_997), .C2 (n_990));
INV_X1 i_604 (.ZN (n_983), .A (n_985));
NOR2_X2 i_603 (.ZN (n_982), .A1 (n_938), .A2 (n_896));
OAI21_X4 i_602 (.ZN (n_981), .A (n_1000), .B1 (n_983), .B2 (n_982));
OAI21_X4 i_601 (.ZN (n_980), .A (n_1001), .B1 (n_981), .B2 (n_945));
NOR2_X4 i_600 (.ZN (n_979), .A1 (slo__sro_n464), .A2 (n_937));
NAND2_X2 i_599 (.ZN (n_978), .A1 (n_937), .A2 (slo__sro_n464));
OAI21_X1 i_598 (.ZN (n_977), .A (n_978), .B1 (n_937), .B2 (slo__sro_n464));
XOR2_X2 i_597 (.Z (\aggregated_res[14] [36] ), .A (n_980), .B (n_977));
XOR2_X1 i_596 (.Z (n_976), .A (p_3[36]), .B (p_2[36]));
XNOR2_X1 i_595 (.ZN (n_895), .A (p_1[36]), .B (n_976));
INV_X1 slo__sro_c810 (.ZN (slo__sro_n499), .A (n_1026));
FA_X1 i_593 (.CO (n_974), .S (n_546), .A (n_921), .B (n_542), .CI (slo__sro_n1255));
FA_X1 i_592 (.CO (n_973), .S (n_542), .A (n_928), .B (n_920), .CI (n_536));
FA_X1 i_591 (.CO (n_972), .S (n_536), .A (n_957), .B (n_933), .CI (n_532));
FA_X1 i_590 (.CO (n_971), .S (n_532), .A (p_13[36]), .B (p_14[36]), .CI (n_923));
FA_X1 i_589 (.CO (n_970), .S (n_544), .A (n_934), .B (n_538), .CI (n_540));
FA_X1 i_588 (.CO (n_969), .S (n_540), .A (n_895), .B (n_929), .CI (n_534));
FA_X1 i_587 (.CO (n_968), .S (n_534), .A (n_924), .B (n_925), .CI (n_919));
FA_X1 i_586 (.CO (n_967), .S (n_538), .A (n_530), .B (n_528), .CI (n_526));
FA_X1 i_585 (.CO (n_966), .S (n_526), .A (p_4[36]), .B (p_5[36]), .CI (p_6[36]));
FA_X1 i_584 (.CO (n_965), .S (n_528), .A (p_7[36]), .B (p_8[36]), .CI (p_9[36]));
FA_X1 i_583 (.CO (n_964), .S (n_530), .A (p_10[36]), .B (p_11[36]), .CI (p_12[36]));
INV_X1 i_582 (.ZN (n_963), .A (p_1[35]));
INV_X1 i_581 (.ZN (n_962), .A (p_1[34]));
INV_X1 i_580 (.ZN (n_960), .A (p_2[35]));
NAND2_X1 i_579 (.ZN (n_957), .A1 (n_963), .A2 (n_960));
NOR2_X4 i_578 (.ZN (n_954), .A1 (n_524), .A2 (slo__sro_n1538));
NAND2_X1 i_577 (.ZN (n_946), .A1 (n_524), .A2 (slo__sro_n1538));
INV_X1 i_576 (.ZN (n_945), .A (n_946));
NOR2_X1 i_575 (.ZN (n_944), .A1 (n_954), .A2 (n_945));
OAI21_X1 i_574 (.ZN (n_898), .A (n_957), .B1 (n_963), .B2 (n_960));
NOR2_X1 i_573 (.ZN (n_942), .A1 (n_962), .A2 (p_0[34]));
AOI21_X1 i_572 (.ZN (n_940), .A (n_942), .B1 (n_962), .B2 (p_0[34]));
XOR2_X1 i_571 (.Z (n_900), .A (p_2[34]), .B (n_940));
NOR2_X1 i_570 (.ZN (n_939), .A1 (p_2[34]), .A2 (n_942));
AOI21_X1 i_569 (.ZN (n_902), .A (n_939), .B1 (n_962), .B2 (p_0[34]));
NAND2_X1 slo__sro_c2239 (.ZN (slo__sro_n1550), .A1 (n_492), .A2 (n_886));
HA_X1 i_567 (.CO (n_937), .S (n_524), .A (slo__sro_n1548), .B (slo__sro_n1267));
INV_X1 slo__sro_c1853 (.ZN (slo__sro_n1282), .A (n_174));
NAND2_X1 slo__sro_c1841 (.ZN (slo__sro_n1270), .A1 (n_518), .A2 (n_495));
FA_X1 i_564 (.CO (n_934), .S (n_516), .A (n_510), .B (n_508), .CI (n_489));
FA_X1 i_563 (.CO (n_933), .S (n_508), .A (n_481), .B (n_479), .CI (n_477));
FA_X1 i_562 (.CO (n_929), .S (n_510), .A (n_475), .B (n_902), .CI (n_483));
FA_X1 i_561 (.CO (n_928), .S (n_512), .A (n_506), .B (n_504), .CI (n_502));
FA_X1 i_560 (.CO (n_925), .S (n_502), .A (p_6[35]), .B (p_7[35]), .CI (p_8[35]));
FA_X1 i_559 (.CO (n_924), .S (n_504), .A (p_9[35]), .B (p_10[35]), .CI (p_11[35]));
FA_X1 i_558 (.CO (n_923), .S (n_506), .A (p_12[35]), .B (p_13[35]), .CI (p_14[35]));
FA_X1 i_557 (.CO (n_495), .S (n_494), .A (n_488), .B (n_486), .CI (n_490));
FA_X1 i_556 (.CO (n_489), .S (n_488), .A (n_476), .B (n_474), .CI (n_900));
FA_X1 i_555 (.CO (n_475), .S (n_474), .A (p_3[34]), .B (p_4[34]), .CI (p_5[34]));
FA_X1 i_554 (.CO (n_477), .S (n_476), .A (p_6[34]), .B (p_7[34]), .CI (p_8[34]));
INV_X1 slo__sro_c2419 (.ZN (slo__sro_n1655), .A (n_482));
FA_X1 i_552 (.CO (n_920), .S (n_514), .A (n_500), .B (n_898), .CI (n_485));
FA_X1 i_551 (.CO (n_919), .S (n_500), .A (p_3[35]), .B (p_4[35]), .CI (p_5[35]));
INV_X1 slo__sro_c2437 (.ZN (slo__sro_n1665), .A (n_877));
FA_X1 i_549 (.CO (n_483), .S (n_482), .A (n_859), .B (n_864), .CI (n_866));
BUF_X2 slo__c2475 (.Z (n_1208), .A (slo__n1685));
FA_X1 i_547 (.CO (n_487), .S (n_486), .A (n_881), .B (n_480), .CI (n_478));
FA_X1 i_546 (.CO (n_479), .S (n_478), .A (p_9[34]), .B (p_10[34]), .CI (p_11[34]));
FA_X1 i_545 (.CO (n_481), .S (n_480), .A (p_12[34]), .B (p_13[34]), .CI (p_14[34]));
NAND2_X1 slo__sro_c2276 (.ZN (slo__sro_n1572), .A1 (p_6[14]), .A2 (p_15[14]));
FA_X1 i_543 (.CO (n_493), .S (n_492), .A (n_861), .B (n_884), .CI (n_879));
INV_X1 i_542 (.ZN (n_917), .A (p_0[33]));
INV_X1 i_541 (.ZN (n_916), .A (p_1[33]));
INV_X1 i_540 (.ZN (n_911), .A (n_844));
NAND2_X1 i_539 (.ZN (n_909), .A1 (n_917), .A2 (n_916));
NAND2_X1 i_538 (.ZN (n_908), .A1 (CLOCK_sgo__sro_n2583), .A2 (n_833));
OAI21_X1 i_537 (.ZN (n_906), .A (n_908), .B1 (CLOCK_sgo__sro_n2583), .B2 (n_833));
AOI21_X2 i_536 (.ZN (n_904), .A (n_911), .B1 (n_839), .B2 (n_841));
XNOR2_X2 i_535 (.ZN (\aggregated_res[14] [33] ), .A (n_904), .B (n_906));
NAND2_X1 i_534 (.ZN (n_901), .A1 (n_851), .A2 (n_779));
OAI21_X1 i_533 (.ZN (n_899), .A (p_14[32]), .B1 (n_851), .B2 (n_779));
NAND2_X1 i_532 (.ZN (n_905), .A1 (n_901), .A2 (n_899));
OAI21_X1 i_531 (.ZN (n_903), .A (n_909), .B1 (n_917), .B2 (n_916));
OR2_X1 CLOCK_sgo__sro_c3511 (.ZN (CLOCK_sgo__sro_n2608), .A1 (n_405), .A2 (n_411));
FA_X1 i_529 (.CO (n_891), .S (n_470), .A (n_466), .B (n_831), .CI (n_468));
FA_X1 i_528 (.CO (n_886), .S (n_468), .A (n_462), .B (n_464), .CI (n_813));
FA_X1 i_527 (.CO (n_884), .S (n_464), .A (n_454), .B (n_812), .CI (n_822));
FA_X1 i_526 (.CO (n_881), .S (n_454), .A (p_14[33]), .B (n_814), .CI (n_818));
FA_X1 i_525 (.CO (n_879), .S (n_462), .A (n_903), .B (n_807), .CI (n_456));
FA_X1 i_524 (.CO (n_877), .S (n_456), .A (n_809), .B (n_811), .CI (n_846));
FA_X1 i_523 (.CO (n_876), .S (n_466), .A (n_458), .B (n_829), .CI (n_460));
FA_X1 i_522 (.CO (n_874), .S (n_460), .A (n_450), .B (n_448), .CI (n_446));
FA_X1 i_521 (.CO (n_871), .S (n_446), .A (p_2[33]), .B (p_3[33]), .CI (p_4[33]));
FA_X1 i_520 (.CO (n_866), .S (n_448), .A (p_5[33]), .B (p_6[33]), .CI (p_7[33]));
FA_X1 i_519 (.CO (n_864), .S (n_450), .A (p_8[33]), .B (p_9[33]), .CI (p_10[33]));
FA_X1 i_518 (.CO (n_861), .S (n_458), .A (n_828), .B (n_905), .CI (n_452));
FA_X1 i_517 (.CO (n_859), .S (n_452), .A (p_11[33]), .B (p_12[33]), .CI (p_13[33]));
INV_X1 i_516 (.ZN (n_856), .A (p_0[32]));
INV_X1 i_515 (.ZN (n_854), .A (p_1[32]));
INV_X1 i_514 (.ZN (n_851), .A (p_15[32]));
NAND2_X1 i_513 (.ZN (n_846), .A1 (n_856), .A2 (n_854));
NOR3_X2 sgo__c185 (.ZN (sgo__n107), .A1 (n_1022), .A2 (n_979), .A3 (n_954));
NAND2_X1 i_511 (.ZN (n_841), .A1 (n_795), .A2 (n_444));
INV_X1 CLOCK_slo__xsl_c3842 (.ZN (CLOCK_slo__xsl_n2800), .A (CLOCK_slo__xsl_n2801));
NAND2_X1 i_509 (.ZN (n_836), .A1 (n_844), .A2 (n_841));
XOR2_X2 i_508 (.Z (\aggregated_res[14] [32] ), .A (n_839), .B (n_836));
OAI21_X1 i_507 (.ZN (n_910), .A (n_846), .B1 (n_856), .B2 (n_854));
XOR2_X1 i_506 (.Z (n_835), .A (n_779), .B (p_14[32]));
XNOR2_X1 i_505 (.ZN (n_907), .A (n_835), .B (p_15[32]));
INV_X1 sgo__sro_c172 (.ZN (sgo__sro_n101), .A (sgo__sro_n102));
INV_X1 slo__sro_c1760 (.ZN (slo__sro_n1212), .A (n_685));
FA_X1 i_502 (.CO (n_831), .S (n_440), .A (n_432), .B (n_783), .CI (n_436));
FA_X1 i_501 (.CO (n_829), .S (n_436), .A (n_428), .B (n_776), .CI (n_781));
FA_X1 i_500 (.CO (n_828), .S (n_428), .A (n_771), .B (n_773), .CI (n_775));
FA_X1 i_499 (.CO (n_822), .S (n_432), .A (n_907), .B (n_426), .CI (n_424));
FA_X1 i_498 (.CO (n_818), .S (n_424), .A (p_8[32]), .B (p_9[32]), .CI (p_10[32]));
FA_X1 i_497 (.CO (n_814), .S (n_426), .A (p_11[32]), .B (p_12[32]), .CI (p_13[32]));
FA_X1 i_496 (.CO (n_813), .S (n_438), .A (n_430), .B (n_789), .CI (n_434));
FA_X1 i_495 (.CO (n_812), .S (n_434), .A (n_422), .B (n_420), .CI (n_910));
FA_X1 i_494 (.CO (n_811), .S (n_420), .A (p_2[32]), .B (p_3[32]), .CI (p_4[32]));
FA_X1 i_493 (.CO (n_809), .S (n_422), .A (p_5[32]), .B (p_6[32]), .CI (p_7[32]));
FA_X1 i_492 (.CO (n_807), .S (n_430), .A (n_785), .B (n_786), .CI (n_787));
XNOR2_X1 i_491 (.ZN (\aggregated_res[14] [31] ), .A (n_799), .B (n_805));
OAI21_X1 i_490 (.ZN (n_805), .A (slo__xsl_n988), .B1 (n_793), .B2 (n_711));
NAND2_X1 slo__sro_c1505 (.ZN (slo__sro_n1023), .A1 (n_1037), .A2 (n_1042));
NAND2_X1 slo__sro_c1507 (.ZN (slo__sro_n1021), .A1 (n_1035), .A2 (slo__sro_n1022));
NAND2_X2 i_487 (.ZN (n_799), .A1 (n_797), .A2 (n_715));
OAI21_X1 i_486 (.ZN (n_797), .A (n_717), .B1 (n_663), .B2 (opt_ipo_n1924));
INV_X1 slo__sro_c1325 (.ZN (slo__sro_n910), .A (n_322));
FA_X1 i_484 (.CO (n_791), .S (n_416), .A (n_412), .B (n_410), .CI (n_687));
FA_X1 i_483 (.CO (n_789), .S (n_410), .A (n_392), .B (n_404), .CI (n_402));
FA_X1 i_482 (.CO (n_787), .S (n_402), .A (p_15[31]), .B (n_675), .CI (n_677));
FA_X1 i_481 (.CO (n_786), .S (n_404), .A (n_667), .B (n_669), .CI (n_671));
FA_X1 i_480 (.CO (n_785), .S (n_392), .A (p_0[31]), .B (p_1[31]), .CI (p_2[31]));
FA_X1 i_479 (.CO (n_783), .S (n_412), .A (n_673), .B (n_679), .CI (n_406));
FA_X1 i_478 (.CO (n_781), .S (n_406), .A (n_681), .B (n_683), .CI (slo__sro_n1241));
NAND2_X1 slo__sro_c1827 (.ZN (slo__sro_n1258), .A1 (n_493), .A2 (n_512));
NAND2_X1 slo__sro_c1808 (.ZN (slo__sro_n1244), .A1 (p_12[31]), .A2 (p_13[31]));
FA_X1 i_475 (.CO (n_776), .S (n_408), .A (n_398), .B (n_396), .CI (n_394));
FA_X1 i_474 (.CO (n_775), .S (n_394), .A (p_3[31]), .B (p_4[31]), .CI (p_5[31]));
FA_X1 i_473 (.CO (n_773), .S (n_396), .A (p_6[31]), .B (p_7[31]), .CI (p_8[31]));
FA_X1 i_472 (.CO (n_771), .S (n_398), .A (p_9[31]), .B (p_10[31]), .CI (p_11[31]));
XNOR2_X2 slo__sro_c1317 (.ZN (n_793), .A (slo__sro_n901), .B (n_416));
NAND2_X1 slo__sro_c1315 (.ZN (n_795), .A1 (slo__sro_n902), .A2 (slo__sro_n903));
NOR2_X2 i_468 (.ZN (n_752), .A1 (n_336), .A2 (slo__sro_n1747));
INV_X2 i_467 (.ZN (n_739), .A (n_752));
AND2_X1 slo__sro_c618 (.ZN (slo__sro_n333), .A1 (n_1072), .A2 (n_1096));
NOR2_X2 slo__c736 (.ZN (slo__n419), .A1 (slo__sro_n692), .A2 (n_555));
OR2_X2 i_464 (.ZN (n_735), .A1 (n_590), .A2 (n_553));
NAND2_X1 i_463 (.ZN (n_733), .A1 (n_665), .A2 (n_592));
NAND2_X1 i_461 (.ZN (n_729), .A1 (slo__sro_n704), .A2 (n_337));
NAND2_X1 i_460 (.ZN (n_727), .A1 (n_336), .A2 (slo__sro_n1747));
OAI21_X4 i_459 (.ZN (n_725), .A (slo__n638), .B1 (opt_ipo_n2117), .B2 (opt_ipo_n2154));
INV_X1 sgo__sro_c347 (.ZN (sgo__sro_n187), .A (n_974));
INV_X1 i_457 (.ZN (n_721), .A (n_723));
NAND2_X1 i_456 (.ZN (n_719), .A1 (n_616), .A2 (n_735));
OAI21_X2 i_455 (.ZN (n_717), .A (n_721), .B1 (n_719), .B2 (slo__xsl_n395));
NAND2_X1 i_454 (.ZN (n_715), .A1 (n_663), .A2 (opt_ipo_n1924));
OAI21_X1 i_453 (.ZN (n_712), .A (n_715), .B1 (n_663), .B2 (opt_ipo_n1924));
XNOR2_X1 i_452 (.ZN (\aggregated_res[14] [30] ), .A (n_717), .B (n_712));
HA_X1 i_451 (.CO (n_711), .S (n_693), .A (n_386), .B (slo__sro_n915));
NAND2_X1 slo__sro_c1351 (.ZN (slo__sro_n931), .A1 (n_331), .A2 (n_356));
FA_X1 i_449 (.CO (n_689), .S (n_384), .A (n_353), .B (n_355), .CI (n_357));
FA_X1 i_448 (.CO (n_325), .S (n_324), .A (n_289), .B (n_299), .CI (n_297));
FA_X1 i_447 (.CO (n_297), .S (n_296), .A (p_12[27]), .B (p_15[27]), .CI (n_567));
FA_X1 i_446 (.CO (n_299), .S (n_298), .A (n_557), .B (n_559), .CI (n_561));
FA_X1 i_445 (.CO (n_289), .S (n_288), .A (p_0[27]), .B (p_1[27]), .CI (p_2[27]));
FA_X1 i_444 (.CO (n_687), .S (n_386), .A (n_380), .B (n_378), .CI (n_382));
FA_X1 i_443 (.CO (n_685), .S (n_382), .A (n_351), .B (n_376), .CI (n_374));
FA_X1 i_442 (.CO (n_683), .S (n_374), .A (p_15[30]), .B (n_347), .CI (n_345));
FA_X1 i_441 (.CO (n_345), .S (n_344), .A (p_9[29]), .B (p_10[29]), .CI (p_11[29]));
FA_X1 i_440 (.CO (n_347), .S (n_346), .A (p_12[29]), .B (p_13[29]), .CI (p_15[29]));
FA_X1 i_439 (.CO (n_681), .S (n_376), .A (n_343), .B (n_341), .CI (n_339));
FA_X1 i_438 (.CO (n_339), .S (n_338), .A (p_0[29]), .B (p_1[29]), .CI (p_2[29]));
FA_X1 i_437 (.CO (n_341), .S (n_340), .A (p_3[29]), .B (p_4[29]), .CI (p_5[29]));
FA_X1 i_436 (.CO (n_343), .S (n_342), .A (p_6[29]), .B (p_7[29]), .CI (p_8[29]));
FA_X1 i_435 (.CO (n_351), .S (n_350), .A (n_315), .B (n_313), .CI (n_323));
NAND2_X1 slo__sro_c1385 (.ZN (slo__sro_n954), .A1 (n_326), .A2 (n_328));
FA_X1 i_433 (.CO (n_291), .S (n_290), .A (p_3[27]), .B (p_4[27]), .CI (p_5[27]));
FA_X1 i_432 (.CO (n_293), .S (n_292), .A (p_6[27]), .B (p_7[27]), .CI (p_8[27]));
FA_X1 i_431 (.CO (n_295), .S (n_294), .A (p_9[27]), .B (p_10[27]), .CI (p_11[27]));
FA_X1 i_430 (.CO (n_313), .S (n_312), .A (p_0[28]), .B (p_1[28]), .CI (p_2[28]));
FA_X1 i_429 (.CO (n_315), .S (n_314), .A (p_3[28]), .B (p_4[28]), .CI (p_5[28]));
FA_X1 i_428 (.CO (n_679), .S (n_378), .A (n_349), .B (n_372), .CI (n_370));
FA_X1 i_427 (.CO (n_677), .S (n_370), .A (p_9[30]), .B (p_10[30]), .CI (p_11[30]));
FA_X1 i_426 (.CO (n_675), .S (n_372), .A (p_12[30]), .B (p_13[30]), .CI (p_14[30]));
FA_X1 i_425 (.CO (n_349), .S (n_348), .A (n_321), .B (n_319), .CI (n_317));
FA_X1 i_424 (.CO (n_317), .S (n_316), .A (p_6[28]), .B (p_7[28]), .CI (p_8[28]));
FA_X1 i_423 (.CO (n_319), .S (n_318), .A (p_9[28]), .B (p_10[28]), .CI (p_11[28]));
FA_X1 i_422 (.CO (n_321), .S (n_320), .A (p_12[28]), .B (p_13[28]), .CI (p_15[28]));
FA_X1 i_421 (.CO (n_673), .S (n_380), .A (n_368), .B (n_366), .CI (n_364));
FA_X1 i_420 (.CO (n_671), .S (n_364), .A (p_0[30]), .B (p_1[30]), .CI (p_2[30]));
FA_X1 i_419 (.CO (n_669), .S (n_366), .A (p_3[30]), .B (p_4[30]), .CI (p_5[30]));
FA_X1 i_418 (.CO (n_667), .S (n_368), .A (p_6[30]), .B (p_7[30]), .CI (p_8[30]));
INV_X1 slo__sro_c2572 (.ZN (slo__sro_n1762), .A (n_139));
FA_X1 i_416 (.CO (n_303), .S (n_302), .A (n_294), .B (n_292), .CI (n_290));
FA_X1 i_415 (.CO (n_301), .S (n_300), .A (n_572), .B (n_565), .CI (n_296));
HA_X1 i_414 (.CO (n_337), .S (n_336), .A (slo__sro_n951), .B (n_334));
FA_X1 i_413 (.CO (n_327), .S (n_326), .A (n_320), .B (n_318), .CI (n_316));
FA_X1 i_412 (.CO (n_305), .S (n_304), .A (n_288), .B (n_298), .CI (n_563));
NAND2_X1 slo__sro_c1045 (.ZN (slo__sro_n719), .A1 (n_216), .A2 (n_214));
INV_X1 slo__sro_c1367 (.ZN (slo__sro_n944), .A (n_295));
NAND2_X1 slo__sro_c1397 (.ZN (slo__sro_n961), .A1 (n_1068), .A2 (n_1031));
FA_X1 i_408 (.CO (n_357), .S (n_356), .A (n_350), .B (n_348), .CI (n_327));
INV_X1 slo__sro_c2132 (.ZN (slo__sro_n1481), .A (n_970));
FA_X1 i_406 (.CO (n_309), .S (n_308), .A (n_302), .B (n_304), .CI (n_571));
FA_X1 i_405 (.CO (n_331), .S (n_330), .A (n_303), .B (n_301), .CI (n_324));
FA_X1 i_404 (.CO (n_307), .S (n_306), .A (n_569), .B (n_300), .CI (n_573));
FA_X1 i_403 (.CO (n_359), .S (n_358), .A (n_329), .B (n_354), .CI (n_352));
FA_X1 i_402 (.CO (n_353), .S (n_352), .A (n_346), .B (n_344), .CI (n_342));
FA_X1 i_401 (.CO (n_355), .S (n_354), .A (n_340), .B (n_338), .CI (n_325));
NAND2_X1 slo__sro_c1339 (.ZN (slo__sro_n919), .A1 (n_384), .A2 (n_359));
NOR2_X1 i_399 (.ZN (n_661), .A1 (slo__sro_n692), .A2 (n_555));
NOR2_X1 i_398 (.ZN (n_659), .A1 (n_240), .A2 (n_219));
INV_X1 i_397 (.ZN (n_657), .A (n_659));
NOR2_X1 i_396 (.ZN (n_655), .A1 (slo__sro_n716), .A2 (n_503));
INV_X1 i_395 (.ZN (n_653), .A (n_655));
NAND2_X1 i_394 (.ZN (n_651), .A1 (n_503), .A2 (slo__sro_n716));
AND2_X1 i_393 (.ZN (n_649), .A1 (n_240), .A2 (n_219));
AND2_X1 i_392 (.ZN (n_647), .A1 (n_511), .A2 (n_651));
NAND3_X2 sgo__c341 (.ZN (sgo__n185), .A1 (n_1397), .A2 (opt_ipo_n1940), .A3 (n_513));
AOI21_X1 i_390 (.ZN (n_643), .A (n_649), .B1 (slo__sro_n692), .B2 (n_555));
OAI22_X2 i_389 (.ZN (n_641), .A1 (opt_ipo_n1967), .A2 (n_647), .B1 (n_661), .B2 (n_643));
NOR2_X1 i_387 (.ZN (n_636), .A1 (n_501), .A2 (n_457));
INV_X1 slo__sro_c2695 (.ZN (slo__sro_n1859), .A (n_761));
NOR3_X1 slo__c829 (.ZN (slo__n521), .A1 (sgo__sro_n14), .A2 (opt_ipo_n2168), .A3 (n_1104));
NAND2_X1 i_384 (.ZN (n_614), .A1 (n_553), .A2 (n_590));
OAI21_X1 i_383 (.ZN (n_594), .A (opt_ipo_n2116), .B1 (n_553), .B2 (n_590));
XNOR2_X1 i_382 (.ZN (\aggregated_res[14] [26] ), .A (n_616), .B (n_594));
HA_X1 i_381 (.CO (n_592), .S (n_590), .A (n_282), .B (n_284));
FA_X1 i_380 (.CO (n_588), .S (n_284), .A (slo__sro_n1800), .B (n_280), .CI (n_261));
FA_X1 i_379 (.CO (n_573), .S (n_280), .A (slo__sro_n752), .B (n_274), .CI (n_255));
FA_X1 i_378 (.CO (n_572), .S (n_274), .A (n_247), .B (n_245), .CI (n_243));
FA_X1 i_377 (.CO (n_245), .S (n_244), .A (p_3[25]), .B (p_4[25]), .CI (p_5[25]));
FA_X1 i_376 (.CO (n_247), .S (n_246), .A (p_6[25]), .B (p_7[25]), .CI (p_8[25]));
FA_X1 i_375 (.CO (n_571), .S (n_282), .A (n_257), .B (n_278), .CI (n_276));
FA_X1 i_374 (.CO (n_569), .S (n_276), .A (n_251), .B (n_272), .CI (n_270));
FA_X1 i_373 (.CO (n_567), .S (n_270), .A (p_9[26]), .B (p_10[26]), .CI (p_11[26]));
FA_X1 i_372 (.CO (n_565), .S (n_272), .A (p_12[26]), .B (p_15[26]), .CI (n_249));
FA_X1 i_371 (.CO (n_249), .S (n_248), .A (p_9[25]), .B (p_10[25]), .CI (p_11[25]));
FA_X1 i_370 (.CO (n_225), .S (n_224), .A (p_6[24]), .B (p_7[24]), .CI (p_8[24]));
FA_X1 i_369 (.CO (n_227), .S (n_226), .A (p_9[24]), .B (p_10[24]), .CI (p_11[24]));
FA_X1 i_368 (.CO (n_563), .S (n_278), .A (n_268), .B (n_266), .CI (n_264));
FA_X1 i_367 (.CO (n_561), .S (n_264), .A (p_0[26]), .B (p_1[26]), .CI (p_2[26]));
FA_X1 i_366 (.CO (n_559), .S (n_266), .A (p_3[26]), .B (p_4[26]), .CI (p_5[26]));
FA_X1 i_365 (.CO (n_557), .S (n_268), .A (p_6[26]), .B (p_7[26]), .CI (p_8[26]));
AND2_X2 CLOCK_sgo__sro_c3464 (.ZN (n_896), .A1 (n_470), .A2 (n_832));
NAND2_X1 slo__sro_c1135 (.ZN (slo__sro_n793), .A1 (n_170), .A2 (n_162));
FA_X1 i_362 (.CO (n_205), .S (n_204), .A (p_6[23]), .B (p_7[23]), .CI (p_8[23]));
FA_X1 i_361 (.CO (n_207), .S (n_206), .A (p_9[23]), .B (p_10[23]), .CI (p_15[23]));
FA_X1 i_360 (.CO (n_221), .S (n_220), .A (p_0[24]), .B (p_1[24]), .CI (p_2[24]));
FA_X1 i_359 (.CO (n_223), .S (n_222), .A (p_3[24]), .B (p_4[24]), .CI (p_5[24]));
INV_X1 slo__sro_c2665 (.ZN (slo__sro_n1835), .A (n_220));
FA_X1 i_357 (.CO (n_201), .S (n_200), .A (p_0[23]), .B (p_1[23]), .CI (p_2[23]));
FA_X1 i_356 (.CO (n_203), .S (n_202), .A (p_3[23]), .B (p_4[23]), .CI (p_5[23]));
FA_X1 i_355 (.CO (n_243), .S (n_242), .A (p_0[25]), .B (p_1[25]), .CI (p_2[25]));
INV_X1 slo__sro_c1057 (.ZN (slo__sro_n730), .A (slo__sro_n791));
FA_X1 i_353 (.CO (n_215), .S (n_214), .A (n_208), .B (n_471), .CI (n_465));
FA_X1 i_352 (.CO (n_209), .S (n_208), .A (n_467), .B (n_469), .CI (n_461));
INV_X2 sgo__sro_c582 (.ZN (sgo__sro_n311), .A (n_665));
FA_X1 i_350 (.CO (n_217), .S (n_216), .A (n_210), .B (n_212), .CI (n_473));
FA_X1 i_349 (.CO (n_213), .S (n_212), .A (n_204), .B (n_202), .CI (n_200));
NAND2_X1 slo__sro_c2558 (.ZN (slo__sro_n1749), .A1 (n_308), .A2 (n_306));
INV_X1 slo__sro_c1031 (.ZN (slo__sro_n708), .A (n_335));
FA_X1 i_346 (.CO (n_261), .S (n_260), .A (n_254), .B (n_256), .CI (n_237));
FA_X1 i_345 (.CO (n_257), .S (n_256), .A (n_242), .B (slo__sro_n1818), .CI (slo__sro_n750));
FA_X1 i_344 (.CO (n_255), .S (n_254), .A (n_248), .B (n_246), .CI (n_244));
NAND2_X1 slo__sro_c1119 (.ZN (slo__sro_n780), .A1 (n_207), .A2 (p_15[24]));
INV_X1 slo__sro_c1089 (.ZN (slo__sro_n755), .A (slo__sro_n777));
INV_X1 slo__sro_c2651 (.ZN (slo__sro_n1821), .A (n_209));
BUF_X1 slo__c2689 (.Z (sgo__n228), .A (slo__n1848));
FA_X1 i_339 (.CO (n_233), .S (n_232), .A (n_226), .B (n_224), .CI (n_222));
FA_X1 i_338 (.CO (n_251), .S (n_250), .A (p_15[25]), .B (n_227), .CI (n_225));
INV_X1 i_337 (.ZN (n_549), .A (n_459));
INV_X1 i_336 (.ZN (n_547), .A (n_407));
INV_X2 sgo__sro_c9 (.ZN (sgo__sro_n8), .A (sgo__sro_n9));
NOR2_X4 i_334 (.ZN (n_543), .A1 (n_455), .A2 (n_447));
INV_X4 i_333 (.ZN (n_541), .A (n_543));
NAND2_X1 i_332 (.ZN (n_539), .A1 (n_429), .A2 (n_127));
NAND2_X1 i_331 (.ZN (n_537), .A1 (n_459), .A2 (n_407));
NOR2_X2 i_330 (.ZN (n_535), .A1 (n_429), .A2 (n_127));
INV_X4 i_329 (.ZN (n_533), .A (n_535));
NAND3_X4 i_328 (.ZN (n_531), .A1 (n_533), .A2 (n_453), .A3 (n_541));
AOI21_X4 i_327 (.ZN (n_529), .A (n_531), .B1 (n_539), .B2 (n_537));
INV_X1 CLOCK_slo__sro_c3951 (.ZN (CLOCK_slo__sro_n2897), .A (n_495));
INV_X1 slo__sro_c914 (.ZN (slo__sro_n604), .A (n_1218));
NAND2_X2 i_323 (.ZN (n_521), .A1 (n_421), .A2 (n_419));
BUF_X1 CLOCK_sgo__c3557 (.Z (n_459), .A (CLOCK_sgo__n2634));
AOI21_X2 i_321 (.ZN (n_517), .A (n_519), .B1 (n_549), .B2 (n_547));
INV_X1 i_320 (.ZN (n_515), .A (n_517));
AOI22_X4 i_319 (.ZN (n_513), .A1 (CLOCK_spw__n3015), .A2 (n_447), .B1 (n_541), .B2 (n_1137));
NAND2_X2 i_318 (.ZN (n_511), .A1 (n_457), .A2 (n_501));
NOR2_X1 slo__c868 (.ZN (slo__n557), .A1 (n_1092), .A2 (sgo__sro_n16));
INV_X2 i_316 (.ZN (n_507), .A (n_509));
OAI21_X1 i_315 (.ZN (n_505), .A (n_511), .B1 (n_457), .B2 (n_501));
XNOR2_X1 i_314 (.ZN (\aggregated_res[14] [22] ), .A (n_509), .B (n_505));
HA_X1 i_313 (.CO (n_503), .S (spw__n3514), .A (n_177), .B (n_196));
FA_X1 i_312 (.CO (n_498), .S (n_196), .A (n_192), .B (n_190), .CI (slo__sro_n726));
INV_X1 slo__sro_c1075 (.ZN (slo__sro_n745), .A (n_215));
FA_X1 i_310 (.CO (n_472), .S (n_188), .A (n_167), .B (n_165), .CI (n_163));
FA_X1 i_309 (.CO (n_471), .S (n_190), .A (n_169), .B (n_186), .CI (n_184));
FA_X1 i_308 (.CO (n_469), .S (n_184), .A (p_6[22]), .B (p_7[22]), .CI (p_8[22]));
FA_X1 i_307 (.CO (n_467), .S (n_186), .A (p_9[22]), .B (p_10[22]), .CI (p_15[22]));
FA_X1 i_306 (.CO (n_465), .S (n_192), .A (n_182), .B (n_180), .CI (n_171));
FA_X1 i_305 (.CO (n_463), .S (n_180), .A (p_0[22]), .B (p_1[22]), .CI (p_2[22]));
FA_X1 i_304 (.CO (n_461), .S (n_182), .A (p_3[22]), .B (p_4[22]), .CI (p_5[22]));
HA_X1 i_303 (.CO (n_127), .S (CLOCK_sgo__n2634), .A (n_427), .B (n_425));
INV_X1 slo__sro_c1871 (.ZN (slo__sro_n1292), .A (n_135));
INV_X1 slo__sro_c1928 (.ZN (slo__sro_n1334), .A (n_699));
FA_X1 i_300 (.CO (n_173), .S (n_172), .A (n_168), .B (n_166), .CI (n_164));
FA_X1 i_299 (.CO (n_165), .S (n_164), .A (p_3[21]), .B (p_4[21]), .CI (p_5[21]));
FA_X1 i_298 (.CO (n_167), .S (n_166), .A (p_6[21]), .B (p_7[21]), .CI (p_8[21]));
FA_X1 i_297 (.CO (n_169), .S (n_168), .A (p_9[21]), .B (p_15[21]), .CI (n_439));
NAND2_X1 slo__sro_c1149 (.ZN (slo__sro_n804), .A1 (n_1146), .A2 (n_1144));
FA_X1 i_295 (.CO (n_171), .S (n_170), .A (n_441), .B (n_431), .CI (n_437));
FA_X1 i_294 (.CO (n_163), .S (n_162), .A (p_0[21]), .B (p_1[21]), .CI (p_2[21]));
OR2_X4 i_293 (.ZN (n_453), .A1 (n_143), .A2 (n_160));
NAND2_X1 i_292 (.ZN (n_451), .A1 (n_143), .A2 (n_160));
NAND2_X1 i_291 (.ZN (n_449), .A1 (n_453), .A2 (n_451));
HA_X1 i_290 (.CO (n_447), .S (n_160), .A (n_156), .B (slo__sro_n1756));
INV_X1 slo__sro_c2601 (.ZN (slo__sro_n1781), .A (n_119));
FA_X1 i_288 (.CO (n_443), .S (n_154), .A (n_150), .B (n_148), .CI (n_146));
FA_X1 i_287 (.CO (n_441), .S (n_146), .A (p_3[20]), .B (p_4[20]), .CI (p_5[20]));
FA_X1 i_286 (.CO (n_439), .S (n_148), .A (p_6[20]), .B (p_7[20]), .CI (p_8[20]));
FA_X1 i_285 (.CO (n_437), .S (n_150), .A (p_9[20]), .B (p_15[20]), .CI (n_133));
FA_X1 i_284 (.CO (n_435), .S (n_156), .A (n_144), .B (n_152), .CI (n_137));
INV_X1 slo__sro_c1885 (.ZN (slo__sro_n1300), .A (n_435));
FA_X1 i_282 (.CO (n_431), .S (n_144), .A (p_0[20]), .B (p_1[20]), .CI (p_2[20]));
FA_X1 i_281 (.CO (n_143), .S (n_429), .A (n_138), .B (n_125), .CI (n_140));
FA_X1 i_280 (.CO (n_141), .S (n_140), .A (n_121), .B (n_136), .CI (n_123));
FA_X1 i_279 (.CO (n_123), .S (n_427), .A (n_114), .B (n_112), .CI (n_118));
INV_X1 slo__sro_c2633 (.ZN (slo__sro_n1805), .A (n_250));
FA_X1 i_277 (.CO (n_133), .S (n_132), .A (p_6[19]), .B (p_7[19]), .CI (p_8[19]));
FA_X1 i_276 (.CO (n_119), .S (n_118), .A (p_15[18]), .B (n_393), .CI (n_395));
FA_X1 i_275 (.CO (n_113), .S (n_112), .A (p_0[18]), .B (p_1[18]), .CI (p_2[18]));
FA_X1 i_274 (.CO (n_125), .S (n_425), .A (n_399), .B (n_120), .CI (n_403));
FA_X1 i_273 (.CO (n_121), .S (n_120), .A (n_397), .B (n_401), .CI (n_116));
FA_X1 i_272 (.CO (n_139), .S (n_138), .A (n_130), .B (n_128), .CI (n_134));
FA_X1 i_271 (.CO (n_135), .S (n_134), .A (p_15[19]), .B (n_117), .CI (n_115));
FA_X1 i_270 (.CO (n_115), .S (n_114), .A (p_3[18]), .B (p_4[18]), .CI (p_5[18]));
FA_X1 i_269 (.CO (n_117), .S (n_116), .A (p_6[18]), .B (p_7[18]), .CI (p_8[18]));
FA_X1 i_268 (.CO (n_129), .S (n_128), .A (p_0[19]), .B (p_1[19]), .CI (p_2[19]));
FA_X1 i_267 (.CO (n_131), .S (n_130), .A (p_3[19]), .B (p_4[19]), .CI (p_5[19]));
OAI21_X4 sgo__sro_c10 (.ZN (n_1116), .A (sgo__sro_n8), .B1 (opt_ipo_n2091), .B2 (n_1109));
NAND2_X2 i_265 (.ZN (n_421), .A1 (n_405), .A2 (n_411));
NAND2_X1 i_264 (.ZN (n_419), .A1 (n_409), .A2 (n_379));
INV_X1 i_263 (.ZN (n_418), .A (n_419));
AOI21_X1 i_262 (.ZN (n_417), .A (n_391), .B1 (opt_ipo_n1948), .B2 (n_390));
OAI21_X1 i_261 (.ZN (n_415), .A (n_421), .B1 (n_405), .B2 (n_411));
OAI22_X1 i_260 (.ZN (n_413), .A1 (n_409), .A2 (n_379), .B1 (n_418), .B2 (n_417));
XOR2_X1 i_259 (.Z (\aggregated_res[14] [17] ), .A (n_415), .B (n_413));
NAND2_X2 slo__mro_c672 (.ZN (n_1073), .A1 (sgo__sro_n149), .A2 (n_1392));
FA_X1 i_257 (.CO (n_407), .S (n_405), .A (n_106), .B (n_95), .CI (n_108));
FA_X1 i_256 (.CO (n_403), .S (n_108), .A (n_91), .B (n_104), .CI (n_93));
FA_X1 i_255 (.CO (n_93), .S (n_92), .A (n_88), .B (n_86), .CI (n_84));
FA_X1 i_254 (.CO (n_401), .S (n_104), .A (n_89), .B (n_87), .CI (n_85));
FA_X1 i_253 (.CO (n_85), .S (n_84), .A (p_0[16]), .B (p_1[16]), .CI (p_2[16]));
FA_X1 i_252 (.CO (n_87), .S (n_86), .A (p_3[16]), .B (p_4[16]), .CI (p_5[16]));
FA_X1 i_251 (.CO (n_89), .S (n_88), .A (p_6[16]), .B (p_7[16]), .CI (p_15[16]));
FA_X1 i_250 (.CO (n_95), .S (n_94), .A (n_90), .B (n_371), .CI (n_377));
FA_X1 i_249 (.CO (n_91), .S (n_90), .A (n_373), .B (n_375), .CI (n_369));
FA_X1 i_248 (.CO (n_399), .S (n_106), .A (n_102), .B (n_100), .CI (n_98));
FA_X1 i_247 (.CO (n_397), .S (n_98), .A (p_0[17]), .B (p_1[17]), .CI (p_2[17]));
FA_X1 i_246 (.CO (n_395), .S (n_100), .A (p_3[17]), .B (p_4[17]), .CI (p_5[17]));
FA_X1 i_245 (.CO (n_393), .S (n_102), .A (p_6[17]), .B (p_7[17]), .CI (p_15[17]));
NOR2_X2 i_244 (.ZN (n_391), .A1 (n_310), .A2 (n_82));
NAND2_X1 i_243 (.ZN (n_390), .A1 (n_310), .A2 (n_82));
NAND2_X2 i_242 (.ZN (n_389), .A1 (n_262), .A2 (n_241));
OAI21_X2 i_241 (.ZN (n_387), .A (n_389), .B1 (n_187), .B2 (n_197));
OAI21_X4 i_240 (.ZN (n_385), .A (n_367), .B1 (n_387), .B2 (n_365));
AOI21_X1 i_238 (.ZN (n_381), .A (n_391), .B1 (n_310), .B2 (n_82));
XNOR2_X1 i_237 (.ZN (\aggregated_res[14] [15] ), .A (opt_ipo_n1948), .B (n_381));
FA_X1 i_236 (.CO (n_379), .S (n_82), .A (n_78), .B (n_287), .CI (n_80));
FA_X1 i_235 (.CO (n_377), .S (n_80), .A (n_74), .B (n_72), .CI (n_283));
FA_X1 i_234 (.CO (n_375), .S (n_72), .A (p_0[15]), .B (p_1[15]), .CI (p_2[15]));
FA_X1 i_233 (.CO (n_373), .S (n_74), .A (p_3[15]), .B (p_4[15]), .CI (p_5[15]));
FA_X1 i_232 (.CO (n_371), .S (n_78), .A (n_286), .B (n_281), .CI (n_76));
FA_X1 i_231 (.CO (n_369), .S (n_76), .A (p_6[15]), .B (p_15[15]), .CI (n_285));
NAND2_X2 i_230 (.ZN (n_367), .A1 (n_198), .A2 (opt_ipo_n2150));
NOR2_X2 i_229 (.ZN (n_365), .A1 (n_198), .A2 (opt_ipo_n2150));
OAI21_X1 i_228 (.ZN (n_363), .A (n_367), .B1 (n_198), .B2 (opt_ipo_n2150));
HA_X1 i_227 (.CO (n_310), .S (n_70), .A (n_66), .B (n_68));
FA_X1 i_226 (.CO (n_287), .S (n_68), .A (n_62), .B (n_60), .CI (n_195));
FA_X1 i_225 (.CO (n_286), .S (n_60), .A (p_0[14]), .B (p_1[14]), .CI (p_2[14]));
FA_X1 i_224 (.CO (n_285), .S (n_62), .A (p_3[14]), .B (p_4[14]), .CI (p_5[14]));
FA_X1 i_223 (.CO (n_283), .S (n_66), .A (n_193), .B (n_189), .CI (n_64));
BUF_X4 slo__c2295 (.Z (\aggregated_res[14] [35] ), .A (slo__n1579));
INV_X1 i_221 (.ZN (n_279), .A (n_48));
INV_X1 i_220 (.ZN (n_277), .A (n_46));
NAND2_X1 i_219 (.ZN (n_275), .A1 (n_279), .A2 (n_277));
AOI21_X2 i_218 (.ZN (n_273), .A (n_155), .B1 (n_157), .B2 (n_153));
NOR2_X1 i_217 (.ZN (n_271), .A1 (n_185), .A2 (n_145));
AOI21_X1 i_216 (.ZN (n_269), .A (n_273), .B1 (n_185), .B2 (n_145));
NOR2_X2 i_215 (.ZN (n_267), .A1 (n_271), .A2 (n_269));
NOR2_X2 i_214 (.ZN (n_265), .A1 (n_279), .A2 (n_277));
INV_X1 i_213 (.ZN (n_263), .A (n_265));
OAI21_X2 i_212 (.ZN (n_262), .A (n_275), .B1 (n_267), .B2 (n_265));
NAND2_X1 i_211 (.ZN (n_241), .A1 (n_187), .A2 (n_197));
OAI21_X1 i_210 (.ZN (n_199), .A (n_241), .B1 (n_187), .B2 (n_197));
XOR2_X1 i_209 (.Z (\aggregated_res[14] [13] ), .A (n_262), .B (n_199));
FA_X1 i_208 (.CO (n_198), .S (n_197), .A (n_54), .B (n_47), .CI (n_56));
FA_X1 i_207 (.CO (n_195), .S (n_56), .A (n_45), .B (n_52), .CI (n_50));
FA_X1 i_206 (.CO (n_193), .S (n_50), .A (p_0[13]), .B (p_1[13]), .CI (p_2[13]));
FA_X1 i_205 (.CO (n_191), .S (n_52), .A (p_3[13]), .B (p_4[13]), .CI (p_5[13]));
FA_X1 i_204 (.CO (n_189), .S (n_54), .A (p_15[13]), .B (n_43), .CI (n_41));
FA_X1 i_203 (.CO (n_47), .S (n_46), .A (n_42), .B (n_40), .CI (n_44));
FA_X1 i_202 (.CO (n_45), .S (n_44), .A (p_15[12]), .B (n_35), .CI (n_33));
FA_X1 i_201 (.CO (n_41), .S (n_40), .A (p_0[12]), .B (p_1[12]), .CI (p_2[12]));
FA_X1 i_200 (.CO (n_43), .S (n_42), .A (p_3[12]), .B (p_4[12]), .CI (p_5[12]));
HA_X1 i_199 (.CO (n_187), .S (n_48), .A (n_37), .B (n_39));
NAND2_X1 slo__sro_c2318 (.ZN (slo__sro_n1595), .A1 (n_34), .A2 (n_147));
FA_X1 i_197 (.CO (n_33), .S (n_32), .A (p_0[11]), .B (p_1[11]), .CI (p_2[11]));
NAND2_X1 slo__sro_c2330 (.ZN (slo__sro_n1601), .A1 (p_0[10]), .A2 (p_1[10]));
FA_X1 i_195 (.CO (n_35), .S (n_34), .A (p_3[11]), .B (p_4[11]), .CI (p_15[11]));
INV_X1 i_194 (.ZN (n_183), .A (n_105));
INV_X1 i_193 (.ZN (n_181), .A (n_126));
OAI211_X1 i_192 (.ZN (n_179), .A (n_71), .B (n_103), .C1 (n_73), .C2 (n_101));
INV_X1 i_191 (.ZN (n_178), .A (n_179));
OAI21_X1 i_190 (.ZN (n_161), .A (n_183), .B1 (n_53), .B2 (n_57));
OAI211_X2 i_189 (.ZN (n_159), .A (n_63), .B (n_124), .C1 (n_178), .C2 (n_161));
NAND2_X2 i_188 (.ZN (n_157), .A1 (n_159), .A2 (n_181));
NOR2_X2 i_187 (.ZN (n_155), .A1 (opt_ipo_n2336), .A2 (n_28));
NAND2_X2 i_186 (.ZN (n_153), .A1 (opt_ipo_n2336), .A2 (n_28));
OAI21_X1 i_185 (.ZN (n_151), .A (n_153), .B1 (opt_ipo_n2336), .B2 (n_28));
XOR2_X1 i_184 (.Z (\aggregated_res[14] [10] ), .A (n_157), .B (n_151));
FA_X1 i_183 (.CO (n_149), .S (n_28), .A (n_109), .B (n_107), .CI (n_26));
FA_X1 i_182 (.CO (n_147), .S (n_26), .A (p_3[10]), .B (p_4[10]), .CI (p_15[10]));
HA_X1 i_181 (.CO (n_145), .S (n_30), .A (n_24), .B (slo__sro_n847));
NAND2_X1 slo__sro_c2342 (.ZN (slo__sro_n1607), .A1 (n_646), .A2 (n_648));
NOR2_X1 i_179 (.ZN (n_126), .A1 (n_55), .A2 (n_22));
NAND2_X1 i_178 (.ZN (n_124), .A1 (n_55), .A2 (n_22));
AOI21_X1 i_177 (.ZN (n_122), .A (n_126), .B1 (n_55), .B2 (n_22));
OAI22_X1 i_176 (.ZN (n_111), .A1 (n_57), .A2 (n_53), .B1 (n_61), .B2 (n_65));
XNOR2_X1 i_175 (.ZN (\aggregated_res[14] [9] ), .A (n_122), .B (n_111));
NAND2_X1 slo__sro_c1229 (.ZN (slo__sro_n856), .A1 (slo__sro_n814), .A2 (n_1084));
FA_X1 i_173 (.CO (n_109), .S (n_18), .A (p_0[9]), .B (p_1[9]), .CI (p_2[9]));
FA_X1 i_172 (.CO (n_107), .S (n_20), .A (p_3[9]), .B (p_15[9]), .CI (n_58));
NOR2_X2 i_171 (.ZN (n_105), .A1 (n_29), .A2 (n_31));
NAND2_X1 i_170 (.ZN (n_103), .A1 (n_29), .A2 (n_31));
NOR2_X1 i_169 (.ZN (n_101), .A1 (n_23), .A2 (n_27));
NAND2_X1 i_168 (.ZN (n_99), .A1 (n_38), .A2 (p_15[4]));
NAND2_X1 i_167 (.ZN (n_97), .A1 (p_0[2]), .A2 (p_15[2]));
NAND2_X1 i_166 (.ZN (n_96), .A1 (p_0[3]), .A2 (p_15[3]));
NOR2_X1 i_165 (.ZN (n_83), .A1 (p_0[3]), .A2 (p_15[3]));
AOI21_X1 i_164 (.ZN (n_81), .A (n_83), .B1 (n_97), .B2 (n_96));
OAI21_X1 i_163 (.ZN (n_79), .A (n_81), .B1 (n_38), .B2 (p_15[4]));
NAND2_X1 i_162 (.ZN (n_77), .A1 (n_99), .A2 (n_79));
AND2_X1 i_161 (.ZN (n_75), .A1 (n_25), .A2 (n_49));
OAI22_X1 i_160 (.ZN (n_73), .A1 (n_25), .A2 (n_49), .B1 (n_77), .B2 (n_75));
NAND2_X1 i_159 (.ZN (n_71), .A1 (n_23), .A2 (n_27));
AOI21_X1 i_158 (.ZN (n_69), .A (n_101), .B1 (n_73), .B2 (n_71));
INV_X1 i_157 (.ZN (n_67), .A (n_69));
AOI21_X1 i_156 (.ZN (n_65), .A (n_105), .B1 (n_103), .B2 (n_67));
NAND2_X1 i_155 (.ZN (n_63), .A1 (n_53), .A2 (n_57));
INV_X1 i_154 (.ZN (n_61), .A (n_63));
OAI21_X1 i_153 (.ZN (n_59), .A (n_63), .B1 (n_53), .B2 (n_57));
XNOR2_X1 i_152 (.ZN (\aggregated_res[14] [8] ), .A (n_65), .B (n_59));
FA_X1 i_151 (.CO (n_58), .S (n_57), .A (p_0[8]), .B (p_1[8]), .CI (p_2[8]));
HA_X1 i_150 (.CO (n_55), .S (n_53), .A (n_13), .B (slo__sro_n1181));
NAND2_X1 slo__sro_c1738 (.ZN (slo__sro_n1196), .A1 (n_440), .A2 (n_777));
HA_X1 i_148 (.CO (n_49), .S (n_38), .A (p_0[4]), .B (p_1[4]));
FA_X1 i_147 (.CO (n_14), .S (n_31), .A (p_0[7]), .B (p_1[7]), .CI (p_2[7]));
FA_X1 i_146 (.CO (n_13), .S (n_29), .A (p_15[7]), .B (n_10), .CI (n_12));
HA_X1 i_145 (.CO (n_12), .S (n_27), .A (p_15[6]), .B (n_11));
FA_X1 i_144 (.CO (n_11), .S (n_25), .A (p_0[5]), .B (p_1[5]), .CI (p_15[5]));
FA_X1 i_143 (.CO (n_10), .S (n_23), .A (p_0[6]), .B (p_1[6]), .CI (p_2[6]));
NAND2_X1 i_142 (.ZN (n_9), .A1 (n_1283), .A2 (p_14[62]));
NOR2_X2 i_141 (.ZN (n_8), .A1 (n_1238), .A2 (n_1274));
NAND2_X1 slo__sro_c775 (.ZN (slo__sro_n468), .A1 (n_546), .A2 (n_544));
OAI221_X2 i_139 (.ZN (n_6), .A (n_1145), .B1 (n_1287), .B2 (n_1306), .C1 (n_1238), .C2 (n_1235));
OR2_X1 i_138 (.ZN (n_5), .A1 (n_1384), .A2 (n_1293));
NOR2_X2 sgo__c163 (.ZN (sgo__n97), .A1 (n_444), .A2 (n_795));
INV_X1 i_136 (.ZN (n_3), .A (n_1376));
NAND2_X1 i_135 (.ZN (n_2), .A1 (n_1348), .A2 (n_3));
AOI21_X4 i_134 (.ZN (n_1), .A (n_2), .B1 (sgo__sro_n32), .B2 (n_1386));
OAI21_X4 i_133 (.ZN (\aggregated_res[14] [63] ), .A (n_9), .B1 (n_1), .B2 (n_1373));
NAND2_X4 i_132 (.ZN (n_0), .A1 (sgo__sro_n32), .A2 (n_1386));
XNOR2_X1 i_131 (.ZN (n_1398), .A (n_0), .B (n_1346));
INV_X1 i_130 (.ZN (\aggregated_res[14] [58] ), .A (n_1398));
XNOR2_X2 i_129 (.ZN (\aggregated_res[14] [44] ), .A (n_1174), .B (n_1067));
NAND2_X1 i_128 (.ZN (n_1367), .A1 (n_1033), .A2 (n_1070));
NOR3_X4 sgo__sro_c22 (.ZN (n_1254), .A1 (sgo__sro_n14), .A2 (opt_ipo_n2168), .A3 (n_1104));
NOR2_X1 i_126 (.ZN (n_1365), .A1 (n_1078), .A2 (n_1018));
NAND2_X1 i_125 (.ZN (n_1072), .A1 (n_1078), .A2 (n_1018));
INV_X1 slo__sro_c659 (.ZN (slo__sro_n366), .A (n_92));
NAND2_X2 i_123 (.ZN (n_1362), .A1 (slo__sro_n332), .A2 (n_1095));
AOI21_X2 i_122 (.ZN (n_1361), .A (n_1077), .B1 (n_1362), .B2 (n_1367));
XNOR2_X2 i_121 (.ZN (\aggregated_res[14] [41] ), .A (n_1361), .B (n_1056));
NAND2_X1 i_120 (.ZN (n_1342), .A1 (n_767), .A2 (n_729));
INV_X1 i_119 (.ZN (n_1131), .A (n_727));
NOR2_X1 i_118 (.ZN (n_1160), .A1 (n_665), .A2 (n_592));
OAI21_X1 i_117 (.ZN (n_1341), .A (n_616), .B1 (n_553), .B2 (n_590));
NAND2_X2 i_116 (.ZN (n_961), .A1 (n_1341), .A2 (opt_ipo_n2116));
INV_X1 i_115 (.ZN (n_1340), .A (n_961));
AOI21_X4 i_114 (.ZN (n_959), .A (n_1160), .B1 (n_1340), .B2 (opt_ipo_n2153));
INV_X2 CLOCK_slo__c3941 (.ZN (n_767), .A (CLOCK_slo__n2890));
INV_X1 CLOCK_slo__xsl_c3907 (.ZN (CLOCK_slo__xsl_n2867), .A (n_525));
NOR2_X4 i_111 (.ZN (n_1047), .A1 (n_7), .A2 (n_6));
INV_X1 i_110 (.ZN (n_1331), .A (n_1));
INV_X1 i_109 (.ZN (n_1241), .A (n_1269));
NAND2_X1 i_108 (.ZN (n_1145), .A1 (n_1281), .A2 (n_1292));
XNOR2_X1 i_107 (.ZN (n_1130), .A (n_1283), .B (p_14[62]));
AOI21_X2 i_106 (.ZN (n_1127), .A (n_1130), .B1 (n_1331), .B2 (n_1374));
INV_X1 CLOCK_sgo__sro_c3685 (.ZN (CLOCK_sgo__sro_n2705), .A (n_663));
NOR2_X4 slo__c965 (.ZN (slo__n651), .A1 (n_1257), .A2 (n_1255));
NOR2_X4 i_103 (.ZN (\aggregated_res[14] [62] ), .A1 (n_1126), .A2 (n_1127));
NAND2_X1 i_102 (.ZN (n_1124), .A1 (n_1378), .A2 (n_1379));
INV_X1 i_101 (.ZN (n_1120), .A (n_1124));
OR2_X1 i_100 (.ZN (n_1118), .A1 (n_1377), .A2 (n_1355));
NAND2_X4 i_99 (.ZN (n_1117), .A1 (n_0), .A2 (n_1348));
NAND3_X2 i_98 (.ZN (n_1114), .A1 (n_1117), .A2 (n_1347), .A3 (n_1368));
NAND2_X1 i_97 (.ZN (n_1113), .A1 (n_1114), .A2 (n_1118));
NAND2_X1 i_96 (.ZN (n_1111), .A1 (n_1113), .A2 (n_1120));
NAND3_X1 i_95 (.ZN (n_1110), .A1 (n_1114), .A2 (n_1124), .A3 (n_1118));
NAND2_X2 i_94 (.ZN (\aggregated_res[14] [61] ), .A1 (n_1111), .A2 (n_1110));
NAND3_X2 i_93 (.ZN (n_1107), .A1 (n_1117), .A2 (n_1371), .A3 (n_1347));
OR2_X1 i_92 (.ZN (n_1101), .A1 (n_1344), .A2 (n_1350));
NAND3_X2 i_91 (.ZN (n_1100), .A1 (n_1107), .A2 (n_1352), .A3 (n_1101));
NAND2_X1 i_90 (.ZN (n_1099), .A1 (n_1107), .A2 (n_1101));
NAND2_X2 i_89 (.ZN (n_1098), .A1 (n_1099), .A2 (n_1353));
NAND2_X4 i_88 (.ZN (\aggregated_res[14] [60] ), .A1 (n_1098), .A2 (n_1100));
INV_X1 i_87 (.ZN (n_1091), .A (n_1396));
NOR2_X1 i_86 (.ZN (n_1090), .A1 (n_1384), .A2 (n_1293));
NAND2_X1 i_85 (.ZN (n_1250), .A1 (n_1384), .A2 (n_1293));
NOR3_X4 sgo__c305 (.ZN (sgo__n168), .A1 (slo__n419), .A2 (n_659), .A3 (n_655));
AOI21_X4 i_83 (.ZN (n_1081), .A (n_1091), .B1 (sgo__sro_n149), .B2 (n_1392));
NOR2_X1 i_82 (.ZN (n_1080), .A1 (n_1081), .A2 (n_1391));
NAND2_X2 i_81 (.ZN (n_1076), .A1 (n_1080), .A2 (n_1327));
OAI21_X2 i_80 (.ZN (n_1074), .A (n_1328), .B1 (n_1081), .B2 (n_1391));
NAND2_X4 i_79 (.ZN (\aggregated_res[14] [57] ), .A1 (n_1076), .A2 (n_1074));
AOI21_X2 slo__c733 (.ZN (slo__n416), .A (n_1156), .B1 (n_1129), .B2 (n_1133));
NOR2_X1 i_77 (.ZN (n_1071), .A1 (n_1391), .A2 (n_1091));
INV_X1 slo__xsl_c705 (.ZN (slo__xsl_n395), .A (n_738));
NAND2_X1 i_75 (.ZN (n_1067), .A1 (n_1169), .A2 (n_1173));
NAND2_X1 i_74 (.ZN (n_1059), .A1 (n_1075), .A2 (n_1367));
INV_X1 CLOCK_slo__mro_c3867 (.ZN (CLOCK_slo__mro_n2829), .A (n_1342));
INV_X1 i_685 (.ZN (n_21), .A (p_1[36]));
INV_X1 i_674 (.ZN (n_19), .A (p_5[42]));
INV_X1 i_72 (.ZN (n_1044), .A (p_4[42]));
AOI21_X1 i_71 (.ZN (n_17), .A (p_6[42]), .B1 (p_5[42]), .B2 (n_1044));
OAI21_X1 i_70 (.ZN (n_991), .A (n_1072), .B1 (n_1123), .B2 (n_1365));
OAI21_X1 i_69 (.ZN (n_1029), .A (n_1250), .B1 (n_1047), .B2 (n_1090));
NAND2_X1 i_68 (.ZN (n_1040), .A1 (n_1117), .A2 (n_1347));
INV_X1 i_67 (.ZN (n_1039), .A (n_1040));
XOR2_X1 i_66 (.Z (\aggregated_res[14] [14] ), .A (n_387), .B (n_363));
NAND2_X1 i_65 (.ZN (n_994), .A1 (n_275), .A2 (n_263));
XNOR2_X1 i_64 (.ZN (\aggregated_res[14] [12] ), .A (n_267), .B (n_994));
AOI21_X2 i_63 (.ZN (n_931), .A (n_517), .B1 (n_407), .B2 (n_459));
AOI21_X2 i_62 (.ZN (n_943), .A (CLOCK_slo__xsl_n2800), .B1 (n_931), .B2 (n_539));
XNOR2_X1 i_61 (.ZN (\aggregated_res[14] [20] ), .A (n_449), .B (n_943));
NAND2_X1 i_60 (.ZN (n_930), .A1 (n_533), .A2 (n_539));
XOR2_X1 i_59 (.Z (\aggregated_res[14] [19] ), .A (n_931), .B (n_930));
NAND2_X1 i_58 (.ZN (n_927), .A1 (n_1400), .A2 (n_537));
XOR2_X1 i_57 (.Z (\aggregated_res[14] [18] ), .A (n_519), .B (n_927));
INV_X1 i_56 (.ZN (n_1137), .A (n_451));
INV_X1 i_55 (.ZN (n_1315), .A (p_6[44]));
INV_X1 i_54 (.ZN (n_1283), .A (p_14[61]));
OAI211_X1 i_53 (.ZN (n_1238), .A (n_1309), .B (n_1241), .C1 (n_1281), .C2 (n_1292));
AOI21_X1 i_52 (.ZN (n_1235), .A (n_1267), .B1 (n_1207), .B2 (n_1237));
INV_X1 i_51 (.ZN (n_1121), .A (n_651));
NAND2_X1 slo__sro_c1724 (.ZN (slo__sro_n1185), .A1 (p_15[8]), .A2 (p_3[8]));
OAI21_X1 i_49 (.ZN (n_1030), .A (n_1250), .B1 (n_1293), .B2 (n_1384));
NOR2_X1 i_48 (.ZN (n_1026), .A1 (n_1393), .A2 (n_1394));
CLKBUF_X1 slo___L1_c819 (.Z (slo___n509), .A (n_1245));
XOR2_X1 i_46 (.Z (\aggregated_res[14] [54] ), .A (n_1047), .B (n_1030));
INV_X2 i_45 (.ZN (n_1007), .A (n_1217));
NOR2_X1 i_44 (.ZN (n_1003), .A1 (n_1216), .A2 (n_1221));
INV_X2 sgo__sro_c254 (.ZN (sgo__sro_n137), .A (sgo__sro_n138));
XNOR2_X2 i_42 (.ZN (\aggregated_res[14] [48] ), .A (n_1002), .B (n_1003));
AND3_X2 slo__c935 (.ZN (n_1126), .A1 (n_1331), .A2 (n_1374), .A3 (n_1130));
OAI21_X1 i_40 (.ZN (n_992), .A (n_1072), .B1 (n_1018), .B2 (n_1078));
NOR2_X1 i_39 (.ZN (n_988), .A1 (n_1094), .A2 (n_1097));
XOR2_X1 i_38 (.Z (\aggregated_res[14] [39] ), .A (n_991), .B (n_988));
XOR2_X1 i_37 (.Z (\aggregated_res[14] [38] ), .A (n_1123), .B (n_992));
OAI21_X1 i_36 (.ZN (n_984), .A (n_1000), .B1 (n_896), .B2 (n_938));
XOR2_X1 i_35 (.Z (slo__n1579), .A (n_981), .B (n_944));
XOR2_X1 i_34 (.Z (\aggregated_res[14] [34] ), .A (n_983), .B (n_984));
NOR2_X1 i_33 (.ZN (n_958), .A1 (n_1160), .A2 (opt_ipo_n2152));
NOR2_X1 i_32 (.ZN (n_956), .A1 (n_752), .A2 (n_1131));
XOR2_X2 i_31 (.Z (\aggregated_res[14] [28] ), .A (n_959), .B (n_956));
XOR2_X1 i_30 (.Z (\aggregated_res[14] [27] ), .A (n_961), .B (n_958));
AOI21_X1 i_29 (.ZN (n_955), .A (n_661), .B1 (n_555), .B2 (slo__sro_n692));
AOI21_X1 i_28 (.ZN (n_953), .A (n_636), .B1 (n_507), .B2 (n_511));
OAI21_X2 i_27 (.ZN (n_952), .A (n_653), .B1 (slo__n539), .B2 (n_1121));
INV_X2 i_26 (.ZN (n_951), .A (n_952));
NOR2_X1 i_25 (.ZN (n_950), .A1 (n_655), .A2 (n_1121));
AOI21_X2 slo__c846 (.ZN (slo__n539), .A (n_636), .B1 (n_507), .B2 (n_511));
XNOR2_X2 i_23 (.ZN (\aggregated_res[14] [25] ), .A (n_955), .B (slo__sro_n535));
NOR2_X1 i_22 (.ZN (n_948), .A1 (n_659), .A2 (n_649));
XOR2_X2 i_21 (.Z (\aggregated_res[14] [24] ), .A (n_951), .B (n_948));
XOR2_X2 i_20 (.Z (\aggregated_res[14] [23] ), .A (n_953), .B (n_950));
AOI21_X1 i_19 (.ZN (n_947), .A (n_543), .B1 (n_447), .B2 (n_455));
OAI21_X2 i_18 (.ZN (n_941), .A (n_453), .B1 (n_943), .B2 (n_1137));
XNOR2_X2 i_17 (.ZN (\aggregated_res[14] [21] ), .A (n_947), .B (n_941));
NOR2_X1 i_16 (.ZN (n_932), .A1 (CLOCK_slo__xsl_n2867), .A2 (n_418));
XOR2_X1 i_15 (.Z (\aggregated_res[14] [16] ), .A (n_417), .B (n_932));
AOI21_X1 i_14 (.ZN (n_926), .A (n_271), .B1 (n_145), .B2 (n_185));
XOR2_X1 i_13 (.Z (\aggregated_res[14] [11] ), .A (n_273), .B (n_926));
OAI21_X1 i_12 (.ZN (n_922), .A (n_71), .B1 (n_23), .B2 (n_27));
AOI21_X1 i_11 (.ZN (n_918), .A (n_105), .B1 (n_31), .B2 (n_29));
XOR2_X1 i_10 (.Z (\aggregated_res[14] [7] ), .A (n_69), .B (n_918));
XOR2_X1 i_9 (.Z (\aggregated_res[14] [6] ), .A (n_73), .B (n_922));
XOR2_X1 i_8 (.Z (n_915), .A (n_49), .B (n_25));
XOR2_X1 i_7 (.Z (\aggregated_res[14] [5] ), .A (n_77), .B (n_915));
OAI21_X1 i_6 (.ZN (n_914), .A (n_99), .B1 (p_15[4]), .B2 (n_38));
XNOR2_X1 i_5 (.ZN (\aggregated_res[14] [4] ), .A (n_81), .B (n_914));
OAI21_X1 i_4 (.ZN (n_913), .A (n_96), .B1 (p_0[3]), .B2 (p_15[3]));
XOR2_X1 i_3 (.Z (\aggregated_res[14] [3] ), .A (n_97), .B (n_913));
OAI21_X1 i_2 (.ZN (n_912), .A (n_97), .B1 (p_0[2]), .B2 (p_15[2]));
INV_X1 i_1 (.ZN (\aggregated_res[14] [2] ), .A (n_912));
OAI222_X2 i_0 (.ZN (n_16), .A1 (p_5[44]), .A2 (n_1175), .B1 (n_1315), .B2 (p_5[44])
    , .C1 (n_1315), .C2 (n_1175));
INV_X1 sgo__sro_c27 (.ZN (sgo__sro_n18), .A (n_1089));
NAND2_X1 sgo__sro_c28 (.ZN (sgo__sro_n17), .A1 (n_690), .A2 (n_1089));
INV_X1 sgo__sro_c29 (.ZN (n_1147), .A (sgo__sro_n17));
XNOR2_X1 sgo__sro_c30 (.ZN (sgo__sro_n16), .A (n_690), .B (sgo__sro_n18));
INV_X1 sgo__sro_c141 (.ZN (sgo__sro_n87), .A (n_791));
AND2_X2 sgo__sro_c142 (.ZN (n_833), .A1 (slo__sro_n1193), .A2 (n_791));
XNOR2_X2 sgo__sro_c143 (.ZN (n_444), .A (slo__sro_n1193), .B (sgo__sro_n87));
OAI21_X4 sgo__sro_c173 (.ZN (n_1217), .A (sgo__sro_n101), .B1 (n_1189), .B2 (n_1225));
OR2_X1 sgo__sro_c179 (.ZN (sgo__sro_n105), .A1 (n_1184), .A2 (n_1208));
OAI21_X2 sgo__sro_c180 (.ZN (n_1002), .A (sgo__sro_n105), .B1 (n_1007), .B2 (n_1219));
NAND2_X1 sgo__sro_c54 (.ZN (sgo__sro_n34), .A1 (n_1389), .A2 (n_5));
INV_X1 sgo__sro_c55 (.ZN (sgo__sro_n33), .A (sgo__sro_n34));
OAI21_X4 sgo__sro_c56 (.ZN (sgo__sro_n32), .A (sgo__sro_n33), .B1 (slo__n432), .B2 (n_6));
INV_X2 sgo__c165 (.ZN (n_844), .A (sgo__n97));
AND2_X1 sgo__sro_c348 (.ZN (n_1018), .A1 (slo__sro_n1474), .A2 (n_974));
NOR2_X4 sgo__c203 (.ZN (sgo__n115), .A1 (n_1195), .A2 (n_1132));
NAND3_X4 sgo__c299 (.ZN (sgo__n166), .A1 (n_738), .A2 (n_995), .A3 (n_735));
XNOR2_X2 CLOCK_sgo__sro_c3576 (.ZN (n_1069), .A (slo__sro_n1339), .B (CLOCK_sgo__sro_n2645));
NAND2_X1 sgo__sro_c275 (.ZN (sgo__sro_n151), .A1 (n_1250), .A2 (n_1395));
INV_X1 sgo__sro_c276 (.ZN (sgo__sro_n150), .A (sgo__sro_n151));
OAI21_X4 sgo__sro_c277 (.ZN (sgo__sro_n149), .A (sgo__sro_n150), .B1 (n_1047), .B2 (n_1090));
INV_X4 sgo__c343 (.ZN (n_996), .A (sgo__n185));
INV_X1 CLOCK_slo__xsl_c3841 (.ZN (CLOCK_slo__xsl_n2801), .A (n_535));
NOR3_X4 sgo__sro_c361 (.ZN (n_1119), .A1 (sgo__sro_n191), .A2 (n_979), .A3 (n_954));
AND2_X1 sgo__sro_c554 (.ZN (n_555), .A1 (slo__sro_n764), .A2 (n_217));
XNOR2_X1 sgo__sro_c555 (.ZN (n_240), .A (slo__sro_n764), .B (sgo__sro_n293));
INV_X1 sgo__sro_c583 (.ZN (sgo__sro_n310), .A (n_592));
NOR2_X2 sgo__c494 (.ZN (sgo__n265), .A1 (n_1214), .A2 (n_1221));
INV_X1 sgo__c496 (.ZN (n_1213), .A (sgo__n265));
AND2_X4 slo__c750 (.ZN (slo__n432), .A1 (n_1245), .A2 (n_8));
OAI21_X2 slo__sro_c619 (.ZN (slo__sro_n332), .A (slo__sro_n333), .B1 (n_1123), .B2 (n_1365));
AND2_X1 slo__sro_c660 (.ZN (n_411), .A1 (n_94), .A2 (n_92));
XNOR2_X2 slo__sro_c661 (.ZN (n_409), .A (n_94), .B (slo__sro_n366));
XNOR2_X2 slo__mro_c673 (.ZN (\aggregated_res[14] [56] ), .A (n_1073), .B (n_1071));
AND3_X2 slo__xsl_c708 (.ZN (n_738), .A1 (sgo__sro_n309), .A2 (n_739), .A3 (n_767));
INV_X1 slo__sro_c754 (.ZN (slo__sro_n442), .A (n_1215));
XNOR2_X2 slo__sro_c755 (.ZN (\aggregated_res[14] [49] ), .A (n_1213), .B (slo__sro_n442));
INV_X4 slo__sro_c770 (.ZN (n_7), .A (slo__sro_n460));
OAI21_X1 slo__sro_c776 (.ZN (slo__sro_n467), .A (n_936), .B1 (n_546), .B2 (n_544));
NAND2_X2 slo__sro_c777 (.ZN (slo__sro_n466), .A1 (slo__sro_n467), .A2 (slo__sro_n468));
XNOR2_X1 slo__sro_c778 (.ZN (slo__sro_n465), .A (n_936), .B (n_544));
XNOR2_X2 slo__sro_c779 (.ZN (slo__sro_n464), .A (n_546), .B (slo__sro_n465));
XNOR2_X1 slo__sro_c811 (.ZN (\aggregated_res[14] [55] ), .A (n_1029), .B (slo__sro_n499));
OAI21_X2 slo__sro_c822 (.ZN (n_616), .A (opt_ipo_n2338), .B1 (n_507), .B2 (opt_ipo_n1965));
OAI21_X1 slo__sro_c842 (.ZN (slo__sro_n535), .A (n_657), .B1 (n_951), .B2 (n_649));
INV_X1 slo__sro_c851 (.ZN (slo__sro_n546), .A (n_531));
INV_X2 slo__sro_c852 (.ZN (slo__sro_n545), .A (n_515));
NAND2_X2 slo__sro_c853 (.ZN (slo__sro_n544), .A1 (slo__sro_n545), .A2 (slo__sro_n546));
NAND3_X2 slo__sro_c854 (.ZN (n_509), .A1 (slo__sro_n544), .A2 (opt_ipo_n1940), .A3 (n_513));
AND2_X1 slo__sro_c881 (.ZN (slo__sro_n568), .A1 (n_1134), .A2 (n_1149));
NOR2_X1 slo__sro_c882 (.ZN (slo__sro_n567), .A1 (n_1195), .A2 (slo__sro_n568));
INV_X4 slo__sro_c902 (.ZN (slo__sro_n589), .A (n_391));
NAND2_X4 slo__sro_c903 (.ZN (slo__sro_n588), .A1 (slo__sro_n589), .A2 (n_525));
AOI21_X4 slo__sro_c904 (.ZN (slo__sro_n587), .A (slo__sro_n588), .B1 (opt_ipo_n1948), .B2 (n_390));
XNOR2_X2 slo__sro_c915 (.ZN (\aggregated_res[14] [47] ), .A (n_1007), .B (slo__sro_n604));
INV_X2 slo__c967 (.ZN (sgo__sro_n14), .A (slo__n651));
OAI21_X1 slo__sro_c1018 (.ZN (slo__sro_n694), .A (n_239), .B1 (n_260), .B2 (slo__sro_n1798));
NAND2_X1 slo__sro_c1019 (.ZN (n_553), .A1 (slo__sro_n694), .A2 (slo__sro_n695));
XNOR2_X2 slo__sro_c1020 (.ZN (slo__sro_n693), .A (n_239), .B (slo__sro_n1798));
XNOR2_X2 slo__sro_c1021 (.ZN (slo__sro_n692), .A (slo__sro_n693), .B (n_260));
NAND2_X1 slo__sro_c1032 (.ZN (slo__sro_n707), .A1 (slo__sro_n927), .A2 (n_358));
NOR2_X1 slo__sro_c1033 (.ZN (slo__sro_n706), .A1 (slo__sro_n927), .A2 (n_358));
OAI21_X4 slo__sro_c1034 (.ZN (n_663), .A (slo__sro_n707), .B1 (slo__sro_n708), .B2 (slo__sro_n706));
XNOR2_X2 slo__sro_c1035 (.ZN (slo__sro_n705), .A (n_358), .B (slo__sro_n927));
XNOR2_X2 slo__sro_c1036 (.ZN (slo__sro_n704), .A (slo__sro_n705), .B (n_335));
OAI21_X1 slo__sro_c1046 (.ZN (slo__sro_n718), .A (n_498), .B1 (n_216), .B2 (n_214));
NAND2_X1 slo__sro_c1047 (.ZN (n_219), .A1 (slo__sro_n718), .A2 (slo__sro_n719));
XNOR2_X1 slo__sro_c1048 (.ZN (slo__sro_n717), .A (n_498), .B (n_214));
XNOR2_X1 slo__sro_c1049 (.ZN (slo__sro_n716), .A (slo__sro_n717), .B (n_216));
NAND2_X1 slo__sro_c1058 (.ZN (slo__sro_n729), .A1 (n_173), .A2 (n_188));
NOR2_X1 slo__sro_c1059 (.ZN (slo__sro_n728), .A1 (n_173), .A2 (n_188));
OAI21_X1 slo__sro_c1060 (.ZN (n_473), .A (slo__sro_n729), .B1 (slo__sro_n730), .B2 (slo__sro_n728));
XNOR2_X2 slo__sro_c1061 (.ZN (slo__sro_n727), .A (n_173), .B (n_188));
XNOR2_X2 slo__sro_c1062 (.ZN (slo__sro_n726), .A (slo__sro_n791), .B (slo__sro_n727));
NAND2_X1 slo__sro_c1076 (.ZN (slo__sro_n744), .A1 (n_211), .A2 (n_213));
NOR2_X1 slo__sro_c1077 (.ZN (slo__sro_n743), .A1 (n_213), .A2 (n_211));
OAI21_X1 slo__sro_c1078 (.ZN (n_237), .A (slo__sro_n744), .B1 (slo__sro_n745), .B2 (slo__sro_n743));
XNOR2_X1 slo__sro_c1079 (.ZN (slo__sro_n742), .A (n_211), .B (n_213));
XNOR2_X1 slo__sro_c1080 (.ZN (n_236), .A (slo__sro_n742), .B (n_215));
NAND2_X1 slo__sro_c1090 (.ZN (slo__sro_n754), .A1 (n_221), .A2 (n_223));
NOR2_X1 slo__sro_c1091 (.ZN (slo__sro_n753), .A1 (n_221), .A2 (n_223));
OAI21_X1 slo__sro_c1092 (.ZN (slo__sro_n752), .A (slo__sro_n754), .B1 (slo__sro_n755), .B2 (slo__sro_n753));
XNOR2_X1 slo__sro_c1093 (.ZN (slo__sro_n751), .A (n_221), .B (n_223));
XNOR2_X1 slo__sro_c1094 (.ZN (slo__sro_n750), .A (slo__sro_n751), .B (slo__sro_n777));
NAND2_X1 slo__sro_c1104 (.ZN (slo__sro_n767), .A1 (n_236), .A2 (n_232));
AOI22_X1 slo__sro_c1105 (.ZN (slo__sro_n766), .A1 (n_236), .A2 (n_234), .B1 (n_234), .B2 (n_232));
NAND2_X2 slo__sro_c1106 (.ZN (n_239), .A1 (slo__sro_n766), .A2 (slo__sro_n767));
XNOR2_X1 slo__sro_c1107 (.ZN (slo__sro_n765), .A (n_234), .B (n_232));
XNOR2_X1 slo__sro_c1108 (.ZN (slo__sro_n764), .A (slo__sro_n765), .B (n_236));
NAND2_X1 slo__sro_c1120 (.ZN (slo__sro_n779), .A1 (n_205), .A2 (p_15[24]));
NAND2_X1 slo__sro_c1121 (.ZN (slo__sro_n778), .A1 (n_207), .A2 (n_205));
NAND3_X1 slo__sro_c1122 (.ZN (slo__sro_n777), .A1 (slo__sro_n780), .A2 (slo__sro_n778), .A3 (slo__sro_n779));
XNOR2_X1 slo__sro_c1123 (.ZN (slo__sro_n776), .A (n_205), .B (p_15[24]));
XNOR2_X1 slo__sro_c1124 (.ZN (n_228), .A (slo__sro_n776), .B (n_207));
OAI21_X1 slo__sro_c1136 (.ZN (slo__sro_n792), .A (n_433), .B1 (n_170), .B2 (n_162));
NAND2_X1 slo__sro_c1137 (.ZN (slo__sro_n791), .A1 (slo__sro_n793), .A2 (slo__sro_n792));
XNOR2_X1 slo__sro_c1138 (.ZN (slo__sro_n790), .A (n_170), .B (n_162));
XNOR2_X2 slo__sro_c1139 (.ZN (n_174), .A (slo__sro_n790), .B (n_433));
AOI22_X1 slo__sro_c1150 (.ZN (slo__sro_n803), .A1 (n_1146), .A2 (slo__sro_n1688), .B1 (slo__sro_n1688), .B2 (n_1144));
NAND2_X1 slo__sro_c1151 (.ZN (n_709), .A1 (slo__sro_n803), .A2 (slo__sro_n804));
XNOR2_X1 slo__sro_c1152 (.ZN (slo__sro_n802), .A (slo__sro_n1688), .B (n_1144));
XNOR2_X1 slo__sro_c1153 (.ZN (n_708), .A (slo__sro_n802), .B (n_1146));
NOR2_X1 slo__sro_c1171 (.ZN (slo__sro_n819), .A1 (n_878), .A2 (n_676));
INV_X1 slo__sro_c1172 (.ZN (slo__sro_n818), .A (slo__sro_n819));
NAND2_X1 slo__sro_c1173 (.ZN (slo__sro_n817), .A1 (slo__sro_n818), .A2 (n_682));
NAND2_X1 slo__sro_c1174 (.ZN (slo__sro_n816), .A1 (slo__sro_n817), .A2 (slo__sro_n820));
XNOR2_X1 slo__sro_c1175 (.ZN (slo__sro_n815), .A (n_878), .B (n_676));
XNOR2_X1 slo__sro_c1176 (.ZN (slo__sro_n814), .A (n_682), .B (slo__sro_n815));
NAND2_X1 slo__sro_c1192 (.ZN (slo__sro_n834), .A1 (n_882), .A2 (n_1079));
NOR2_X1 slo__sro_c1193 (.ZN (slo__sro_n833), .A1 (n_882), .A2 (n_1079));
OAI21_X1 slo__sro_c1194 (.ZN (n_1142), .A (slo__sro_n834), .B1 (slo__sro_n835), .B2 (slo__sro_n833));
XNOR2_X1 slo__sro_c1195 (.ZN (slo__sro_n832), .A (n_882), .B (n_1079));
XNOR2_X1 slo__sro_c1196 (.ZN (n_682), .A (slo__sro_n832), .B (n_1082));
OAI21_X1 slo__sro_c1206 (.ZN (slo__sro_n841), .A (n_1088), .B1 (n_688), .B2 (n_684));
NAND2_X1 slo__sro_c1207 (.ZN (n_1146), .A1 (slo__sro_n842), .A2 (slo__sro_n841));
XNOR2_X1 slo__sro_c1208 (.ZN (slo__sro_n840), .A (n_1088), .B (n_684));
XNOR2_X1 slo__sro_c1209 (.ZN (n_690), .A (slo__sro_n840), .B (n_688));
OAI21_X2 slo__sro_c1218 (.ZN (slo__sro_n848), .A (n_18), .B1 (n_20), .B2 (n_51));
NAND2_X1 slo__sro_c1219 (.ZN (slo__sro_n847), .A1 (slo__sro_n848), .A2 (slo__sro_n849));
XNOR2_X1 slo__sro_c1220 (.ZN (slo__sro_n846), .A (n_51), .B (n_18));
XNOR2_X1 slo__sro_c1221 (.ZN (n_22), .A (slo__sro_n846), .B (n_20));
OAI21_X1 slo__sro_c1230 (.ZN (slo__sro_n855), .A (n_1087), .B1 (n_1084), .B2 (slo__sro_n814));
NAND2_X1 slo__sro_c1231 (.ZN (n_1144), .A1 (slo__sro_n855), .A2 (slo__sro_n856));
XNOR2_X1 slo__sro_c1232 (.ZN (slo__sro_n854), .A (slo__sro_n814), .B (n_1084));
XNOR2_X1 slo__sro_c1233 (.ZN (n_688), .A (slo__sro_n854), .B (n_1087));
OAI21_X1 slo__sro_c1314 (.ZN (slo__sro_n902), .A (slo__sro_n917), .B1 (n_416), .B2 (n_414));
XNOR2_X2 slo__sro_c1316 (.ZN (slo__sro_n901), .A (slo__sro_n917), .B (n_414));
INV_X1 slo__xsl_c1260 (.ZN (slo__xsl_n869), .A (n_767));
INV_X1 CLOCK_slo__sro_c3950 (.ZN (CLOCK_slo__sro_n2898), .A (n_518));
NAND2_X1 slo__sro_c1326 (.ZN (slo__sro_n909), .A1 (n_312), .A2 (n_314));
NOR2_X1 slo__sro_c1327 (.ZN (slo__sro_n908), .A1 (n_312), .A2 (n_314));
OAI21_X1 slo__sro_c1328 (.ZN (n_329), .A (slo__sro_n909), .B1 (slo__sro_n910), .B2 (slo__sro_n908));
XNOR2_X1 slo__sro_c1329 (.ZN (slo__sro_n907), .A (n_312), .B (n_314));
XNOR2_X1 slo__sro_c1330 (.ZN (n_328), .A (slo__sro_n907), .B (n_322));
OAI21_X2 slo__sro_c1340 (.ZN (slo__sro_n918), .A (n_361), .B1 (n_359), .B2 (n_384));
NAND2_X2 slo__sro_c1341 (.ZN (slo__sro_n917), .A1 (slo__sro_n918), .A2 (slo__sro_n919));
XNOR2_X1 slo__sro_c1342 (.ZN (slo__sro_n916), .A (n_359), .B (n_361));
XNOR2_X1 slo__sro_c1343 (.ZN (slo__sro_n915), .A (slo__sro_n916), .B (n_384));
NAND2_X1 slo__sro_c1352 (.ZN (slo__sro_n930), .A1 (n_333), .A2 (n_331));
NAND2_X1 slo__sro_c1353 (.ZN (slo__sro_n929), .A1 (n_333), .A2 (n_356));
NAND3_X2 slo__sro_c1354 (.ZN (n_361), .A1 (slo__sro_n929), .A2 (slo__sro_n931), .A3 (slo__sro_n930));
XNOR2_X1 slo__sro_c1355 (.ZN (slo__sro_n928), .A (n_333), .B (n_331));
XNOR2_X2 slo__sro_c1356 (.ZN (slo__sro_n927), .A (slo__sro_n928), .B (n_356));
INV_X1 slo__sro_c1368 (.ZN (slo__sro_n943), .A (n_293));
NAND2_X1 slo__sro_c1369 (.ZN (slo__sro_n942), .A1 (n_295), .A2 (n_293));
NAND2_X1 slo__sro_c1370 (.ZN (slo__sro_n941), .A1 (slo__sro_n944), .A2 (slo__sro_n943));
NAND2_X1 slo__sro_c1371 (.ZN (slo__sro_n940), .A1 (slo__sro_n941), .A2 (n_291));
NAND2_X2 slo__sro_c1372 (.ZN (n_323), .A1 (slo__sro_n940), .A2 (slo__sro_n942));
XNOR2_X1 slo__sro_c1373 (.ZN (slo__sro_n939), .A (n_295), .B (n_293));
XNOR2_X1 slo__sro_c1374 (.ZN (n_322), .A (slo__sro_n939), .B (n_291));
OAI21_X1 slo__sro_c1386 (.ZN (slo__sro_n953), .A (n_305), .B1 (n_326), .B2 (n_328));
NAND2_X1 slo__sro_c1387 (.ZN (n_333), .A1 (slo__sro_n953), .A2 (slo__sro_n954));
XNOR2_X1 slo__sro_c1388 (.ZN (slo__sro_n952), .A (n_305), .B (n_328));
XNOR2_X1 slo__sro_c1389 (.ZN (slo__sro_n951), .A (slo__sro_n952), .B (n_326));
OAI21_X1 slo__sro_c1398 (.ZN (slo__sro_n960), .A (slo__sro_n1476), .B1 (n_1068), .B2 (n_1031));
NAND2_X1 slo__sro_c1399 (.ZN (n_595), .A1 (slo__sro_n960), .A2 (slo__sro_n961));
XNOR2_X1 slo__sro_c1400 (.ZN (slo__sro_n959), .A (slo__sro_n1476), .B (n_1031));
XNOR2_X2 slo__sro_c1401 (.ZN (n_1078), .A (slo__sro_n959), .B (n_1068));
NAND2_X1 slo__sro_c1410 (.ZN (slo__sro_n967), .A1 (n_1006), .A2 (n_1028));
NOR2_X1 slo__sro_c1411 (.ZN (slo__sro_n966), .A1 (n_1006), .A2 (n_1028));
OAI21_X1 slo__sro_c1412 (.ZN (n_593), .A (slo__sro_n967), .B1 (slo__sro_n968), .B2 (slo__sro_n966));
XNOR2_X1 slo__sro_c1413 (.ZN (slo__sro_n965), .A (n_1006), .B (n_1028));
XNOR2_X1 slo__sro_c1414 (.ZN (n_1068), .A (n_1015), .B (slo__sro_n965));
INV_X1 slo__sro_c1504 (.ZN (slo__sro_n1024), .A (n_1037));
NAND2_X1 slo__sro_c1506 (.ZN (slo__sro_n1022), .A1 (slo__sro_n1024), .A2 (slo__sro_n1025));
INV_X1 slo__xsl_c1447 (.ZN (slo__xsl_n988), .A (n_801));
AND2_X4 slo__xsl_c1450 (.ZN (n_801), .A1 (n_793), .A2 (n_711));
NAND2_X1 slo__sro_c1508 (.ZN (n_1088), .A1 (slo__sro_n1023), .A2 (slo__sro_n1021));
XNOR2_X1 slo__sro_c1509 (.ZN (slo__sro_n1020), .A (n_1037), .B (n_1042));
XNOR2_X1 slo__sro_c1510 (.ZN (n_670), .A (slo__sro_n1020), .B (n_1035));
OAI21_X1 slo__sro_c1522 (.ZN (slo__sro_n1033), .A (slo__sro_n1622), .B1 (slo__sro_n1040), .B2 (n_1043));
NAND2_X1 slo__sro_c1523 (.ZN (n_1092), .A1 (slo__sro_n1033), .A2 (slo__sro_n1034));
XNOR2_X1 slo__sro_c1524 (.ZN (slo__sro_n1032), .A (slo__sro_n1622), .B (n_1043));
XNOR2_X1 slo__sro_c1525 (.ZN (n_674), .A (slo__sro_n1032), .B (slo__sro_n1040));
INV_X1 slo__sro_c1536 (.ZN (slo__sro_n1045), .A (n_666));
NAND2_X1 slo__sro_c1537 (.ZN (slo__sro_n1044), .A1 (n_666), .A2 (n_668));
NAND2_X1 slo__sro_c1538 (.ZN (slo__sro_n1043), .A1 (slo__sro_n1045), .A2 (slo__sro_n1046));
NAND2_X1 slo__sro_c1539 (.ZN (slo__sro_n1042), .A1 (n_670), .A2 (slo__sro_n1043));
NAND2_X1 slo__sro_c1540 (.ZN (n_1089), .A1 (slo__sro_n1042), .A2 (slo__sro_n1044));
XNOR2_X1 slo__sro_c1541 (.ZN (slo__sro_n1041), .A (n_666), .B (n_668));
XNOR2_X1 slo__sro_c1542 (.ZN (slo__sro_n1040), .A (n_670), .B (slo__sro_n1041));
AND2_X1 slo__sro_c1607 (.ZN (slo__sro_n1091), .A1 (n_1302), .A2 (n_1304));
INV_X1 slo__xsl_c1566 (.ZN (slo__xsl_n1064), .A (n_1192));
INV_X1 slo__xsl_c1567 (.ZN (slo__xsl_n1063), .A (slo__xsl_n1064));
NOR3_X2 slo__sro_c1608 (.ZN (\aggregated_res[14] [53] ), .A1 (n_1299), .A2 (n_1294), .A3 (slo__sro_n1091));
NAND2_X1 slo__sro_c1635 (.ZN (n_637), .A1 (slo__sro_n1107), .A2 (slo__sro_n1108));
XNOR2_X2 slo__sro_c1636 (.ZN (slo__sro_n1106), .A (slo__sro_n1341), .B (n_632));
XNOR2_X2 slo__sro_c1637 (.ZN (n_1033), .A (slo__sro_n1106), .B (slo__sro_n1130));
NAND2_X1 slo__sro_c1655 (.ZN (slo__sro_n1121), .A1 (n_581), .A2 (n_575));
NAND2_X1 slo__sro_c1656 (.ZN (slo__sro_n1120), .A1 (n_581), .A2 (n_892));
NAND3_X1 slo__sro_c1657 (.ZN (n_605), .A1 (slo__sro_n1121), .A2 (slo__sro_n1120), .A3 (slo__sro_n1122));
XNOR2_X2 slo__sro_c1658 (.ZN (slo__sro_n1119), .A (n_892), .B (n_575));
XNOR2_X2 slo__sro_c1659 (.ZN (slo__sro_n1118), .A (slo__sro_n1119), .B (n_581));
NAND2_X1 slo__sro_c1669 (.ZN (slo__sro_n1134), .A1 (n_613), .A2 (n_630));
NOR2_X1 slo__sro_c1670 (.ZN (slo__sro_n1133), .A1 (n_613), .A2 (n_630));
OAI21_X1 slo__sro_c1671 (.ZN (slo__sro_n1132), .A (slo__sro_n1134), .B1 (slo__sro_n1133), .B2 (slo__sro_n1135));
XNOR2_X1 slo__sro_c1672 (.ZN (slo__sro_n1131), .A (n_613), .B (n_630));
XNOR2_X2 slo__sro_c1673 (.ZN (slo__sro_n1130), .A (slo__sro_n1131), .B (n_611));
NAND2_X1 slo__sro_c1694 (.ZN (slo__sro_n1154), .A1 (slo__sro_n1118), .A2 (n_888));
NOR2_X1 slo__sro_c1695 (.ZN (slo__sro_n1153), .A1 (slo__sro_n1118), .A2 (n_888));
OAI21_X1 slo__sro_c1696 (.ZN (slo__sro_n1152), .A (slo__sro_n1154), .B1 (slo__sro_n1153), .B2 (slo__sro_n1155));
XNOR2_X1 slo__sro_c1697 (.ZN (slo__sro_n1151), .A (slo__sro_n1118), .B (n_888));
XNOR2_X1 slo__sro_c1698 (.ZN (slo__sro_n1150), .A (slo__sro_n1151), .B (slo__sro_n1357));
AOI21_X4 slo__sro_c1708 (.ZN (\aggregated_res[14] [59] ), .A (slo__sro_n1166), .B1 (n_1039), .B2 (n_1369));
OR2_X1 slo__sro_c1725 (.ZN (slo__sro_n1184), .A1 (p_15[8]), .A2 (p_3[8]));
NAND2_X1 slo__sro_c1726 (.ZN (slo__sro_n1183), .A1 (slo__sro_n1184), .A2 (n_14));
NAND2_X1 slo__sro_c1727 (.ZN (n_51), .A1 (slo__sro_n1183), .A2 (slo__sro_n1185));
XNOR2_X1 slo__sro_c1728 (.ZN (slo__sro_n1182), .A (p_15[8]), .B (p_3[8]));
XNOR2_X1 slo__sro_c1729 (.ZN (slo__sro_n1181), .A (slo__sro_n1182), .B (n_14));
OAI21_X1 slo__sro_c1739 (.ZN (slo__sro_n1195), .A (n_438), .B1 (n_440), .B2 (n_777));
NAND2_X1 slo__sro_c1740 (.ZN (n_832), .A1 (slo__sro_n1195), .A2 (slo__sro_n1196));
XNOR2_X2 slo__sro_c1741 (.ZN (slo__sro_n1194), .A (n_777), .B (n_438));
XNOR2_X2 slo__sro_c1742 (.ZN (slo__sro_n1193), .A (n_440), .B (slo__sro_n1194));
INV_X1 slo__sro_c1761 (.ZN (slo__sro_n1211), .A (n_408));
NAND2_X1 slo__sro_c1762 (.ZN (slo__sro_n1210), .A1 (n_685), .A2 (n_408));
NAND2_X1 slo__sro_c1763 (.ZN (slo__sro_n1209), .A1 (slo__sro_n1212), .A2 (slo__sro_n1211));
NAND2_X2 slo__sro_c1764 (.ZN (slo__sro_n1208), .A1 (n_689), .A2 (slo__sro_n1209));
NAND2_X2 slo__sro_c1765 (.ZN (n_777), .A1 (slo__sro_n1210), .A2 (slo__sro_n1208));
XNOR2_X1 slo__sro_c1766 (.ZN (slo__sro_n1207), .A (n_685), .B (n_408));
XNOR2_X2 slo__sro_c1767 (.ZN (n_414), .A (n_689), .B (slo__sro_n1207));
OAI21_X1 slo__sro_c1809 (.ZN (slo__sro_n1243), .A (p_14[31]), .B1 (p_12[31]), .B2 (p_13[31]));
NAND2_X2 slo__sro_c1810 (.ZN (n_779), .A1 (slo__sro_n1243), .A2 (slo__sro_n1244));
XNOR2_X1 slo__sro_c1811 (.ZN (slo__sro_n1242), .A (p_14[31]), .B (p_13[31]));
XNOR2_X1 slo__sro_c1812 (.ZN (slo__sro_n1241), .A (slo__sro_n1242), .B (p_12[31]));
NAND2_X1 slo__sro_c1828 (.ZN (slo__sro_n1257), .A1 (n_516), .A2 (n_512));
NAND2_X1 slo__sro_c1829 (.ZN (slo__sro_n1256), .A1 (n_516), .A2 (n_493));
NAND3_X1 slo__sro_c1830 (.ZN (slo__sro_n1255), .A1 (slo__sro_n1257), .A2 (slo__sro_n1256), .A3 (slo__sro_n1258));
XNOR2_X2 slo__sro_c1831 (.ZN (slo__sro_n1254), .A (n_493), .B (n_512));
XNOR2_X2 slo__sro_c1832 (.ZN (slo__sro_n1253), .A (slo__sro_n1254), .B (n_516));
NAND2_X2 slo__sro_c1843 (.ZN (n_936), .A1 (CLOCK_slo__sro_n2895), .A2 (slo__sro_n1270));
XNOR2_X1 slo__sro_c1844 (.ZN (slo__sro_n1268), .A (n_495), .B (n_518));
XNOR2_X2 slo__sro_c1845 (.ZN (slo__sro_n1267), .A (slo__sro_n1268), .B (slo__sro_n1253));
INV_X1 slo__sro_c1854 (.ZN (slo__sro_n1281), .A (n_445));
NAND2_X1 slo__sro_c1855 (.ZN (slo__sro_n1280), .A1 (n_445), .A2 (n_174));
NAND2_X1 slo__sro_c1856 (.ZN (slo__sro_n1279), .A1 (slo__sro_n1282), .A2 (slo__sro_n1281));
NAND2_X1 slo__sro_c1857 (.ZN (slo__sro_n1278), .A1 (slo__sro_n1279), .A2 (n_176));
NAND2_X1 slo__sro_c1858 (.ZN (n_457), .A1 (slo__sro_n1278), .A2 (slo__sro_n1280));
XNOR2_X2 slo__sro_c1859 (.ZN (slo__sro_n1277), .A (n_445), .B (n_174));
XNOR2_X2 slo__sro_c1860 (.ZN (n_455), .A (slo__sro_n1277), .B (n_176));
NAND2_X1 slo__sro_c1872 (.ZN (slo__sro_n1291), .A1 (n_129), .A2 (n_131));
NOR2_X1 slo__sro_c1873 (.ZN (slo__sro_n1290), .A1 (n_129), .A2 (n_131));
OAI21_X2 slo__sro_c1874 (.ZN (n_433), .A (slo__sro_n1291), .B1 (slo__sro_n1292), .B2 (slo__sro_n1290));
XNOR2_X1 slo__sro_c1875 (.ZN (slo__sro_n1289), .A (n_129), .B (n_131));
XNOR2_X1 slo__sro_c1876 (.ZN (n_152), .A (slo__sro_n1289), .B (n_135));
NAND2_X1 slo__sro_c1886 (.ZN (slo__sro_n1299), .A1 (n_443), .A2 (n_172));
NOR2_X1 slo__sro_c1887 (.ZN (slo__sro_n1298), .A1 (n_172), .A2 (n_443));
OAI21_X1 slo__sro_c1888 (.ZN (n_177), .A (slo__sro_n1299), .B1 (slo__sro_n1300), .B2 (slo__sro_n1298));
XNOR2_X1 slo__sro_c1889 (.ZN (slo__sro_n1297), .A (n_172), .B (n_443));
XNOR2_X2 slo__sro_c1890 (.ZN (n_176), .A (slo__sro_n1297), .B (n_435));
NAND2_X1 slo__sro_c1929 (.ZN (slo__sro_n1333), .A1 (n_16), .A2 (n_1176));
NOR2_X1 slo__sro_c1930 (.ZN (slo__sro_n1332), .A1 (n_16), .A2 (n_1176));
OAI21_X1 slo__sro_c1931 (.ZN (n_1161), .A (slo__sro_n1333), .B1 (slo__sro_n1332), .B2 (slo__sro_n1334));
XNOR2_X2 slo__sro_c1932 (.ZN (slo__sro_n1331), .A (n_16), .B (n_1176));
XNOR2_X2 slo__sro_c1933 (.ZN (n_716), .A (slo__sro_n1331), .B (n_699));
OAI21_X2 slo__sro_c1943 (.ZN (slo__sro_n1342), .A (n_591), .B1 (n_612), .B2 (n_610));
NAND2_X2 slo__sro_c1944 (.ZN (slo__sro_n1341), .A1 (slo__sro_n1342), .A2 (slo__sro_n1343));
XNOR2_X2 slo__sro_c1945 (.ZN (slo__sro_n1340), .A (n_612), .B (n_591));
XNOR2_X2 slo__sro_c1946 (.ZN (slo__sro_n1339), .A (slo__sro_n1340), .B (n_610));
AOI22_X1 slo__sro_c1959 (.ZN (slo__sro_n1358), .A1 (n_1012), .A2 (n_1023), .B1 (n_1023), .B2 (n_1010));
NAND2_X1 slo__sro_c1960 (.ZN (slo__sro_n1357), .A1 (slo__sro_n1358), .A2 (slo__sro_n1359));
XNOR2_X1 slo__sro_c1961 (.ZN (slo__sro_n1356), .A (n_1023), .B (n_1010));
XNOR2_X1 slo__sro_c1962 (.ZN (slo__sro_n1355), .A (slo__sro_n1356), .B (n_1012));
INV_X1 slo__sro_c1971 (.ZN (slo__sro_n1371), .A (n_584));
NAND2_X1 slo__sro_c1972 (.ZN (slo__sro_n1370), .A1 (n_1014), .A2 (n_584));
NAND2_X1 slo__sro_c1973 (.ZN (slo__sro_n1369), .A1 (slo__sro_n1372), .A2 (slo__sro_n1371));
NAND2_X1 slo__sro_c1974 (.ZN (slo__sro_n1368), .A1 (slo__sro_n1379), .A2 (slo__sro_n1369));
NAND2_X1 slo__sro_c1975 (.ZN (n_591), .A1 (slo__sro_n1368), .A2 (slo__sro_n1370));
XNOR2_X1 slo__sro_c1976 (.ZN (slo__sro_n1367), .A (n_1014), .B (n_584));
XNOR2_X1 slo__sro_c1977 (.ZN (n_1031), .A (slo__sro_n1379), .B (slo__sro_n1367));
NAND2_X1 slo__sro_c1989 (.ZN (slo__sro_n1383), .A1 (n_574), .A2 (n_890));
OR2_X1 slo__sro_c1990 (.ZN (slo__sro_n1382), .A1 (n_574), .A2 (n_890));
NAND2_X1 slo__sro_c1991 (.ZN (slo__sro_n1381), .A1 (slo__sro_n1355), .A2 (slo__sro_n1382));
NAND2_X1 slo__sro_c1992 (.ZN (n_587), .A1 (slo__sro_n1381), .A2 (slo__sro_n1383));
XNOR2_X1 slo__sro_c1993 (.ZN (slo__sro_n1380), .A (n_574), .B (n_890));
XNOR2_X1 slo__sro_c1994 (.ZN (slo__sro_n1379), .A (slo__sro_n1355), .B (slo__sro_n1380));
OAI21_X1 slo__sro_c2005 (.ZN (slo__sro_n1395), .A (n_966), .B1 (n_897), .B2 (n_965));
NAND2_X1 slo__sro_c2006 (.ZN (n_1012), .A1 (slo__sro_n1395), .A2 (slo__sro_n1396));
XNOR2_X1 slo__sro_c2007 (.ZN (slo__sro_n1394), .A (n_965), .B (n_966));
XNOR2_X1 slo__sro_c2008 (.ZN (slo__sro_n1393), .A (slo__sro_n1394), .B (n_897));
NAND2_X1 slo__sro_c2017 (.ZN (slo__sro_n1404), .A1 (n_716), .A2 (n_701));
NOR2_X1 slo__sro_c2018 (.ZN (slo__sro_n1403), .A1 (n_716), .A2 (n_701));
OAI21_X1 slo__sro_c2019 (.ZN (slo__sro_n1402), .A (slo__sro_n1404), .B1 (slo__sro_n1403), .B2 (slo__sro_n1405));
XNOR2_X1 slo__sro_c2020 (.ZN (slo__sro_n1401), .A (n_716), .B (n_701));
XNOR2_X1 slo__sro_c2021 (.ZN (n_720), .A (slo__sro_n1401), .B (n_703));
NAND2_X1 slo__sro_c2074 (.ZN (slo__sro_n1441), .A1 (n_330), .A2 (n_307));
NOR2_X1 slo__sro_c2075 (.ZN (slo__sro_n1440), .A1 (n_307), .A2 (n_330));
OAI21_X1 slo__sro_c2076 (.ZN (n_335), .A (slo__sro_n1441), .B1 (slo__sro_n1442), .B2 (slo__sro_n1440));
XNOR2_X2 slo__sro_c2077 (.ZN (slo__sro_n1439), .A (n_330), .B (n_307));
XNOR2_X2 slo__sro_c2078 (.ZN (n_334), .A (slo__sro_n1439), .B (n_309));
INV_X1 slo__sro_c2133 (.ZN (slo__sro_n1480), .A (n_566));
NAND2_X1 slo__sro_c2134 (.ZN (slo__sro_n1479), .A1 (n_566), .A2 (n_970));
NAND2_X1 slo__sro_c2135 (.ZN (slo__sro_n1478), .A1 (slo__sro_n1480), .A2 (slo__sro_n1481));
NAND2_X1 slo__sro_c2136 (.ZN (slo__sro_n1477), .A1 (n_568), .A2 (slo__sro_n1478));
NAND2_X1 slo__sro_c2137 (.ZN (slo__sro_n1476), .A1 (slo__sro_n1477), .A2 (slo__sro_n1479));
XNOR2_X1 slo__sro_c2138 (.ZN (slo__sro_n1475), .A (n_566), .B (n_970));
XNOR2_X1 slo__sro_c2139 (.ZN (slo__sro_n1474), .A (n_568), .B (slo__sro_n1475));
NAND2_X1 slo__sro_c2153 (.ZN (slo__sro_n1496), .A1 (n_564), .A2 (n_562));
NOR2_X1 slo__sro_c2154 (.ZN (slo__sro_n1495), .A1 (n_564), .A2 (n_562));
OAI21_X1 slo__sro_c2155 (.ZN (n_1015), .A (slo__sro_n1496), .B1 (slo__sro_n1497), .B2 (slo__sro_n1495));
XNOR2_X1 slo__sro_c2156 (.ZN (slo__sro_n1494), .A (n_564), .B (n_562));
XNOR2_X1 slo__sro_c2157 (.ZN (n_568), .A (slo__sro_n1494), .B (n_973));
INV_X1 slo__sro_c2189 (.ZN (slo__sro_n1522), .A (n_749));
NAND2_X1 slo__sro_c2190 (.ZN (slo__sro_n1521), .A1 (n_747), .A2 (n_758));
NOR2_X1 slo__sro_c2191 (.ZN (slo__sro_n1520), .A1 (n_758), .A2 (n_747));
OAI21_X1 slo__sro_c2192 (.ZN (n_763), .A (slo__sro_n1521), .B1 (slo__sro_n1522), .B2 (slo__sro_n1520));
XNOR2_X2 slo__sro_c2193 (.ZN (slo__sro_n1519), .A (n_758), .B (n_747));
XNOR2_X2 slo__sro_c2194 (.ZN (n_762), .A (slo__sro_n1519), .B (n_749));
OAI21_X1 slo__sro_c2223 (.ZN (slo__sro_n1539), .A (n_891), .B1 (n_496), .B2 (n_494));
NAND2_X1 slo__sro_c2224 (.ZN (slo__sro_n1538), .A1 (slo__sro_n1539), .A2 (slo__sro_n1540));
XNOR2_X2 slo__sro_c2225 (.ZN (slo__sro_n1537), .A (n_891), .B (n_494));
XNOR2_X2 slo__sro_c2226 (.ZN (n_938), .A (slo__sro_n1537), .B (n_496));
OAI21_X1 slo__sro_c2240 (.ZN (slo__sro_n1549), .A (n_876), .B1 (n_886), .B2 (n_492));
NAND2_X1 slo__sro_c2241 (.ZN (slo__sro_n1548), .A1 (slo__sro_n1549), .A2 (slo__sro_n1550));
XNOR2_X1 slo__sro_c2242 (.ZN (slo__sro_n1547), .A (n_876), .B (n_886));
XNOR2_X1 slo__sro_c2243 (.ZN (n_496), .A (slo__sro_n1547), .B (n_492));
OR2_X1 slo__sro_c2277 (.ZN (slo__sro_n1571), .A1 (p_15[14]), .A2 (p_6[14]));
NAND2_X1 slo__sro_c2278 (.ZN (slo__sro_n1570), .A1 (n_191), .A2 (slo__sro_n1571));
NAND2_X1 slo__sro_c2279 (.ZN (n_281), .A1 (slo__sro_n1570), .A2 (slo__sro_n1572));
XNOR2_X1 slo__sro_c2280 (.ZN (slo__sro_n1569), .A (p_15[14]), .B (p_6[14]));
XNOR2_X1 slo__sro_c2281 (.ZN (n_64), .A (n_191), .B (slo__sro_n1569));
NAND2_X1 slo__sro_c2306 (.ZN (slo__sro_n1589), .A1 (n_36), .A2 (n_32));
OAI21_X1 slo__sro_c2307 (.ZN (slo__sro_n1588), .A (n_149), .B1 (n_36), .B2 (n_32));
NAND2_X1 slo__sro_c2308 (.ZN (n_39), .A1 (slo__sro_n1588), .A2 (slo__sro_n1589));
XNOR2_X1 slo__sro_c2309 (.ZN (slo__sro_n1587), .A (n_149), .B (n_32));
XNOR2_X1 slo__sro_c2310 (.ZN (n_185), .A (slo__sro_n1587), .B (n_36));
OAI21_X1 slo__sro_c2319 (.ZN (slo__sro_n1594), .A (n_142), .B1 (n_34), .B2 (n_147));
NAND2_X1 slo__sro_c2320 (.ZN (n_37), .A1 (slo__sro_n1595), .A2 (slo__sro_n1594));
XNOR2_X1 slo__sro_c2321 (.ZN (slo__sro_n1593), .A (n_34), .B (n_147));
XNOR2_X1 slo__sro_c2322 (.ZN (n_36), .A (slo__sro_n1593), .B (n_142));
AOI22_X1 slo__sro_c2331 (.ZN (slo__sro_n1600), .A1 (p_0[10]), .A2 (p_2[10]), .B1 (p_1[10]), .B2 (p_2[10]));
NAND2_X1 slo__sro_c2332 (.ZN (n_142), .A1 (slo__sro_n1601), .A2 (slo__sro_n1600));
XNOR2_X1 slo__sro_c2333 (.ZN (slo__sro_n1599), .A (p_2[10]), .B (p_1[10]));
XNOR2_X1 slo__sro_c2334 (.ZN (n_24), .A (slo__sro_n1599), .B (p_0[10]));
OAI21_X1 slo__sro_c2343 (.ZN (slo__sro_n1606), .A (n_631), .B1 (n_646), .B2 (n_648));
NAND2_X1 slo__sro_c2344 (.ZN (n_1043), .A1 (slo__sro_n1606), .A2 (slo__sro_n1607));
XNOR2_X1 slo__sro_c2345 (.ZN (slo__sro_n1605), .A (n_631), .B (n_648));
XNOR2_X2 slo__sro_c2346 (.ZN (n_652), .A (slo__sro_n1605), .B (n_646));
NAND2_X1 slo__sro_c2355 (.ZN (slo__sro_n1614), .A1 (n_599), .A2 (n_601));
NOR2_X1 slo__sro_c2356 (.ZN (slo__sro_n1613), .A1 (n_599), .A2 (n_601));
OAI21_X1 slo__sro_c2357 (.ZN (slo__sro_n1612), .A (slo__sro_n1614), .B1 (slo__sro_n1615), .B2 (slo__sro_n1613));
XNOR2_X1 slo__sro_c2358 (.ZN (slo__sro_n1611), .A (n_599), .B (n_601));
XNOR2_X1 slo__sro_c2359 (.ZN (n_624), .A (slo__sro_n1611), .B (n_597));
AOI22_X1 slo__sro_c2369 (.ZN (slo__sro_n1623), .A1 (n_652), .A2 (n_633), .B1 (n_633), .B2 (n_650));
NAND2_X1 slo__sro_c2370 (.ZN (slo__sro_n1622), .A1 (slo__sro_n1623), .A2 (slo__sro_n1624));
XNOR2_X1 slo__sro_c2371 (.ZN (slo__sro_n1621), .A (n_650), .B (n_633));
XNOR2_X2 slo__sro_c2372 (.ZN (n_654), .A (slo__sro_n1621), .B (n_652));
INV_X2 slo__c2386 (.ZN (n_1058), .A (slo__n1633));
OAI21_X1 slo__sro_c2408 (.ZN (slo__sro_n1645), .A (n_491), .B1 (n_514), .B2 (n_487));
NAND2_X1 slo__sro_c2409 (.ZN (n_921), .A1 (slo__sro_n1645), .A2 (slo__sro_n1646));
XNOR2_X1 slo__sro_c2410 (.ZN (slo__sro_n1644), .A (n_491), .B (n_487));
XNOR2_X1 slo__sro_c2411 (.ZN (n_518), .A (slo__sro_n1644), .B (n_514));
INV_X1 slo__sro_c2420 (.ZN (slo__sro_n1654), .A (n_874));
NAND2_X1 slo__sro_c2421 (.ZN (slo__sro_n1653), .A1 (n_874), .A2 (n_482));
NAND2_X1 slo__sro_c2422 (.ZN (slo__sro_n1652), .A1 (slo__sro_n1654), .A2 (slo__sro_n1655));
NAND2_X1 slo__sro_c2423 (.ZN (slo__sro_n1651), .A1 (n_484), .A2 (slo__sro_n1652));
NAND2_X1 slo__sro_c2424 (.ZN (n_491), .A1 (slo__sro_n1651), .A2 (slo__sro_n1653));
XNOR2_X1 slo__sro_c2425 (.ZN (slo__sro_n1650), .A (n_874), .B (n_482));
XNOR2_X1 slo__sro_c2426 (.ZN (n_490), .A (n_484), .B (slo__sro_n1650));
NAND2_X1 slo__sro_c2438 (.ZN (slo__sro_n1664), .A1 (n_909), .A2 (n_871));
NOR2_X1 slo__sro_c2439 (.ZN (slo__sro_n1663), .A1 (n_871), .A2 (n_909));
OAI21_X1 slo__sro_c2440 (.ZN (n_485), .A (slo__sro_n1664), .B1 (slo__sro_n1665), .B2 (slo__sro_n1663));
XNOR2_X1 slo__sro_c2441 (.ZN (slo__sro_n1662), .A (n_909), .B (n_871));
XNOR2_X1 slo__sro_c2442 (.ZN (n_484), .A (slo__sro_n1662), .B (n_877));
NAND2_X1 slo__sro_c2478 (.ZN (slo__sro_n1692), .A1 (n_702), .A2 (slo__sro_n816));
OR2_X1 slo__sro_c2479 (.ZN (slo__sro_n1691), .A1 (n_702), .A2 (slo__sro_n816));
NAND2_X1 slo__sro_c2480 (.ZN (slo__sro_n1690), .A1 (slo__sro_n1691), .A2 (n_704));
NAND2_X1 slo__sro_c2481 (.ZN (n_707), .A1 (slo__sro_n1690), .A2 (slo__sro_n1692));
XNOR2_X1 slo__sro_c2482 (.ZN (slo__sro_n1689), .A (n_702), .B (slo__sro_n816));
XNOR2_X1 slo__sro_c2483 (.ZN (slo__sro_n1688), .A (n_704), .B (slo__sro_n1689));
INV_X1 slo__sro_c2493 (.ZN (slo__sro_n1704), .A (n_746));
NAND2_X1 slo__sro_c2494 (.ZN (slo__sro_n1703), .A1 (n_746), .A2 (n_1178));
NAND2_X1 slo__sro_c2495 (.ZN (slo__sro_n1702), .A1 (slo__sro_n1704), .A2 (slo__sro_n1705));
NAND2_X1 slo__sro_c2496 (.ZN (slo__sro_n1701), .A1 (slo__sro_n1702), .A2 (slo__sro_n1714));
NAND2_X1 slo__sro_c2497 (.ZN (n_751), .A1 (slo__sro_n1701), .A2 (slo__sro_n1703));
XNOR2_X2 slo__sro_c2498 (.ZN (slo__sro_n1700), .A (n_746), .B (n_1178));
XNOR2_X1 slo__sro_c2499 (.ZN (n_750), .A (slo__sro_n1714), .B (slo__sro_n1700));
INV_X1 slo__sro_c2513 (.ZN (slo__sro_n1718), .A (n_1181));
NAND2_X1 slo__sro_c2514 (.ZN (slo__sro_n1717), .A1 (n_744), .A2 (n_868));
NOR2_X1 slo__sro_c2515 (.ZN (slo__sro_n1716), .A1 (n_744), .A2 (n_868));
OAI21_X1 slo__sro_c2516 (.ZN (n_749), .A (slo__sro_n1717), .B1 (slo__sro_n1716), .B2 (slo__sro_n1718));
XNOR2_X1 slo__sro_c2517 (.ZN (slo__sro_n1715), .A (n_744), .B (n_868));
XNOR2_X1 slo__sro_c2518 (.ZN (slo__sro_n1714), .A (slo__sro_n1715), .B (n_1181));
INV_X1 slo__sro_c2539 (.ZN (slo__sro_n1736), .A (n_206));
NAND2_X1 slo__sro_c2540 (.ZN (slo__sro_n1735), .A1 (n_463), .A2 (n_206));
NAND2_X1 slo__sro_c2541 (.ZN (slo__sro_n1734), .A1 (slo__sro_n1737), .A2 (slo__sro_n1736));
NAND2_X1 slo__sro_c2542 (.ZN (slo__sro_n1733), .A1 (n_472), .A2 (slo__sro_n1734));
NAND2_X1 slo__sro_c2543 (.ZN (n_211), .A1 (slo__sro_n1735), .A2 (slo__sro_n1733));
XNOR2_X1 slo__sro_c2544 (.ZN (slo__sro_n1732), .A (n_463), .B (n_206));
XNOR2_X1 slo__sro_c2545 (.ZN (n_210), .A (n_472), .B (slo__sro_n1732));
OAI21_X1 slo__sro_c2559 (.ZN (slo__sro_n1748), .A (n_588), .B1 (n_308), .B2 (n_306));
NAND2_X1 slo__sro_c2560 (.ZN (slo__sro_n1747), .A1 (slo__sro_n1748), .A2 (slo__sro_n1749));
XNOR2_X2 slo__sro_c2561 (.ZN (slo__sro_n1746), .A (n_588), .B (n_306));
XNOR2_X2 slo__sro_c2562 (.ZN (n_665), .A (slo__sro_n1746), .B (n_308));
INV_X1 slo__sro_c2573 (.ZN (slo__sro_n1761), .A (n_154));
NAND2_X1 slo__sro_c2574 (.ZN (slo__sro_n1760), .A1 (n_154), .A2 (n_139));
NAND2_X1 slo__sro_c2575 (.ZN (slo__sro_n1759), .A1 (slo__sro_n1761), .A2 (slo__sro_n1762));
NAND2_X2 slo__sro_c2576 (.ZN (slo__sro_n1758), .A1 (n_141), .A2 (slo__sro_n1759));
NAND2_X2 slo__sro_c2577 (.ZN (n_445), .A1 (slo__sro_n1760), .A2 (slo__sro_n1758));
XNOR2_X1 slo__sro_c2578 (.ZN (slo__sro_n1757), .A (n_154), .B (n_139));
XNOR2_X1 slo__sro_c2579 (.ZN (slo__sro_n1756), .A (n_141), .B (slo__sro_n1757));
NAND2_X1 slo__sro_c2602 (.ZN (slo__sro_n1780), .A1 (n_113), .A2 (n_132));
NOR2_X1 slo__sro_c2603 (.ZN (slo__sro_n1779), .A1 (n_113), .A2 (n_132));
OAI21_X1 slo__sro_c2604 (.ZN (n_137), .A (slo__sro_n1780), .B1 (slo__sro_n1781), .B2 (slo__sro_n1779));
XNOR2_X1 slo__sro_c2605 (.ZN (slo__sro_n1778), .A (n_113), .B (n_132));
XNOR2_X1 slo__sro_c2606 (.ZN (n_136), .A (slo__sro_n1778), .B (n_119));
INV_X1 slo__sro_c2634 (.ZN (slo__sro_n1804), .A (n_233));
NAND2_X1 slo__sro_c2635 (.ZN (slo__sro_n1803), .A1 (n_250), .A2 (n_233));
NAND2_X1 slo__sro_c2636 (.ZN (slo__sro_n1802), .A1 (slo__sro_n1805), .A2 (slo__sro_n1804));
NAND2_X1 slo__sro_c2637 (.ZN (slo__sro_n1801), .A1 (n_235), .A2 (slo__sro_n1802));
NAND2_X1 slo__sro_c2638 (.ZN (slo__sro_n1800), .A1 (slo__sro_n1801), .A2 (slo__sro_n1803));
XNOR2_X1 slo__sro_c2639 (.ZN (slo__sro_n1799), .A (n_250), .B (n_233));
XNOR2_X1 slo__sro_c2640 (.ZN (slo__sro_n1798), .A (n_235), .B (slo__sro_n1799));
NAND2_X1 slo__sro_c2652 (.ZN (slo__sro_n1820), .A1 (n_201), .A2 (n_203));
NOR2_X1 slo__sro_c2653 (.ZN (slo__sro_n1819), .A1 (n_201), .A2 (n_203));
OAI21_X1 slo__sro_c2654 (.ZN (slo__sro_n1818), .A (slo__sro_n1820), .B1 (slo__sro_n1821), .B2 (slo__sro_n1819));
XNOR2_X1 slo__sro_c2655 (.ZN (slo__sro_n1817), .A (n_201), .B (n_203));
XNOR2_X1 slo__sro_c2656 (.ZN (slo__sro_n1816), .A (slo__sro_n1817), .B (n_209));
INV_X1 slo__sro_c2666 (.ZN (slo__sro_n1834), .A (n_228));
NAND2_X1 slo__sro_c2667 (.ZN (slo__sro_n1833), .A1 (n_220), .A2 (n_228));
NAND2_X1 slo__sro_c2668 (.ZN (slo__sro_n1832), .A1 (slo__sro_n1834), .A2 (slo__sro_n1835));
NAND2_X1 slo__sro_c2669 (.ZN (slo__sro_n1831), .A1 (slo__sro_n1832), .A2 (slo__sro_n1816));
NAND2_X1 slo__sro_c2670 (.ZN (n_235), .A1 (slo__sro_n1831), .A2 (slo__sro_n1833));
XNOR2_X1 slo__sro_c2671 (.ZN (slo__sro_n1830), .A (n_228), .B (n_220));
XNOR2_X1 slo__sro_c2672 (.ZN (n_234), .A (slo__sro_n1816), .B (slo__sro_n1830));
INV_X1 slo__sro_c2696 (.ZN (slo__sro_n1858), .A (n_770));
NAND2_X1 slo__sro_c2697 (.ZN (slo__sro_n1857), .A1 (n_770), .A2 (n_761));
NAND2_X1 slo__sro_c2698 (.ZN (slo__sro_n1856), .A1 (slo__sro_n1859), .A2 (slo__sro_n1858));
NAND2_X1 slo__sro_c2699 (.ZN (slo__sro_n1855), .A1 (slo__sro_n1856), .A2 (slo__sro_n1868));
NAND2_X1 slo__sro_c2700 (.ZN (n_1205), .A1 (slo__sro_n1855), .A2 (slo__sro_n1857));
XNOR2_X2 slo__sro_c2701 (.ZN (slo__sro_n1854), .A (n_770), .B (n_761));
XNOR2_X2 slo__sro_c2702 (.ZN (n_774), .A (slo__sro_n1868), .B (slo__sro_n1854));
NAND2_X1 slo__sro_c2719 (.ZN (slo__sro_n1872), .A1 (n_863), .A2 (n_766));
NOR2_X1 slo__sro_c2720 (.ZN (slo__sro_n1871), .A1 (n_863), .A2 (n_766));
OAI21_X1 slo__sro_c2721 (.ZN (slo__sro_n1870), .A (slo__sro_n1872), .B1 (slo__sro_n1873), .B2 (slo__sro_n1871));
XNOR2_X1 slo__sro_c2722 (.ZN (slo__sro_n1869), .A (n_766), .B (n_863));
XNOR2_X1 slo__sro_c2723 (.ZN (slo__sro_n1868), .A (n_759), .B (slo__sro_n1869));
INV_X1 CLOCK_sgo__sro_c3574 (.ZN (CLOCK_sgo__sro_n2645), .A (n_593));
AND2_X1 CLOCK_sgo__sro_c3575 (.ZN (n_1070), .A1 (slo__sro_n1339), .A2 (n_593));
INV_X4 opt_ipo_c2755 (.ZN (opt_ipo_n1905), .A (sgo__n166));
INV_X2 CLOCK_sgo__c3792 (.ZN (sgo__sro_n191), .A (CLOCK_sgo__n2761));
INV_X1 CLOCK_sgo__sro_c3684 (.ZN (CLOCK_sgo__sro_n2706), .A (opt_ipo_n1924));
NAND3_X2 CLOCK_sgo__c3551 (.ZN (CLOCK_sgo__n2632), .A1 (sgo__sro_n309), .A2 (n_739), .A3 (n_767));
INV_X4 CLOCK_sgo__c3553 (.ZN (slo__n638), .A (CLOCK_sgo__n2632));
OAI21_X4 CLOCK_sgo__sro_c3687 (.ZN (sgo__sro_n84), .A (CLOCK_sgo__sro_n2704), .B1 (CLOCK_sgo__sro_n2583), .B2 (n_833));
INV_X1 CLOCK_slo__mro_c3861 (.ZN (CLOCK_slo__mro_n2819), .A (n_1059));
BUF_X4 opt_ipo_c2774 (.Z (opt_ipo_n1924), .A (n_693));
XNOR2_X2 CLOCK_slo__mro_c3862 (.ZN (\aggregated_res[14] [40] ), .A (n_1362), .B (CLOCK_slo__mro_n2819));
OAI21_X2 CLOCK_slo__mro_c3868 (.ZN (CLOCK_slo__mro_n2828), .A (n_739), .B1 (n_959), .B2 (n_1131));
XNOR2_X2 CLOCK_slo__mro_c3869 (.ZN (\aggregated_res[14] [29] ), .A (CLOCK_slo__mro_n2828), .B (CLOCK_slo__mro_n2829));
OR2_X4 CLOCK_slo__xsl_c3910 (.ZN (n_525), .A1 (n_379), .A2 (n_409));
NAND2_X1 CLOCK_slo__sro_c3952 (.ZN (CLOCK_slo__sro_n2896), .A1 (CLOCK_slo__sro_n2898), .A2 (CLOCK_slo__sro_n2897));
NAND2_X2 CLOCK_slo__sro_c3953 (.ZN (CLOCK_slo__sro_n2895), .A1 (slo__sro_n1253), .A2 (CLOCK_slo__sro_n2896));
INV_X4 opt_ipo_c2790 (.ZN (opt_ipo_n1940), .A (n_529));
BUF_X4 opt_ipo_c3184 (.Z (opt_ipo_n2336), .A (n_30));
INV_X2 opt_ipo_c3186 (.ZN (opt_ipo_n2338), .A (n_641));
INV_X4 opt_ipo_c2798 (.ZN (opt_ipo_n1948), .A (n_385));
BUF_X4 spw__c4560 (.Z (n_501), .A (spw__n3514));
INV_X2 opt_ipo_c2815 (.ZN (opt_ipo_n1965), .A (sgo__n199));
INV_X4 opt_ipo_c2817 (.ZN (opt_ipo_n1967), .A (sgo__n168));
INV_X4 opt_ipo_c2871 (.ZN (opt_ipo_n2021), .A (sgo__sro_n84));
INV_X1 opt_ipo_c2941 (.ZN (opt_ipo_n2091), .A (sgo__n107));
INV_X1 opt_ipo_c2966 (.ZN (opt_ipo_n2116), .A (opt_ipo_n2117));
INV_X2 opt_ipo_c2967 (.ZN (opt_ipo_n2117), .A (n_614));
BUF_X2 opt_ipo_c3000 (.Z (opt_ipo_n2150), .A (n_70));
INV_X1 opt_ipo_c3002 (.ZN (opt_ipo_n2152), .A (opt_ipo_n2153));
INV_X1 opt_ipo_c3003 (.ZN (opt_ipo_n2153), .A (opt_ipo_n2154));
INV_X2 opt_ipo_c3004 (.ZN (opt_ipo_n2154), .A (n_733));
CLKBUF_X1 CLOCK_spw__L1_c4066 (.Z (CLOCK_spw__n3015), .A (n_455));
INV_X4 opt_ipo_c3018 (.ZN (opt_ipo_n2168), .A (sgo__n115));

endmodule //datapath__0_67

module datapath__0_1 (B_in, p_0);

output [31:0] p_0;
input [31:0] B_in;
wire slo__sro_n738;
wire n_3;
wire n_37;
wire n_2;
wire n_13;
wire n_15;
wire n_26;
wire slo__xsl_n137;
wire n_14;
wire n_11;
wire n_25;
wire n_9;
wire n_10;
wire n_24;
wire n_8;
wire n_66;
wire n_19;
wire n_39;
wire n_41;
wire n_23;
wire n_51;
wire n_21;
wire n_22;
wire n_55;
wire n_20;
wire n_61;
wire n_56;
wire n_78;
wire n_63;
wire n_69;
wire n_70;
wire n_47;
wire n_48;
wire n_50;
wire n_76;
wire n_49;
wire n_75;
wire n_79;
wire n_71;
wire n_1;
wire n_4;
wire n_5;
wire n_6;
wire slo__n495;
wire n_12;
wire n_16;
wire n_17;
wire n_18;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_36;
wire n_34;
wire n_35;
wire n_38;
wire n_42;
wire n_43;
wire n_44;
wire n_53;
wire n_46;
wire n_52;
wire n_57;
wire n_54;
wire n_58;
wire n_59;
wire n_60;
wire n_65;
wire n_64;
wire n_67;
wire n_68;
wire n_72;
wire n_73;
wire n_74;
wire n_77;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire sgo__n14;
wire slo__xsl_n50;
wire slo__n253;
wire slo__n364;
wire slo__sro_n739;
wire CLOCK_sgo__sro_n1049;
wire CLOCK_sgo__sro_n1048;
wire CLOCK_sgo__sro_n1050;


XOR2_X1 i_114 (.Z (p_0[31]), .A (n_81), .B (B_in[31]));
AOI21_X1 i_113 (.ZN (p_0[30]), .A (n_82), .B1 (n_83), .B2 (B_in[30]));
NAND4_X1 i_112 (.ZN (n_83), .A1 (n_79), .A2 (n_63), .A3 (n_76), .A4 (n_71));
INV_X1 i_111 (.ZN (n_82), .A (n_81));
NAND4_X2 i_110 (.ZN (n_81), .A1 (n_78), .A2 (n_80), .A3 (n_79), .A4 (n_76));
INV_X1 i_109 (.ZN (n_80), .A (B_in[30]));
NOR2_X1 i_108 (.ZN (n_79), .A1 (B_in[29]), .A2 (B_in[28]));
INV_X2 i_107 (.ZN (n_78), .A (n_70));
INV_X1 i_106 (.ZN (n_77), .A (n_73));
NOR2_X1 i_105 (.ZN (n_76), .A1 (n_74), .A2 (B_in[27]));
NOR3_X1 i_104 (.ZN (n_75), .A1 (n_70), .A2 (B_in[27]), .A3 (n_74));
AOI21_X1 i_103 (.ZN (p_0[27]), .A (n_75), .B1 (n_77), .B2 (B_in[27]));
OR3_X1 i_102 (.ZN (n_74), .A1 (B_in[26]), .A2 (B_in[24]), .A3 (B_in[25]));
NOR2_X1 i_101 (.ZN (n_73), .A1 (n_70), .A2 (n_74));
AOI21_X1 i_100 (.ZN (p_0[26]), .A (n_73), .B1 (B_in[26]), .B2 (n_68));
INV_X1 i_99 (.ZN (n_72), .A (B_in[25]));
INV_X1 i_98 (.ZN (n_71), .A (B_in[23]));
NOR3_X1 CLOCK_sgo__sro_c1312 (.ZN (CLOCK_sgo__sro_n1050), .A1 (B_in[13]), .A2 (B_in[12]), .A3 (B_in[14]));
NOR2_X4 i_96 (.ZN (n_69), .A1 (n_70), .A2 (B_in[24]));
NAND2_X2 i_95 (.ZN (n_68), .A1 (n_72), .A2 (n_69));
OAI21_X1 i_94 (.ZN (n_67), .A (n_68), .B1 (n_72), .B2 (n_69));
INV_X1 i_93 (.ZN (p_0[25]), .A (n_67));
INV_X2 i_92 (.ZN (n_66), .A (n_33));
INV_X1 i_91 (.ZN (n_65), .A (n_59));
NOR3_X1 i_90 (.ZN (n_64), .A1 (B_in[22]), .A2 (B_in[20]), .A3 (B_in[21]));
NOR2_X1 slo__c462 (.ZN (slo__n364), .A1 (n_41), .A2 (B_in[13]));
AOI21_X1 i_87 (.ZN (p_0[22]), .A (n_63), .B1 (B_in[22]), .B2 (n_65));
NOR2_X2 i_86 (.ZN (n_61), .A1 (n_56), .A2 (B_in[20]));
INV_X2 i_85 (.ZN (n_60), .A (n_61));
NOR2_X4 i_84 (.ZN (n_59), .A1 (n_60), .A2 (B_in[21]));
OR3_X2 i_82 (.ZN (n_58), .A1 (B_in[17]), .A2 (B_in[16]), .A3 (B_in[18]));
NOR2_X2 i_81 (.ZN (n_57), .A1 (B_in[19]), .A2 (n_58));
NAND2_X2 i_80 (.ZN (n_56), .A1 (n_46), .A2 (n_57));
NOR2_X1 i_79 (.ZN (n_55), .A1 (n_51), .A2 (n_58));
INV_X1 i_78 (.ZN (n_54), .A (n_55));
AOI22_X1 i_77 (.ZN (p_0[19]), .A1 (n_46), .A2 (n_57), .B1 (n_54), .B2 (B_in[19]));
INV_X1 i_76 (.ZN (n_53), .A (B_in[15]));
AND4_X2 i_75 (.ZN (n_52), .A1 (n_43), .A2 (n_42), .A3 (n_53), .A4 (n_44));
NAND4_X4 i_74 (.ZN (n_51), .A1 (n_37), .A2 (n_36), .A3 (n_34), .A4 (n_52));
INV_X2 i_73 (.ZN (n_46), .A (n_51));
OAI21_X1 i_72 (.ZN (p_0[15]), .A (n_51), .B1 (CLOCK_sgo__sro_n1048), .B2 (n_53));
INV_X1 i_70 (.ZN (n_44), .A (B_in[14]));
INV_X1 i_69 (.ZN (n_43), .A (B_in[13]));
INV_X1 i_68 (.ZN (n_42), .A (B_in[12]));
INV_X2 i_67 (.ZN (n_41), .A (n_32));
NOR2_X1 i_65 (.ZN (n_39), .A1 (n_41), .A2 (B_in[13]));
INV_X1 i_64 (.ZN (n_38), .A (slo__n364));
AOI21_X2 i_63 (.ZN (p_0[14]), .A (CLOCK_sgo__sro_n1048), .B1 (B_in[14]), .B2 (n_38));
INV_X4 i_62 (.ZN (n_37), .A (slo__n253));
INV_X2 i_61 (.ZN (n_36), .A (n_27));
INV_X1 i_60 (.ZN (n_35), .A (B_in[11]));
AND4_X2 i_59 (.ZN (n_34), .A1 (n_30), .A2 (n_29), .A3 (n_35), .A4 (n_31));
NAND3_X4 i_58 (.ZN (n_33), .A1 (n_37), .A2 (n_36), .A3 (n_34));
NOR2_X4 i_57 (.ZN (n_32), .A1 (n_33), .A2 (B_in[12]));
AOI21_X1 i_56 (.ZN (p_0[12]), .A (n_32), .B1 (B_in[12]), .B2 (n_33));
INV_X1 i_55 (.ZN (n_31), .A (B_in[10]));
INV_X1 i_54 (.ZN (n_30), .A (B_in[9]));
INV_X1 i_53 (.ZN (n_29), .A (B_in[8]));
INV_X1 i_52 (.ZN (n_28), .A (B_in[7]));
NAND4_X2 i_51 (.ZN (n_27), .A1 (n_17), .A2 (n_16), .A3 (n_28), .A4 (n_18));
NOR2_X1 i_50 (.ZN (n_26), .A1 (n_6), .A2 (n_27));
INV_X2 i_49 (.ZN (n_25), .A (slo__n495));
NOR4_X4 i_48 (.ZN (n_24), .A1 (n_25), .A2 (B_in[9]), .A3 (B_in[8]), .A4 (B_in[10]));
INV_X1 i_47 (.ZN (n_19), .A (n_24));
INV_X1 i_46 (.ZN (n_18), .A (B_in[6]));
INV_X1 i_45 (.ZN (n_17), .A (B_in[5]));
INV_X1 i_44 (.ZN (n_16), .A (B_in[4]));
INV_X1 i_42 (.ZN (n_15), .A (n_5));
NOR2_X2 i_40 (.ZN (n_13), .A1 (B_in[5]), .A2 (n_15));
INV_X1 i_39 (.ZN (n_12), .A (n_13));
AOI21_X1 i_38 (.ZN (p_0[6]), .A (slo__xsl_n50), .B1 (B_in[6]), .B2 (n_12));
AND2_X1 slo__sro_c945 (.ZN (slo__sro_n739), .A1 (n_64), .A2 (n_71));
INV_X1 slo__xsl_c199 (.ZN (slo__xsl_n137), .A (n_63));
NOR2_X1 i_35 (.ZN (n_5), .A1 (B_in[4]), .A2 (slo__n253));
AOI21_X1 i_32 (.ZN (p_0[4]), .A (n_5), .B1 (B_in[4]), .B2 (n_6));
INV_X1 i_31 (.ZN (n_4), .A (B_in[2]));
NOR2_X1 i_30 (.ZN (n_3), .A1 (B_in[0]), .A2 (B_in[1]));
NAND2_X1 i_29 (.ZN (n_2), .A1 (n_4), .A2 (n_3));
OAI21_X1 i_28 (.ZN (n_1), .A (n_2), .B1 (n_4), .B2 (n_3));
INV_X1 i_27 (.ZN (p_0[2]), .A (n_1));
INV_X1 i_26 (.ZN (n_50), .A (B_in[28]));
NAND4_X2 i_25 (.ZN (n_49), .A1 (n_63), .A2 (n_50), .A3 (n_71), .A4 (n_76));
AOI22_X2 i_23 (.ZN (p_0[29]), .A1 (n_49), .A2 (B_in[29]), .B1 (n_75), .B2 (n_79));
INV_X1 i_22 (.ZN (n_48), .A (n_49));
AOI21_X1 i_21 (.ZN (n_47), .A (n_50), .B1 (n_78), .B2 (n_76));
NOR2_X1 i_20 (.ZN (p_0[28]), .A1 (n_47), .A2 (n_48));
AOI21_X1 i_19 (.ZN (p_0[24]), .A (n_69), .B1 (B_in[24]), .B2 (n_70));
AOI21_X1 i_18 (.ZN (p_0[23]), .A (n_78), .B1 (B_in[23]), .B2 (slo__xsl_n137));
AOI21_X1 i_43 (.ZN (p_0[20]), .A (n_61), .B1 (B_in[20]), .B2 (n_56));
NOR2_X2 i_17 (.ZN (n_23), .A1 (n_51), .A2 (B_in[16]));
INV_X2 i_16 (.ZN (n_22), .A (n_23));
NOR2_X4 i_15 (.ZN (n_21), .A1 (n_22), .A2 (B_in[17]));
INV_X1 i_14 (.ZN (n_20), .A (n_21));
AOI21_X1 i_13 (.ZN (p_0[18]), .A (n_55), .B1 (B_in[18]), .B2 (n_20));
AOI21_X1 i_34 (.ZN (p_0[17]), .A (n_21), .B1 (B_in[17]), .B2 (n_22));
AOI21_X1 i_33 (.ZN (p_0[16]), .A (n_23), .B1 (B_in[16]), .B2 (n_51));
AOI21_X1 i_24 (.ZN (p_0[13]), .A (n_39), .B1 (n_41), .B2 (B_in[13]));
NOR2_X2 i_12 (.ZN (n_11), .A1 (n_25), .A2 (B_in[8]));
INV_X2 i_11 (.ZN (n_10), .A (n_11));
NOR2_X4 i_10 (.ZN (n_9), .A1 (n_10), .A2 (B_in[9]));
INV_X1 i_9 (.ZN (n_8), .A (n_9));
AOI21_X1 i_8 (.ZN (p_0[11]), .A (n_66), .B1 (n_19), .B2 (B_in[11]));
AOI21_X1 i_7 (.ZN (p_0[10]), .A (n_24), .B1 (n_8), .B2 (B_in[10]));
AOI21_X1 i_5 (.ZN (p_0[8]), .A (n_11), .B1 (B_in[8]), .B2 (n_25));
AOI21_X2 i_3 (.ZN (p_0[7]), .A (n_26), .B1 (n_14), .B2 (B_in[7]));
AOI21_X1 i_2 (.ZN (p_0[5]), .A (n_13), .B1 (B_in[5]), .B2 (n_15));
AOI21_X1 i_1 (.ZN (p_0[3]), .A (n_37), .B1 (B_in[3]), .B2 (n_2));
AOI21_X1 i_0 (.ZN (p_0[1]), .A (n_3), .B1 (B_in[1]), .B2 (B_in[0]));
NOR2_X2 slo__c634 (.ZN (slo__n495), .A1 (n_6), .A2 (n_27));
NOR4_X4 sgo__c13 (.ZN (sgo__n14), .A1 (B_in[0]), .A2 (B_in[2]), .A3 (B_in[3]), .A4 (B_in[1]));
INV_X1 sgo__c15 (.ZN (n_6), .A (sgo__n14));
INV_X1 slo__xsl_c63 (.ZN (slo__xsl_n50), .A (n_14));
OR4_X2 slo__xsl_c66 (.ZN (n_14), .A1 (n_6), .A2 (B_in[5]), .A3 (B_in[4]), .A4 (B_in[6]));
AND4_X4 slo__xsl_c202 (.ZN (n_63), .A1 (n_66), .A2 (n_57), .A3 (n_52), .A4 (n_64));
INV_X2 slo__c334 (.ZN (slo__n253), .A (sgo__n14));
AOI21_X1 slo__sro_c715 (.ZN (p_0[21]), .A (n_59), .B1 (n_60), .B2 (B_in[21]));
AOI21_X1 slo__sro_c673 (.ZN (p_0[9]), .A (n_9), .B1 (n_10), .B2 (B_in[9]));
NAND2_X4 slo__sro_c947 (.ZN (n_70), .A1 (n_46), .A2 (slo__sro_n738));
AND2_X1 slo__sro_c946 (.ZN (slo__sro_n738), .A1 (n_57), .A2 (slo__sro_n739));
NOR2_X1 CLOCK_sgo__sro_c1314 (.ZN (CLOCK_sgo__sro_n1048), .A1 (n_33), .A2 (CLOCK_sgo__sro_n1049));
INV_X1 CLOCK_sgo__sro_c1313 (.ZN (CLOCK_sgo__sro_n1049), .A (CLOCK_sgo__sro_n1050));

endmodule //datapath__0_1

module datapath__0_0 (opt_ipoPP_2, opt_ipoPP_3, opt_ipoPP_6, opt_ipoPP_7, opt_ipoPP_8, 
    opt_ipoPP_12, opt_ipoPP_13, opt_ipoPP_14, opt_ipoPP_15, opt_ipoPP_17, opt_ipoPP_20, 
    opt_ipoPP_21, opt_ipoPP_22, A_imm, A_imm_2s_complement);

output [31:0] A_imm_2s_complement;
input [31:0] A_imm;
input opt_ipoPP_2;
input opt_ipoPP_3;
input opt_ipoPP_6;
input opt_ipoPP_7;
input opt_ipoPP_8;
input opt_ipoPP_12;
input opt_ipoPP_13;
input opt_ipoPP_14;
input opt_ipoPP_15;
input opt_ipoPP_17;
input opt_ipoPP_20;
input opt_ipoPP_21;
input opt_ipoPP_22;
wire drc_ipo_n39;
wire slo__mro_n456;
wire slo__n890;
wire slo__n1070;
wire slo__n809;
wire opt_ipo_n1512;
wire opt_ipo_n1634;
wire drc_ipo_n41;
wire n_19;
wire n_13;
wire n_55;
wire slo__mro_n524;
wire n_1;
wire n_23;
wire n_45;
wire n_43;
wire slo__xsl_n561;
wire slo__n554;
wire n_7;
wire n_35;
wire n_14;
wire slo__sro_n754;
wire n_8;
wire n_24;
wire n_20;
wire slo__sro_n475;
wire n_21;
wire n_22;
wire n_114;
wire n_113;
wire n_25;
wire n_26;
wire n_28;
wire n_27;
wire n_30;
wire n_29;
wire n_77;
wire n_32;
wire n_50;
wire n_49;
wire n_51;
wire n_54;
wire n_53;
wire n_56;
wire n_40;
wire n_63;
wire n_11;
wire n_65;
wire n_38;
wire n_66;
wire n_67;
wire n_68;
wire n_70;
wire n_60;
wire n_61;
wire n_37;
wire n_79;
wire n_76;
wire n_90;
wire slo__mro_n525;
wire n_85;
wire n_100;
wire n_97;
wire n_91;
wire CLOCK_sgo__sro_n1871;
wire n_6;
wire n_15;
wire n_16;
wire n_36;
wire n_41;
wire n_58;
wire n_42;
wire sgo__sro_n201;
wire n_112;
wire n_62;
wire n_64;
wire n_69;
wire n_71;
wire n_73;
wire slo__n498;
wire n_75;
wire n_81;
wire n_83;
wire n_89;
wire n_86;
wire n_84;
wire sgo__sro_n250;
wire n_88;
wire n_94;
wire n_93;
wire n_95;
wire n_96;
wire n_98;
wire n_101;
wire n_102;
wire n_103;
wire sgo__sro_n249;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_111;
wire n_110;
wire sgo__sro_n148;
wire sgo__n360;
wire sgo__sro_n168;
wire sgo__sro_n149;
wire sgo__sro_n200;
wire sgo__sro_n198;
wire sgo__sro_n199;
wire sgo__sro_n326;
wire sgo__sro_n385;
wire slo__mro_n457;
wire slo__sro_n476;
wire slo__mro_n526;
wire slo__mro_n527;
wire slo__n582;
wire CLOCK_sgo__sro_n1872;
wire slo__sro_n676;
wire slo__sro_n677;
wire opt_ipo_n1387;
wire slo__xsl_n733;
wire slo__sro_n791;
wire slo__sro_n814;
wire slo__sro_n815;
wire slo__n836;
wire slo__n900;
wire opt_ipo_n1651;
wire slo__n970;
wire slo__n977;
wire CLOCK_sgo__sro_n1859;
wire slo__n1024;
wire slo__sro_n1041;
wire slo__sro_n1056;
wire opt_ipo_n1444;
wire opt_ipo_n1481;


INV_X1 i_139 (.ZN (n_114), .A (A_imm[7]));
INV_X1 i_138 (.ZN (n_113), .A (A_imm[6]));
NOR3_X4 i_137 (.ZN (n_112), .A1 (A_imm[8]), .A2 (A_imm[6]), .A3 (A_imm[7]));
NAND2_X2 i_136 (.ZN (n_111), .A1 (n_105), .A2 (n_106));
NAND3_X1 i_135 (.ZN (n_110), .A1 (n_85), .A2 (n_101), .A3 (n_96));
NOR3_X4 i_134 (.ZN (n_109), .A1 (A_imm[31]), .A2 (n_111), .A3 (n_110));
AOI21_X4 i_133 (.ZN (A_imm_2s_complement[31]), .A (n_109), .B1 (A_imm[31]), .B2 (sgo__sro_n148));
AOI21_X4 i_132 (.ZN (A_imm_2s_complement[30]), .A (n_107), .B1 (A_imm[30]), .B2 (n_108));
NAND3_X1 i_131 (.ZN (n_108), .A1 (n_106), .A2 (n_101), .A3 (n_94));
INV_X1 i_130 (.ZN (n_107), .A (sgo__sro_n148));
INV_X1 i_129 (.ZN (n_106), .A (A_imm[29]));
INV_X1 i_128 (.ZN (n_105), .A (A_imm[30]));
NAND2_X1 slo__mro_c589 (.ZN (slo__mro_n525), .A1 (n_43), .A2 (slo__mro_n526));
NOR2_X2 i_126 (.ZN (n_103), .A1 (A_imm[30]), .A2 (A_imm[29]));
NOR2_X1 i_125 (.ZN (n_102), .A1 (n_95), .A2 (A_imm[28]));
XNOR2_X1 i_124 (.ZN (drc_ipo_n39), .A (n_102), .B (A_imm[29]));
INV_X1 i_123 (.ZN (n_101), .A (A_imm[28]));
NOR2_X4 slo__mro_c518 (.ZN (slo__mro_n457), .A1 (A_imm[15]), .A2 (A_imm[18]));
NAND3_X2 i_120 (.ZN (n_98), .A1 (A_imm[25]), .A2 (n_89), .A3 (A_imm[26]));
INV_X1 i_119 (.ZN (n_97), .A (n_98));
NOR2_X4 i_118 (.ZN (n_96), .A1 (n_98), .A2 (A_imm[27]));
NAND4_X2 i_117 (.ZN (n_95), .A1 (n_96), .A2 (n_71), .A3 (sgo__sro_n198), .A4 (n_43));
INV_X2 i_116 (.ZN (n_94), .A (n_95));
NAND2_X1 i_115 (.ZN (n_93), .A1 (n_85), .A2 (n_97));
AOI21_X4 i_114 (.ZN (A_imm_2s_complement[27]), .A (n_94), .B1 (A_imm[27]), .B2 (n_93));
AND2_X1 i_112 (.ZN (n_91), .A1 (opt_ipoPP_15), .A2 (n_89));
NAND2_X4 slo__c922 (.ZN (slo__n890), .A1 (slo__n977), .A2 (n_71));
INV_X2 i_110 (.ZN (n_89), .A (A_imm[24]));
NAND2_X4 i_109 (.ZN (n_88), .A1 (A_imm[19]), .A2 (A_imm[20]));
AND2_X1 sgo__sro_c227 (.ZN (sgo__sro_n249), .A1 (sgo__sro_n198), .A2 (sgo__sro_n250));
CLKBUF_X1 slo__c567 (.Z (slo__n498), .A (A_imm[22]));
INV_X8 i_106 (.ZN (n_85), .A (slo__n890));
NAND2_X1 i_105 (.ZN (n_84), .A1 (n_89), .A2 (n_85));
AOI22_X4 i_104 (.ZN (A_imm_2s_complement[24]), .A1 (n_89), .A2 (n_85), .B1 (n_86), .B2 (A_imm[24]));
NOR2_X1 i_103 (.ZN (n_83), .A1 (A_imm[22]), .A2 (A_imm[21]));
NOR2_X1 i_101 (.ZN (n_81), .A1 (A_imm[21]), .A2 (opt_ipoPP_7));
INV_X1 slo__mro_c588 (.ZN (slo__mro_n526), .A (slo__mro_n527));
INV_X4 i_99 (.ZN (n_79), .A (slo__n1070));
INV_X4 i_97 (.ZN (n_77), .A (n_69));
AOI22_X4 slo__sro_c891 (.ZN (A_imm_2s_complement[25]), .A1 (n_84), .A2 (opt_ipoPP_14)
    , .B1 (n_91), .B2 (n_85));
OAI21_X1 i_95 (.ZN (n_75), .A (opt_ipoPP_7), .B1 (opt_ipoPP_13), .B2 (n_69));
NOR2_X4 slo__c863 (.ZN (slo__n809), .A1 (n_73), .A2 (slo__mro_n456));
NAND4_X4 i_92 (.ZN (n_73), .A1 (n_64), .A2 (n_42), .A3 (n_54), .A4 (n_58));
AND2_X2 sgo__sro_c226 (.ZN (sgo__sro_n250), .A1 (n_29), .A2 (n_30));
AND2_X1 slo__sro_c544 (.ZN (slo__sro_n476), .A1 (n_81), .A2 (opt_ipo_n1481));
NAND3_X4 i_89 (.ZN (n_69), .A1 (slo__n809), .A2 (n_30), .A3 (n_29));
XNOR2_X2 i_88 (.ZN (opt_ipo_n1512), .A (n_69), .B (opt_ipo_n1481));
INV_X1 i_86 (.ZN (n_64), .A (A_imm[16]));
NAND3_X2 i_85 (.ZN (n_62), .A1 (n_43), .A2 (n_54), .A3 (n_41));
XNOR2_X2 slo__sro_c848 (.ZN (slo__sro_n791), .A (n_35), .B (n_7));
XNOR2_X2 i_82 (.ZN (drc_ipo_n41), .A (n_61), .B (A_imm[16]));
INV_X1 i_75 (.ZN (n_60), .A (A_imm[14]));
BUF_X4 drc_ipo_c24 (.Z (A_imm_2s_complement[29]), .A (drc_ipo_n39));
INV_X2 i_73 (.ZN (n_58), .A (A_imm[12]));
NAND2_X4 sgo__sro_c160 (.ZN (sgo__sro_n199), .A1 (sgo__sro_n201), .A2 (sgo__sro_n200));
NAND3_X4 sgo__sro_c110 (.ZN (n_45), .A1 (n_112), .A2 (n_11), .A3 (sgo__sro_n168));
NOR2_X4 i_67 (.ZN (n_43), .A1 (n_45), .A2 (A_imm[9]));
AND2_X4 i_66 (.ZN (n_42), .A1 (A_imm[11]), .A2 (A_imm[10]));
AND2_X2 i_65 (.ZN (n_41), .A1 (n_42), .A2 (n_58));
NAND2_X2 CLOCK_sgo__sro_c1956 (.ZN (CLOCK_sgo__sro_n1871), .A1 (n_77), .A2 (CLOCK_sgo__sro_n1872));
NAND2_X1 sgo__sro_c228 (.ZN (n_86), .A1 (sgo__sro_n249), .A2 (n_71));
NAND2_X2 i_62 (.ZN (n_38), .A1 (n_54), .A2 (n_40));
NAND3_X1 i_60 (.ZN (n_37), .A1 (n_40), .A2 (n_54), .A3 (n_60));
NOR2_X1 i_59 (.ZN (n_36), .A1 (A_imm[2]), .A2 (A_imm[3]));
AND2_X2 i_58 (.ZN (n_35), .A1 (n_15), .A2 (n_36));
NOR2_X1 i_57 (.ZN (n_19), .A1 (A_imm[2]), .A2 (n_13));
INV_X1 i_56 (.ZN (n_16), .A (n_19));
AOI21_X4 i_55 (.ZN (A_imm_2s_complement[3]), .A (n_35), .B1 (slo__n582), .B2 (n_16));
NOR2_X4 i_54 (.ZN (n_15), .A1 (A_imm[1]), .A2 (A_imm[0]));
INV_X1 i_53 (.ZN (n_13), .A (n_15));
AOI21_X4 i_52 (.ZN (A_imm_2s_complement[1]), .A (n_15), .B1 (sgo__n360), .B2 (A_imm[0]));
INV_X2 i_189 (.ZN (n_8), .A (A_imm[5]));
INV_X2 i_188 (.ZN (n_7), .A (A_imm[4]));
NAND2_X2 i_187 (.ZN (n_6), .A1 (n_8), .A2 (n_7));
INV_X2 i_186 (.ZN (n_11), .A (n_6));
BUF_X2 CLOCK_sgo__sro_c1933 (.Z (CLOCK_sgo__sro_n1859), .A (n_53));
NAND2_X1 i_51 (.ZN (n_100), .A1 (n_85), .A2 (n_91));
AOI22_X4 i_50 (.ZN (A_imm_2s_complement[26]), .A1 (n_100), .A2 (opt_ipo_n1444), .B1 (n_85), .B2 (n_97));
AOI21_X4 i_49 (.ZN (A_imm_2s_complement[23]), .A (n_85), .B1 (CLOCK_sgo__sro_n1871), .B2 (A_imm[23]));
INV_X4 i_46 (.ZN (n_90), .A (CLOCK_sgo__sro_n1871));
AOI21_X4 i_45 (.ZN (A_imm_2s_complement[22]), .A (n_90), .B1 (slo__n498), .B2 (slo__sro_n475));
NAND2_X2 slo__c1092 (.ZN (slo__n1070), .A1 (n_77), .A2 (slo__sro_n476));
AOI21_X4 i_87 (.ZN (A_imm_2s_complement[15]), .A (n_61), .B1 (opt_ipoPP_17), .B2 (n_37));
INV_X1 opt_ipo_c1633 (.ZN (opt_ipo_n1651), .A (opt_ipoPP_22));
NAND2_X1 i_81 (.ZN (n_68), .A1 (n_38), .A2 (opt_ipoPP_20));
NAND2_X2 i_80 (.ZN (n_67), .A1 (n_70), .A2 (n_68));
INV_X4 i_79 (.ZN (A_imm_2s_complement[14]), .A (n_67));
NAND2_X1 i_78 (.ZN (n_66), .A1 (slo__xsl_n561), .A2 (A_imm[13]));
NAND2_X2 i_77 (.ZN (n_65), .A1 (n_38), .A2 (n_66));
INV_X4 i_76 (.ZN (A_imm_2s_complement[13]), .A (n_65));
OR2_X1 slo__sro_c823 (.ZN (slo__sro_n754), .A1 (A_imm[14]), .A2 (A_imm[15]));
INV_X1 i_21 (.ZN (n_56), .A (slo__n970));
INV_X16 i_20 (.ZN (n_54), .A (A_imm[13]));
NOR3_X1 i_19 (.ZN (n_53), .A1 (A_imm[14]), .A2 (A_imm[16]), .A3 (A_imm[15]));
NAND3_X1 i_16 (.ZN (n_50), .A1 (n_40), .A2 (n_53), .A3 (n_54));
NAND2_X1 i_15 (.ZN (n_49), .A1 (n_50), .A2 (slo__n970));
NAND2_X2 i_14 (.ZN (A_imm_2s_complement[17]), .A1 (n_49), .A2 (n_51));
NAND2_X1 slo__mro_c587 (.ZN (slo__mro_n527), .A1 (opt_ipoPP_21), .A2 (A_imm[10]));
BUF_X4 drc_ipo_c25 (.Z (A_imm_2s_complement[16]), .A (drc_ipo_n41));
OR2_X1 i_2 (.ZN (n_32), .A1 (n_50), .A2 (slo__n970));
AOI21_X2 i_0 (.ZN (opt_ipo_n1634), .A (n_77), .B1 (n_32), .B2 (A_imm[18]));
INV_X2 i_43 (.ZN (n_30), .A (A_imm[9]));
INV_X2 i_42 (.ZN (n_29), .A (n_45));
NAND4_X1 i_41 (.ZN (n_28), .A1 (opt_ipoPP_3), .A2 (n_30), .A3 (opt_ipoPP_21), .A4 (n_29));
NAND3_X1 i_40 (.ZN (n_27), .A1 (opt_ipoPP_3), .A2 (n_30), .A3 (n_29));
NAND2_X1 i_39 (.ZN (n_26), .A1 (n_27), .A2 (opt_ipoPP_12));
NAND2_X1 i_38 (.ZN (n_25), .A1 (n_26), .A2 (n_28));
INV_X2 i_37 (.ZN (A_imm_2s_complement[11]), .A (n_25));
NAND2_X4 i_36 (.ZN (n_24), .A1 (n_63), .A2 (n_113));
INV_X1 i_35 (.ZN (n_1), .A (n_24));
NAND2_X2 i_34 (.ZN (n_23), .A1 (n_1), .A2 (n_114));
NAND2_X1 i_33 (.ZN (n_22), .A1 (n_23), .A2 (opt_ipo_n1651));
NAND2_X1 i_32 (.ZN (n_21), .A1 (n_22), .A2 (n_45));
INV_X4 i_31 (.ZN (A_imm_2s_complement[8]), .A (n_21));
NAND2_X1 i_30 (.ZN (n_20), .A1 (slo__xsl_n733), .A2 (A_imm[6]));
NAND2_X1 i_29 (.ZN (A_imm_2s_complement[6]), .A1 (n_24), .A2 (n_20));
AND2_X4 slo__sro_c1079 (.ZN (slo__sro_n1056), .A1 (n_76), .A2 (opt_ipo_n1387));
OR2_X1 i_26 (.ZN (n_14), .A1 (n_63), .A2 (slo__sro_n1041));
INV_X4 i_25 (.ZN (A_imm_2s_complement[5]), .A (n_14));
NAND2_X2 slo__sro_c855 (.ZN (A_imm_2s_complement[20]), .A1 (n_76), .A2 (n_75));
INV_X4 i_23 (.ZN (A_imm_2s_complement[4]), .A (slo__sro_n791));
CLKBUF_X1 slo__c617 (.Z (slo__n554), .A (A_imm[7]));
CLKBUF_X1 slo__c653 (.Z (slo__n582), .A (A_imm[3]));
INV_X4 i_11 (.ZN (A_imm_2s_complement[12]), .A (slo__mro_n524));
XNOR2_X2 i_10 (.ZN (A_imm_2s_complement[10]), .A (n_43), .B (opt_ipoPP_3));
XNOR2_X1 i_8 (.ZN (A_imm_2s_complement[9]), .A (n_45), .B (A_imm[9]));
INV_X2 i_3 (.ZN (n_55), .A (n_23));
NOR2_X4 sgo__sro_c161 (.ZN (sgo__sro_n198), .A1 (sgo__sro_n199), .A2 (A_imm[23]));
AOI21_X4 i_6 (.ZN (A_imm_2s_complement[7]), .A (n_55), .B1 (slo__n554), .B2 (n_24));
AOI21_X4 i_1 (.ZN (A_imm_2s_complement[2]), .A (n_19), .B1 (A_imm[2]), .B2 (n_13));
CLKBUF_X1 sgo__c369 (.Z (sgo__n360), .A (A_imm[1]));
NOR2_X4 sgo__sro_c316 (.ZN (sgo__sro_n326), .A1 (A_imm[14]), .A2 (A_imm[17]));
NAND3_X2 sgo__sro_c85 (.ZN (sgo__sro_n148), .A1 (n_103), .A2 (n_85), .A3 (sgo__sro_n149));
AND2_X1 sgo__sro_c84 (.ZN (sgo__sro_n149), .A1 (n_101), .A2 (n_96));
AND2_X1 sgo__sro_c109 (.ZN (sgo__sro_n168), .A1 (slo__n1024), .A2 (n_15));
INV_X4 sgo__sro_c158 (.ZN (sgo__sro_n201), .A (n_88));
NOR2_X4 sgo__sro_c159 (.ZN (sgo__sro_n200), .A1 (A_imm[21]), .A2 (A_imm[22]));
OR2_X1 sgo__sro_c403 (.ZN (sgo__sro_n385), .A1 (n_101), .A2 (n_95));
OAI21_X4 sgo__sro_c404 (.ZN (A_imm_2s_complement[28]), .A (sgo__sro_n385), .B1 (n_94), .B2 (A_imm[28]));
NAND2_X4 slo__mro_c519 (.ZN (slo__mro_n456), .A1 (slo__mro_n457), .A2 (sgo__sro_n326));
NOR2_X2 slo__mro_c520 (.ZN (n_71), .A1 (n_73), .A2 (slo__mro_n456));
NAND2_X1 slo__sro_c545 (.ZN (slo__sro_n475), .A1 (n_77), .A2 (slo__sro_n476));
XNOR2_X2 slo__mro_c590 (.ZN (slo__mro_n524), .A (slo__mro_n525), .B (slo__n900));
INV_X1 slo__xsl_c625 (.ZN (slo__xsl_n561), .A (n_40));
AND2_X4 slo__xsl_c628 (.ZN (n_40), .A1 (n_43), .A2 (n_41));
AND3_X2 CLOCK_sgo__sro_c1955 (.ZN (CLOCK_sgo__sro_n1872), .A1 (n_83), .A2 (opt_ipo_n1481), .A3 (opt_ipoPP_6));
NAND2_X1 slo__sro_c731 (.ZN (slo__sro_n677), .A1 (n_60), .A2 (n_54));
INV_X1 slo__sro_c732 (.ZN (slo__sro_n676), .A (slo__sro_n677));
NAND2_X1 slo__sro_c733 (.ZN (n_70), .A1 (n_40), .A2 (slo__sro_n676));
NAND4_X2 CLOCK_sgo__sro_c1934 (.ZN (n_51), .A1 (n_40), .A2 (n_56), .A3 (n_54), .A4 (CLOCK_sgo__sro_n1859));
NOR2_X4 slo__sro_c824 (.ZN (n_61), .A1 (n_62), .A2 (slo__sro_n754));
INV_X1 slo__xsl_c793 (.ZN (slo__xsl_n733), .A (n_63));
AND2_X4 slo__xsl_c796 (.ZN (n_63), .A1 (n_11), .A2 (slo__n836));
INV_X2 opt_ipo_c1472 (.ZN (opt_ipo_n1387), .A (opt_ipoPP_2));
NAND2_X1 slo__sro_c868 (.ZN (slo__sro_n815), .A1 (opt_ipoPP_6), .A2 (opt_ipo_n1481));
INV_X1 slo__sro_c869 (.ZN (slo__sro_n814), .A (slo__sro_n815));
NAND2_X4 slo__sro_c870 (.ZN (n_76), .A1 (slo__sro_n814), .A2 (n_77));
AND2_X2 slo__c888 (.ZN (slo__n836), .A1 (n_36), .A2 (n_15));
CLKBUF_X1 slo__c932 (.Z (slo__n900), .A (A_imm[12]));
BUF_X8 opt_ipo_c1620 (.Z (A_imm_2s_complement[18]), .A (opt_ipo_n1634));
CLKBUF_X1 slo__c1007 (.Z (slo__n970), .A (A_imm[17]));
AND2_X4 slo__c1014 (.ZN (slo__n977), .A1 (sgo__sro_n198), .A2 (sgo__sro_n250));
NOR2_X2 slo__c1053 (.ZN (slo__n1024), .A1 (A_imm[2]), .A2 (A_imm[3]));
AOI21_X1 slo__sro_c1070 (.ZN (slo__sro_n1041), .A (n_8), .B1 (n_35), .B2 (n_7));
NOR2_X4 slo__sro_c1080 (.ZN (A_imm_2s_complement[21]), .A1 (slo__sro_n1056), .A2 (n_79));
INV_X1 opt_ipo_c1511 (.ZN (opt_ipo_n1444), .A (opt_ipoPP_8));
BUF_X1 opt_ipo_c1532 (.Z (opt_ipo_n1481), .A (A_imm[19]));
BUF_X8 opt_ipo_c1554 (.Z (A_imm_2s_complement[19]), .A (opt_ipo_n1512));

endmodule //datapath__0_0

module datapath (opt_ipoPP_1, opt_ipoPP_13, opt_ipoPP_14, A_in, p_0);

output [31:0] p_0;
input [31:0] A_in;
input opt_ipoPP_1;
input opt_ipoPP_13;
input opt_ipoPP_14;
wire slo__n1059;
wire slo__xsl_n254;
wire n_59;
wire n_55;
wire n_0;
wire n_1;
wire n_52;
wire slo__sro_n289;
wire n_7;
wire n_17;
wire n_51;
wire n_13;
wire n_14;
wire n_49;
wire n_12;
wire n_50;
wire n_15;
wire n_23;
wire n_48;
wire n_19;
wire slo__mro_n189;
wire n_45;
wire n_18;
wire n_46;
wire n_21;
wire n_25;
wire n_44;
wire n_27;
wire n_24;
wire n_43;
wire n_26;
wire n_41;
wire n_42;
wire n_29;
wire slo__mro_n327;
wire n_32;
wire n_30;
wire n_39;
wire n_31;
wire n_47;
wire slo__sro_n397;
wire n_38;
wire slo__sro_n426;
wire n_33;
wire n_37;
wire n_35;
wire n_10;
wire n_22;
wire n_62;
wire n_66;
wire n_94;
wire n_2;
wire n_86;
wire n_3;
wire n_85;
wire n_4;
wire n_54;
wire n_5;
wire n_9;
wire n_8;
wire n_71;
wire n_70;
wire n_69;
wire n_16;
wire n_11;
wire n_28;
wire n_56;
wire n_68;
wire n_53;
wire n_60;
wire n_61;
wire n_64;
wire n_90;
wire n_88;
wire n_67;
wire n_103;
wire n_65;
wire n_96;
wire n_57;
wire sgo__sro_n157;
wire n_98;
wire n_72;
wire n_75;
wire n_76;
wire n_74;
wire n_77;
wire n_104;
wire n_84;
wire n_78;
wire n_79;
wire n_80;
wire slo__xsl_n255;
wire n_83;
wire slo__n1132;
wire n_101;
wire opt_ipo_n1391;
wire n_89;
wire n_87;
wire n_93;
wire n_91;
wire n_100;
wire n_105;
wire slo__sro_n290;
wire slo__sro_n291;
wire slo__sro_n406;
wire slo__sro_n407;
wire sgo__sro_n47;
wire sgo__sro_n48;
wire sgo__sro_n49;
wire slo__sro_n398;
wire slo__sro_n427;
wire slo__sro_n428;
wire slo__mro_n471;
wire slo__xsl_n479;
wire slo__xsl_n480;
wire slo__sro_n527;
wire slo__sro_n528;
wire slo__sro_n529;
wire slo__xsl_n686;
wire slo__xsl_n687;
wire slo__n560;
wire slo__sro_n1119;
wire slo__n753;
wire slo__n646;
wire slo__sro_n937;
wire slo__xsl_n796;
wire slo__n913;
wire slo__sro_n938;
wire slo__n611;
wire opt_ipo_n1484;


INV_X2 i_129 (.ZN (n_103), .A (A_in[10]));
INV_X2 i_128 (.ZN (n_90), .A (A_in[9]));
INV_X4 i_127 (.ZN (n_88), .A (A_in[8]));
NOR3_X1 i_126 (.ZN (n_87), .A1 (A_in[9]), .A2 (A_in[8]), .A3 (A_in[10]));
INV_X4 i_119 (.ZN (n_84), .A (A_in[1]));
INV_X2 i_116 (.ZN (n_77), .A (A_in[0]));
NAND2_X1 i_115 (.ZN (n_74), .A1 (n_84), .A2 (n_77));
AOI22_X1 i_107 (.ZN (p_0[1]), .A1 (n_77), .A2 (n_84), .B1 (A_in[1]), .B2 (A_in[0]));
INV_X1 slo__sro_c424 (.ZN (slo__sro_n291), .A (A_in[28]));
INV_X2 i_138 (.ZN (n_66), .A (A_in[12]));
INV_X4 i_137 (.ZN (n_53), .A (n_65));
INV_X4 i_136 (.ZN (n_105), .A (A_in[3]));
INV_X1 i_135 (.ZN (n_104), .A (A_in[2]));
NOR2_X1 CLOCK_slo__mro_c2341 (.ZN (n_19), .A1 (n_48), .A2 (n_46));
INV_X1 i_95 (.ZN (n_100), .A (A_in[7]));
INV_X4 i_90 (.ZN (n_98), .A (A_in[5]));
INV_X1 slo__sro_c425 (.ZN (slo__sro_n290), .A (n_38));
NAND4_X4 i_88 (.ZN (n_96), .A1 (n_83), .A2 (n_100), .A3 (A_in[6]), .A4 (n_98));
NAND3_X1 sgo__sro_c240 (.ZN (n_86), .A1 (n_101), .A2 (n_68), .A3 (sgo__sro_n157));
NAND4_X1 i_125 (.ZN (n_94), .A1 (slo__n646), .A2 (n_66), .A3 (n_53), .A4 (n_68));
NAND2_X1 i_124 (.ZN (n_93), .A1 (n_94), .A2 (n_62));
INV_X4 i_122 (.ZN (n_55), .A (slo__sro_n1119));
NAND4_X1 i_121 (.ZN (n_91), .A1 (n_55), .A2 (A_in[13]), .A3 (n_66), .A4 (n_53));
NAND2_X2 i_120 (.ZN (p_0[13]), .A1 (n_93), .A2 (n_91));
INV_X1 slo__xsl_c669 (.ZN (slo__xsl_n480), .A (slo__sro_n937));
INV_X1 i_117 (.ZN (n_7), .A (n_89));
NAND3_X4 slo__mro_c289 (.ZN (slo__mro_n189), .A1 (slo__n560), .A2 (slo__n1059), .A3 (n_105));
AOI21_X1 i_113 (.ZN (p_0[10]), .A (n_7), .B1 (n_86), .B2 (A_in[10]));
XNOR2_X2 i_112 (.ZN (p_0[8]), .A (slo__sro_n1119), .B (n_88));
NOR2_X4 i_111 (.ZN (n_52), .A1 (slo__sro_n1119), .A2 (slo__xsl_n686));
INV_X2 i_110 (.ZN (n_51), .A (n_52));
NAND2_X1 i_109 (.ZN (n_85), .A1 (n_55), .A2 (n_88));
INV_X2 i_108 (.ZN (n_57), .A (slo__n913));
NOR2_X4 i_106 (.ZN (n_1), .A1 (n_57), .A2 (n_72));
INV_X4 i_105 (.ZN (n_83), .A (A_in[4]));
INV_X1 slo__xsl_c377 (.ZN (slo__xsl_n255), .A (n_42));
NOR2_X1 slo__c1408 (.ZN (slo__n1132), .A1 (n_44), .A2 (A_in[20]));
AOI21_X2 i_102 (.ZN (p_0[6]), .A (n_1), .B1 (slo__xsl_n479), .B2 (opt_ipoPP_13));
INV_X1 i_101 (.ZN (n_80), .A (slo__sro_n937));
AOI21_X1 i_100 (.ZN (n_79), .A (n_98), .B1 (slo__n646), .B2 (n_83));
NOR2_X1 i_99 (.ZN (p_0[5]), .A1 (n_80), .A2 (n_79));
XNOR2_X1 i_98 (.ZN (n_78), .A (n_57), .B (A_in[4]));
INV_X1 i_97 (.ZN (p_0[4]), .A (n_78));
NAND3_X1 i_96 (.ZN (n_59), .A1 (n_77), .A2 (n_104), .A3 (n_84));
NAND2_X1 i_94 (.ZN (n_76), .A1 (n_74), .A2 (A_in[2]));
NAND2_X1 i_93 (.ZN (n_75), .A1 (n_59), .A2 (n_76));
INV_X1 i_92 (.ZN (p_0[2]), .A (n_75));
NAND3_X1 i_11 (.ZN (n_72), .A1 (n_83), .A2 (A_in[6]), .A3 (n_98));
INV_X1 i_87 (.ZN (n_71), .A (A_in[25]));
INV_X1 i_86 (.ZN (n_70), .A (A_in[24]));
INV_X1 i_85 (.ZN (n_69), .A (A_in[23]));
NOR2_X4 slo__mro_c290 (.ZN (n_101), .A1 (slo__mro_n189), .A2 (A_in[0]));
INV_X4 i_83 (.ZN (n_68), .A (n_96));
INV_X2 i_82 (.ZN (n_67), .A (A_in[11]));
NAND4_X4 i_80 (.ZN (n_65), .A1 (n_90), .A2 (n_88), .A3 (n_67), .A4 (n_103));
INV_X1 i_79 (.ZN (n_64), .A (A_in[15]));
INV_X2 i_76 (.ZN (n_62), .A (A_in[13]));
NAND4_X2 i_75 (.ZN (n_61), .A1 (n_62), .A2 (n_66), .A3 (n_64), .A4 (A_in[14]));
INV_X2 i_74 (.ZN (n_60), .A (n_61));
NAND4_X4 i_73 (.ZN (n_48), .A1 (slo__n611), .A2 (n_68), .A3 (n_53), .A4 (n_60));
INV_X2 i_72 (.ZN (n_49), .A (n_48));
INV_X1 i_71 (.ZN (n_56), .A (A_in[18]));
INV_X2 i_56 (.ZN (n_54), .A (A_in[17]));
INV_X1 i_54 (.ZN (n_28), .A (A_in[16]));
NAND3_X2 i_53 (.ZN (n_46), .A1 (n_54), .A2 (n_28), .A3 (n_56));
OR2_X2 i_52 (.ZN (n_22), .A1 (n_46), .A2 (A_in[19]));
INV_X1 i_42 (.ZN (n_16), .A (n_22));
OR3_X4 i_41 (.ZN (n_11), .A1 (A_in[20]), .A2 (A_in[21]), .A3 (A_in[22]));
INV_X2 i_40 (.ZN (n_10), .A (n_11));
CLKBUF_X1 slo__mro_c654 (.Z (slo__mro_n471), .A (n_87));
INV_X2 i_32 (.ZN (n_41), .A (sgo__sro_n47));
AOI21_X1 i_31 (.ZN (n_9), .A (n_71), .B1 (n_41), .B2 (n_70));
NAND3_X1 i_30 (.ZN (n_30), .A1 (n_41), .A2 (n_71), .A3 (n_70));
INV_X1 i_24 (.ZN (n_8), .A (n_30));
NOR2_X1 i_22 (.ZN (p_0[25]), .A1 (n_8), .A2 (n_9));
NOR2_X2 i_21 (.ZN (n_23), .A1 (n_48), .A2 (A_in[16]));
NAND2_X2 i_20 (.ZN (n_5), .A1 (n_23), .A2 (n_54));
INV_X2 i_19 (.ZN (n_21), .A (n_5));
NOR2_X1 i_18 (.ZN (n_4), .A1 (n_23), .A2 (n_54));
NOR2_X2 i_15 (.ZN (p_0[17]), .A1 (n_21), .A2 (n_4));
NAND2_X1 i_14 (.ZN (n_3), .A1 (n_85), .A2 (A_in[9]));
NAND2_X1 i_13 (.ZN (n_2), .A1 (n_86), .A2 (n_3));
INV_X2 i_12 (.ZN (p_0[9]), .A (n_2));
INV_X1 i_10 (.ZN (n_17), .A (n_94));
NOR2_X1 i_9 (.ZN (n_15), .A1 (n_94), .A2 (A_in[13]));
NAND3_X1 i_8 (.ZN (n_50), .A1 (n_62), .A2 (n_66), .A3 (opt_ipo_n1484));
NOR2_X4 i_5 (.ZN (n_45), .A1 (n_48), .A2 (n_22));
INV_X4 i_4 (.ZN (n_44), .A (n_45));
NAND2_X4 i_3 (.ZN (n_42), .A1 (opt_ipo_n1391), .A2 (n_10));
INV_X2 i_1 (.ZN (n_43), .A (n_42));
NOR2_X1 i_0 (.ZN (n_29), .A1 (sgo__sro_n47), .A2 (A_in[24]));
OR3_X1 i_78 (.ZN (n_47), .A1 (A_in[26]), .A2 (A_in[25]), .A3 (A_in[24]));
NOR3_X2 i_70 (.ZN (n_39), .A1 (sgo__sro_n47), .A2 (n_47), .A3 (A_in[27]));
INV_X2 i_69 (.ZN (n_38), .A (n_39));
NOR4_X4 i_68 (.ZN (n_37), .A1 (n_38), .A2 (A_in[28]), .A3 (A_in[30]), .A4 (A_in[29]));
XNOR2_X2 i_67 (.ZN (p_0[31]), .A (A_in[31]), .B (n_37));
NOR2_X1 slo__sro_c603 (.ZN (slo__sro_n426), .A1 (slo__sro_n427), .A2 (slo__sro_n428));
INV_X1 i_65 (.ZN (n_35), .A (slo__sro_n397));
AOI21_X2 i_64 (.ZN (p_0[30]), .A (n_37), .B1 (A_in[30]), .B2 (n_35));
NOR2_X1 slo__sro_c604 (.ZN (p_0[26]), .A1 (n_32), .A2 (slo__sro_n426));
INV_X1 i_62 (.ZN (n_33), .A (slo__mro_n327));
AOI21_X1 i_61 (.ZN (p_0[29]), .A (slo__sro_n397), .B1 (n_33), .B2 (A_in[29]));
NAND2_X1 slo__sro_c582 (.ZN (slo__sro_n407), .A1 (n_0), .A2 (A_in[7]));
NOR2_X1 i_59 (.ZN (n_32), .A1 (sgo__sro_n47), .A2 (n_47));
INV_X1 i_58 (.ZN (n_31), .A (n_32));
AOI21_X1 i_57 (.ZN (p_0[27]), .A (n_39), .B1 (A_in[27]), .B2 (n_31));
INV_X1 slo__sro_c726 (.ZN (slo__sro_n529), .A (A_in[24]));
AOI21_X2 slo__sro_c1352 (.ZN (p_0[14]), .A (n_13), .B1 (n_14), .B2 (opt_ipoPP_14));
AOI21_X1 i_50 (.ZN (p_0[23]), .A (n_41), .B1 (slo__xsl_n254), .B2 (A_in[23]));
NOR3_X4 i_49 (.ZN (n_27), .A1 (n_44), .A2 (A_in[20]), .A3 (opt_ipoPP_1));
INV_X1 i_48 (.ZN (n_26), .A (n_27));
AOI21_X2 i_47 (.ZN (p_0[22]), .A (n_43), .B1 (A_in[22]), .B2 (n_26));
NOR2_X2 i_46 (.ZN (n_25), .A1 (n_44), .A2 (A_in[20]));
INV_X1 i_45 (.ZN (n_24), .A (slo__n1132));
AOI21_X2 i_44 (.ZN (p_0[21]), .A (n_27), .B1 (n_24), .B2 (opt_ipoPP_1));
AOI21_X1 i_43 (.ZN (p_0[20]), .A (n_25), .B1 (A_in[20]), .B2 (n_44));
AND2_X1 sgo__sro_c239 (.ZN (sgo__sro_n157), .A1 (n_88), .A2 (n_90));
INV_X1 i_37 (.ZN (n_18), .A (n_19));
AOI21_X1 i_36 (.ZN (p_0[19]), .A (opt_ipo_n1391), .B1 (A_in[19]), .B2 (n_18));
AOI21_X1 i_35 (.ZN (p_0[18]), .A (n_19), .B1 (n_5), .B2 (A_in[18]));
AOI21_X1 i_33 (.ZN (p_0[16]), .A (n_23), .B1 (A_in[16]), .B2 (n_48));
INV_X1 i_29 (.ZN (n_14), .A (n_15));
NOR2_X4 i_28 (.ZN (n_13), .A1 (n_51), .A2 (n_50));
INV_X1 i_27 (.ZN (n_12), .A (n_13));
AOI21_X1 i_26 (.ZN (p_0[15]), .A (n_49), .B1 (n_12), .B2 (A_in[15]));
AOI21_X1 i_23 (.ZN (p_0[12]), .A (n_17), .B1 (n_51), .B2 (A_in[12]));
INV_X1 slo__xsl_c378 (.ZN (slo__xsl_n254), .A (slo__xsl_n255));
AOI21_X1 i_16 (.ZN (p_0[11]), .A (n_52), .B1 (n_89), .B2 (A_in[11]));
INV_X1 i_7 (.ZN (n_0), .A (n_1));
INV_X1 slo__sro_c601 (.ZN (slo__sro_n428), .A (A_in[26]));
AOI21_X1 i_2 (.ZN (p_0[3]), .A (n_101), .B1 (n_59), .B2 (A_in[3]));
NOR2_X1 slo__sro_c426 (.ZN (slo__sro_n289), .A1 (slo__sro_n290), .A2 (slo__sro_n291));
NOR2_X1 slo__sro_c427 (.ZN (p_0[28]), .A1 (slo__mro_n327), .A2 (slo__sro_n289));
INV_X1 slo__sro_c583 (.ZN (slo__sro_n406), .A (slo__sro_n407));
NOR2_X2 slo__sro_c584 (.ZN (p_0[7]), .A1 (n_55), .A2 (slo__sro_n406));
INV_X1 slo__sro_c602 (.ZN (slo__sro_n427), .A (n_30));
OR2_X1 slo__sro_c575 (.ZN (slo__sro_n398), .A1 (A_in[28]), .A2 (A_in[29]));
NOR2_X1 slo__mro_c476 (.ZN (slo__mro_n327), .A1 (n_38), .A2 (A_in[28]));
NOR2_X1 slo__sro_c576 (.ZN (slo__sro_n397), .A1 (n_38), .A2 (slo__sro_n398));
INV_X1 slo__sro_c727 (.ZN (slo__sro_n528), .A (sgo__sro_n47));
NAND3_X1 sgo__sro_c68 (.ZN (sgo__sro_n49), .A1 (n_16), .A2 (n_10), .A3 (n_69));
INV_X2 sgo__sro_c69 (.ZN (sgo__sro_n48), .A (sgo__sro_n49));
NAND2_X4 sgo__sro_c70 (.ZN (sgo__sro_n47), .A1 (n_49), .A2 (sgo__sro_n48));
INV_X1 opt_ipo_c1833 (.ZN (opt_ipo_n1484), .A (opt_ipoPP_14));
NAND2_X1 slo__mro_c655 (.ZN (n_89), .A1 (n_55), .A2 (slo__mro_n471));
INV_X1 slo__xsl_c670 (.ZN (slo__xsl_n479), .A (slo__xsl_n480));
NOR2_X1 slo__sro_c728 (.ZN (slo__sro_n527), .A1 (slo__sro_n528), .A2 (slo__sro_n529));
NOR2_X1 slo__sro_c729 (.ZN (p_0[24]), .A1 (n_29), .A2 (slo__sro_n527));
INV_X1 slo__xsl_c883 (.ZN (slo__xsl_n687), .A (n_65));
INV_X1 slo__xsl_c884 (.ZN (slo__xsl_n686), .A (slo__xsl_n687));
INV_X4 slo__c757 (.ZN (slo__n560), .A (A_in[2]));
INV_X4 slo__c1323 (.ZN (slo__n1059), .A (A_in[1]));
INV_X4 opt_ipo_c1774 (.ZN (opt_ipo_n1391), .A (slo__xsl_n796));
NAND3_X4 slo__c972 (.ZN (slo__n753), .A1 (n_84), .A2 (slo__n560), .A3 (n_105));
NAND2_X4 slo__sro_c1392 (.ZN (slo__sro_n1119), .A1 (n_101), .A2 (n_68));
NOR2_X2 slo__c844 (.ZN (slo__n646), .A1 (slo__n753), .A2 (A_in[0]));
AND2_X1 slo__sro_c1196 (.ZN (slo__sro_n938), .A1 (n_83), .A2 (n_98));
INV_X2 slo__xsl_c1021 (.ZN (slo__xsl_n796), .A (n_45));
NAND2_X1 slo__sro_c1197 (.ZN (slo__sro_n937), .A1 (n_101), .A2 (slo__sro_n938));
NOR2_X4 slo__c1166 (.ZN (slo__n913), .A1 (slo__n753), .A2 (A_in[0]));
NOR2_X4 slo__c805 (.ZN (slo__n611), .A1 (slo__mro_n189), .A2 (A_in[0]));

endmodule //datapath

module boothAlgoR4 (Res, OVF, A, B, clk, reset, enable);

output OVF;
output [63:0] Res;
input [31:0] A;
input [31:0] B;
input clk;
input enable;
input reset;
wire opt_ipo_n5239;
wire CLOCK_slh_n7157;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire \A_imm_2s_complement[31] ;
wire \A_imm_2s_complement[30] ;
wire \A_imm_2s_complement[29] ;
wire \A_imm_2s_complement[28] ;
wire \A_imm_2s_complement[27] ;
wire \A_imm_2s_complement[26] ;
wire \A_imm_2s_complement[25] ;
wire \A_imm_2s_complement[24] ;
wire \A_imm_2s_complement[23] ;
wire \A_imm_2s_complement[22] ;
wire \A_imm_2s_complement[21] ;
wire \A_imm_2s_complement[20] ;
wire \A_imm_2s_complement[19] ;
wire \A_imm_2s_complement[18] ;
wire \A_imm_2s_complement[17] ;
wire \A_imm_2s_complement[16] ;
wire \A_imm_2s_complement[15] ;
wire \A_imm_2s_complement[14] ;
wire \A_imm_2s_complement[13] ;
wire \A_imm_2s_complement[12] ;
wire \A_imm_2s_complement[11] ;
wire \A_imm_2s_complement[10] ;
wire \A_imm_2s_complement[9] ;
wire \A_imm_2s_complement[8] ;
wire \A_imm_2s_complement[7] ;
wire \A_imm_2s_complement[6] ;
wire \A_imm_2s_complement[5] ;
wire \A_imm_2s_complement[4] ;
wire \A_imm_2s_complement[3] ;
wire \A_imm_2s_complement[2] ;
wire \A_imm_2s_complement[1] ;
wire hfn_ipo_n45;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire \aggregated_res[14][63] ;
wire \aggregated_res[14][62] ;
wire \aggregated_res[14][61] ;
wire \aggregated_res[14][60] ;
wire \aggregated_res[14][59] ;
wire \aggregated_res[14][58] ;
wire \aggregated_res[14][57] ;
wire \aggregated_res[14][56] ;
wire \aggregated_res[14][55] ;
wire \aggregated_res[14][54] ;
wire \aggregated_res[14][53] ;
wire \aggregated_res[14][52] ;
wire \aggregated_res[14][51] ;
wire \aggregated_res[14][50] ;
wire \aggregated_res[14][49] ;
wire \aggregated_res[14][48] ;
wire \aggregated_res[14][47] ;
wire \aggregated_res[14][46] ;
wire \aggregated_res[14][45] ;
wire \aggregated_res[14][44] ;
wire \aggregated_res[14][43] ;
wire \aggregated_res[14][42] ;
wire \aggregated_res[14][41] ;
wire \aggregated_res[14][40] ;
wire \aggregated_res[14][39] ;
wire \aggregated_res[14][38] ;
wire \aggregated_res[14][37] ;
wire \aggregated_res[14][36] ;
wire \aggregated_res[14][35] ;
wire \aggregated_res[14][34] ;
wire \aggregated_res[14][33] ;
wire \aggregated_res[14][32] ;
wire \aggregated_res[14][31] ;
wire \aggregated_res[14][30] ;
wire \aggregated_res[14][29] ;
wire \aggregated_res[14][28] ;
wire \aggregated_res[14][27] ;
wire \aggregated_res[14][26] ;
wire \aggregated_res[14][25] ;
wire \aggregated_res[14][24] ;
wire \aggregated_res[14][23] ;
wire \aggregated_res[14][22] ;
wire \aggregated_res[14][21] ;
wire \aggregated_res[14][20] ;
wire \aggregated_res[14][19] ;
wire \aggregated_res[14][18] ;
wire \aggregated_res[14][17] ;
wire \aggregated_res[14][16] ;
wire \aggregated_res[14][15] ;
wire \aggregated_res[14][14] ;
wire \aggregated_res[14][13] ;
wire \aggregated_res[14][12] ;
wire \aggregated_res[14][11] ;
wire \aggregated_res[14][10] ;
wire \aggregated_res[14][9] ;
wire \aggregated_res[14][8] ;
wire \aggregated_res[14][7] ;
wire \aggregated_res[14][6] ;
wire \aggregated_res[14][5] ;
wire \aggregated_res[14][4] ;
wire \aggregated_res[14][3] ;
wire \aggregated_res[14][2] ;
wire hfn_ipo_n44;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire A_in;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire B_in;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_169;
wire n_0_170;
wire n_0_171;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_176;
wire n_0_177;
wire n_0_178;
wire n_0_179;
wire n_0_180;
wire n_0_181;
wire n_0_182;
wire n_0_183;
wire n_0_184;
wire n_0_185;
wire n_0_186;
wire n_0_187;
wire n_0_1_74;
wire opt_ipo_n5162;
wire n_0_1_76;
wire n_0_1_77;
wire slo__sro_n1621;
wire CLOCK_slo__sro_n6808;
wire n_0_1_81;
wire sgo__n836;
wire n_0_317;
wire slo__n2107;
wire slo__sro_n2079;
wire n_0_1_91;
wire n_0_319;
wire n_0_1_92;
wire n_0_320;
wire n_0_1_93;
wire n_0_321;
wire n_0_1_94;
wire n_0_322;
wire n_0_1_95;
wire n_0_323;
wire n_0_1_96;
wire n_0_324;
wire n_0_1_97;
wire n_0_325;
wire n_0_1_98;
wire n_0_326;
wire n_0_1_99;
wire n_0_327;
wire n_0_1_100;
wire n_0_328;
wire n_0_1_101;
wire n_0_329;
wire n_0_1_102;
wire n_0_330;
wire n_0_1_103;
wire n_0_331;
wire n_0_1_104;
wire n_0_332;
wire n_0_1_105;
wire n_0_333;
wire n_0_1_106;
wire n_0_334;
wire n_0_1_107;
wire n_0_335;
wire n_0_1_108;
wire n_0_336;
wire n_0_1_109;
wire n_0_337;
wire n_0_1_110;
wire n_0_338;
wire n_0_1_111;
wire n_0_339;
wire n_0_1_112;
wire n_0_340;
wire n_0_1_113;
wire n_0_341;
wire n_0_1_114;
wire n_0_342;
wire n_0_1_115;
wire n_0_343;
wire n_0_1_116;
wire n_0_344;
wire n_0_1_117;
wire n_0_345;
wire n_0_1_118;
wire n_0_346;
wire n_0_1_119;
wire n_0_347;
wire n_0_1_120;
wire n_0_348;
wire n_0_1_121;
wire n_0_349;
wire n_0_1_122;
wire n_0_1_123;
wire n_0_1_124;
wire n_0_1_125;
wire n_0_1_126;
wire n_0_1_127;
wire n_0_1_128;
wire n_0_1_129;
wire n_0_1_130;
wire n_0_1_131;
wire n_0_1_132;
wire n_0_1_133;
wire n_0_350;
wire n_0_351;
wire n_0_1_134;
wire n_0_1_135;
wire n_0_352;
wire n_0_1_136;
wire n_0_353;
wire n_0_1_137;
wire n_0_354;
wire n_0_1_138;
wire n_0_355;
wire n_0_1_139;
wire n_0_356;
wire n_0_1_140;
wire n_0_357;
wire n_0_1_141;
wire n_0_358;
wire n_0_1_142;
wire n_0_359;
wire n_0_1_143;
wire n_0_360;
wire n_0_1_144;
wire n_0_361;
wire n_0_1_145;
wire n_0_362;
wire n_0_1_146;
wire n_0_363;
wire n_0_1_147;
wire n_0_364;
wire n_0_1_148;
wire n_0_365;
wire n_0_1_149;
wire n_0_366;
wire n_0_1_150;
wire n_0_367;
wire n_0_1_151;
wire n_0_368;
wire n_0_1_152;
wire n_0_369;
wire n_0_1_153;
wire n_0_370;
wire n_0_1_154;
wire n_0_371;
wire n_0_1_155;
wire n_0_372;
wire n_0_1_156;
wire n_0_373;
wire n_0_1_157;
wire n_0_374;
wire n_0_1_158;
wire n_0_375;
wire n_0_1_159;
wire n_0_376;
wire n_0_1_160;
wire n_0_377;
wire n_0_1_161;
wire n_0_378;
wire n_0_1_162;
wire n_0_379;
wire n_0_1_163;
wire n_0_380;
wire n_0_1_164;
wire n_0_381;
wire n_0_1_165;
wire n_0_1_166;
wire n_0_1_167;
wire n_0_1_168;
wire n_0_1_169;
wire n_0_1_170;
wire n_0_382;
wire n_0_1_171;
wire n_0_1_172;
wire n_0_1_173;
wire n_0_1_174;
wire n_0_1_175;
wire n_0_1_176;
wire n_0_1_177;
wire n_0_1_178;
wire n_0_1_179;
wire n_0_383;
wire n_0_384;
wire n_0_1_180;
wire n_0_1_181;
wire n_0_385;
wire n_0_1_182;
wire n_0_386;
wire n_0_1_183;
wire n_0_387;
wire n_0_1_184;
wire n_0_388;
wire n_0_1_185;
wire n_0_389;
wire n_0_1_186;
wire n_0_390;
wire n_0_1_187;
wire n_0_391;
wire n_0_1_188;
wire n_0_392;
wire n_0_1_189;
wire n_0_393;
wire n_0_1_190;
wire n_0_394;
wire n_0_1_191;
wire n_0_395;
wire n_0_1_192;
wire n_0_396;
wire n_0_1_193;
wire n_0_397;
wire n_0_1_194;
wire n_0_398;
wire n_0_1_195;
wire n_0_399;
wire n_0_1_196;
wire n_0_400;
wire n_0_1_197;
wire n_0_401;
wire n_0_1_198;
wire n_0_402;
wire n_0_1_199;
wire n_0_403;
wire n_0_1_200;
wire n_0_404;
wire n_0_1_201;
wire n_0_405;
wire n_0_1_202;
wire n_0_406;
wire n_0_1_203;
wire n_0_407;
wire n_0_1_204;
wire n_0_408;
wire n_0_1_205;
wire n_0_409;
wire n_0_1_206;
wire n_0_410;
wire n_0_1_207;
wire n_0_411;
wire n_0_1_208;
wire n_0_412;
wire n_0_1_209;
wire n_0_413;
wire n_0_1_210;
wire n_0_414;
wire n_0_1_211;
wire n_0_1_212;
wire n_0_1_213;
wire n_0_1_214;
wire n_0_1_215;
wire n_0_1_216;
wire n_0_415;
wire n_0_1_217;
wire n_0_1_218;
wire opt_ipo_n5653;
wire n_0_1_220;
wire n_0_1_221;
wire n_0_1_222;
wire n_0_416;
wire n_0_417;
wire n_0_1_223;
wire n_0_1_224;
wire n_0_418;
wire n_0_1_225;
wire n_0_419;
wire n_0_1_226;
wire n_0_420;
wire n_0_1_227;
wire n_0_421;
wire n_0_1_228;
wire n_0_422;
wire n_0_1_229;
wire n_0_423;
wire n_0_1_230;
wire n_0_424;
wire n_0_1_231;
wire n_0_425;
wire n_0_1_232;
wire n_0_426;
wire n_0_1_233;
wire n_0_427;
wire n_0_1_234;
wire n_0_428;
wire n_0_1_235;
wire n_0_429;
wire n_0_1_236;
wire n_0_430;
wire n_0_1_237;
wire n_0_431;
wire n_0_1_238;
wire n_0_432;
wire n_0_1_239;
wire n_0_433;
wire n_0_1_240;
wire n_0_434;
wire n_0_1_241;
wire n_0_435;
wire n_0_1_242;
wire n_0_436;
wire n_0_1_243;
wire n_0_437;
wire n_0_1_244;
wire n_0_438;
wire n_0_1_245;
wire n_0_439;
wire n_0_1_246;
wire n_0_440;
wire n_0_1_247;
wire n_0_441;
wire n_0_1_248;
wire n_0_442;
wire n_0_1_249;
wire n_0_443;
wire n_0_1_250;
wire n_0_444;
wire n_0_1_251;
wire n_0_445;
wire n_0_1_252;
wire n_0_446;
wire n_0_1_253;
wire n_0_447;
wire n_0_1_254;
wire n_0_1_255;
wire n_0_1_256;
wire n_0_1_257;
wire n_0_1_258;
wire n_0_1_259;
wire n_0_448;
wire n_0_1_260;
wire n_0_1_261;
wire n_0_1_262;
wire n_0_1_263;
wire n_0_1_264;
wire n_0_1_265;
wire n_0_449;
wire n_0_450;
wire slo__n3696;
wire n_0_1_267;
wire n_0_451;
wire n_0_1_268;
wire n_0_452;
wire n_0_1_269;
wire n_0_453;
wire n_0_1_270;
wire n_0_454;
wire n_0_1_271;
wire n_0_455;
wire n_0_1_272;
wire n_0_456;
wire n_0_1_273;
wire n_0_457;
wire n_0_1_274;
wire n_0_458;
wire n_0_1_275;
wire n_0_459;
wire n_0_1_276;
wire n_0_460;
wire n_0_1_277;
wire n_0_461;
wire n_0_1_278;
wire n_0_462;
wire n_0_1_279;
wire n_0_463;
wire n_0_1_280;
wire n_0_464;
wire n_0_1_281;
wire n_0_465;
wire n_0_1_282;
wire n_0_466;
wire n_0_1_283;
wire n_0_467;
wire n_0_1_284;
wire n_0_468;
wire n_0_1_285;
wire n_0_469;
wire n_0_1_286;
wire n_0_470;
wire n_0_1_287;
wire n_0_471;
wire n_0_1_288;
wire n_0_472;
wire n_0_1_289;
wire n_0_473;
wire n_0_1_290;
wire n_0_474;
wire n_0_1_291;
wire n_0_475;
wire n_0_1_292;
wire n_0_476;
wire n_0_1_293;
wire n_0_477;
wire n_0_1_294;
wire n_0_478;
wire n_0_1_295;
wire n_0_479;
wire n_0_1_296;
wire n_0_480;
wire n_0_1_297;
wire n_0_1_298;
wire n_0_1_299;
wire n_0_1_300;
wire n_0_1_301;
wire n_0_1_302;
wire n_0_481;
wire n_0_1_303;
wire n_0_1_304;
wire n_0_1_305;
wire n_0_1_306;
wire opt_ipo_n5159;
wire n_0_1_308;
wire n_0_482;
wire n_0_483;
wire n_0_1_309;
wire n_0_1_310;
wire n_0_484;
wire n_0_1_311;
wire n_0_485;
wire n_0_1_312;
wire n_0_486;
wire n_0_1_313;
wire n_0_487;
wire n_0_1_314;
wire n_0_488;
wire n_0_1_315;
wire n_0_489;
wire n_0_1_316;
wire n_0_490;
wire n_0_1_317;
wire n_0_491;
wire n_0_1_318;
wire n_0_492;
wire n_0_1_319;
wire n_0_493;
wire n_0_1_320;
wire n_0_494;
wire n_0_1_321;
wire n_0_495;
wire n_0_1_322;
wire n_0_496;
wire n_0_1_323;
wire n_0_497;
wire n_0_1_324;
wire n_0_498;
wire n_0_1_325;
wire n_0_499;
wire n_0_1_326;
wire n_0_500;
wire n_0_1_327;
wire n_0_501;
wire n_0_1_328;
wire n_0_502;
wire n_0_1_329;
wire n_0_503;
wire n_0_1_330;
wire n_0_504;
wire n_0_1_331;
wire n_0_505;
wire n_0_1_332;
wire n_0_506;
wire n_0_1_333;
wire n_0_507;
wire n_0_1_334;
wire n_0_508;
wire n_0_1_335;
wire n_0_509;
wire n_0_1_336;
wire n_0_510;
wire n_0_1_337;
wire n_0_511;
wire n_0_1_338;
wire n_0_512;
wire n_0_1_339;
wire n_0_513;
wire n_0_1_340;
wire spd__n7595;
wire n_0_1_342;
wire n_0_1_343;
wire n_0_1_344;
wire n_0_1_345;
wire n_0_514;
wire n_0_1_346;
wire n_0_1_347;
wire n_0_1_348;
wire n_0_1_349;
wire n_0_1_350;
wire n_0_1_351;
wire n_0_515;
wire n_0_516;
wire n_0_1_352;
wire n_0_1_353;
wire n_0_517;
wire n_0_1_354;
wire n_0_518;
wire n_0_1_355;
wire n_0_519;
wire n_0_1_356;
wire n_0_520;
wire n_0_1_357;
wire n_0_521;
wire n_0_1_358;
wire n_0_522;
wire n_0_1_359;
wire n_0_523;
wire n_0_1_360;
wire n_0_524;
wire n_0_1_361;
wire n_0_525;
wire n_0_1_362;
wire n_0_526;
wire n_0_1_363;
wire n_0_527;
wire n_0_1_364;
wire n_0_528;
wire n_0_1_365;
wire n_0_529;
wire n_0_1_366;
wire n_0_530;
wire n_0_1_367;
wire n_0_531;
wire n_0_1_368;
wire n_0_532;
wire n_0_1_369;
wire n_0_533;
wire n_0_1_370;
wire n_0_534;
wire n_0_1_371;
wire n_0_535;
wire n_0_1_372;
wire n_0_536;
wire n_0_1_373;
wire n_0_537;
wire n_0_1_374;
wire n_0_538;
wire n_0_1_375;
wire n_0_539;
wire n_0_1_376;
wire n_0_540;
wire n_0_1_377;
wire n_0_541;
wire n_0_1_378;
wire n_0_542;
wire n_0_1_379;
wire n_0_543;
wire n_0_1_380;
wire n_0_544;
wire n_0_1_381;
wire n_0_545;
wire n_0_1_382;
wire n_0_546;
wire n_0_1_383;
wire n_0_1_384;
wire n_0_1_385;
wire n_0_1_386;
wire n_0_1_387;
wire n_0_1_388;
wire n_0_547;
wire n_0_1_389;
wire n_0_1_390;
wire n_0_1_391;
wire n_0_1_392;
wire n_0_1_393;
wire n_0_1_394;
wire n_0_548;
wire n_0_549;
wire n_0_1_395;
wire n_0_1_396;
wire n_0_550;
wire n_0_1_397;
wire n_0_551;
wire sgo__n844;
wire n_0_552;
wire n_0_1_399;
wire n_0_553;
wire n_0_1_400;
wire n_0_554;
wire n_0_1_401;
wire n_0_555;
wire n_0_1_402;
wire n_0_556;
wire n_0_1_403;
wire n_0_557;
wire n_0_1_404;
wire n_0_558;
wire n_0_1_405;
wire n_0_559;
wire n_0_1_406;
wire n_0_560;
wire n_0_1_407;
wire n_0_561;
wire n_0_1_408;
wire n_0_562;
wire n_0_1_409;
wire n_0_563;
wire n_0_1_410;
wire n_0_564;
wire n_0_1_411;
wire n_0_565;
wire n_0_1_412;
wire n_0_566;
wire n_0_1_413;
wire n_0_567;
wire n_0_1_414;
wire n_0_568;
wire n_0_1_415;
wire n_0_569;
wire n_0_1_416;
wire n_0_570;
wire n_0_1_417;
wire n_0_571;
wire n_0_1_418;
wire n_0_572;
wire n_0_1_419;
wire n_0_573;
wire n_0_1_420;
wire n_0_574;
wire n_0_1_421;
wire n_0_575;
wire n_0_1_422;
wire n_0_576;
wire n_0_1_423;
wire n_0_577;
wire n_0_1_424;
wire n_0_578;
wire n_0_1_425;
wire n_0_579;
wire n_0_1_426;
wire n_0_1_427;
wire n_0_1_428;
wire n_0_1_429;
wire n_0_1_430;
wire n_0_1_431;
wire n_0_580;
wire n_0_1_432;
wire n_0_1_433;
wire n_0_1_434;
wire n_0_1_435;
wire n_0_1_436;
wire n_0_1_437;
wire n_0_581;
wire n_0_582;
wire n_0_1_438;
wire n_0_1_439;
wire n_0_583;
wire n_0_1_440;
wire n_0_584;
wire n_0_1_441;
wire n_0_585;
wire n_0_1_442;
wire n_0_586;
wire n_0_1_443;
wire n_0_587;
wire n_0_1_444;
wire n_0_588;
wire n_0_1_445;
wire n_0_589;
wire n_0_1_446;
wire n_0_590;
wire n_0_1_447;
wire n_0_591;
wire n_0_1_448;
wire n_0_592;
wire n_0_1_449;
wire n_0_593;
wire n_0_1_450;
wire n_0_594;
wire n_0_1_451;
wire n_0_595;
wire n_0_1_452;
wire n_0_596;
wire n_0_1_453;
wire n_0_597;
wire n_0_1_454;
wire n_0_598;
wire n_0_1_455;
wire n_0_599;
wire n_0_1_456;
wire n_0_600;
wire n_0_1_457;
wire n_0_601;
wire n_0_1_458;
wire n_0_602;
wire n_0_1_459;
wire n_0_603;
wire n_0_1_460;
wire n_0_604;
wire n_0_1_461;
wire n_0_605;
wire n_0_1_462;
wire n_0_606;
wire n_0_1_463;
wire n_0_607;
wire n_0_1_464;
wire n_0_608;
wire n_0_1_465;
wire n_0_609;
wire n_0_1_466;
wire n_0_610;
wire n_0_1_467;
wire n_0_611;
wire n_0_1_468;
wire n_0_612;
wire n_0_1_469;
wire n_0_1_470;
wire n_0_1_471;
wire n_0_1_472;
wire n_0_1_473;
wire n_0_1_474;
wire n_0_613;
wire n_0_1_475;
wire n_0_1_476;
wire n_0_1_477;
wire n_0_1_478;
wire n_0_1_479;
wire n_0_1_480;
wire n_0_614;
wire n_0_615;
wire n_0_1_481;
wire n_0_1_482;
wire n_0_616;
wire n_0_1_483;
wire n_0_617;
wire n_0_1_484;
wire n_0_618;
wire n_0_1_485;
wire n_0_619;
wire n_0_1_486;
wire n_0_620;
wire n_0_1_487;
wire n_0_621;
wire n_0_1_488;
wire n_0_622;
wire n_0_1_489;
wire n_0_623;
wire n_0_1_490;
wire n_0_624;
wire n_0_1_491;
wire n_0_625;
wire n_0_1_492;
wire n_0_626;
wire n_0_1_493;
wire n_0_627;
wire n_0_1_494;
wire n_0_628;
wire n_0_1_495;
wire n_0_629;
wire n_0_1_496;
wire n_0_630;
wire n_0_1_497;
wire n_0_631;
wire n_0_1_498;
wire n_0_632;
wire n_0_1_499;
wire n_0_633;
wire n_0_1_500;
wire n_0_634;
wire n_0_1_501;
wire n_0_635;
wire n_0_1_502;
wire n_0_636;
wire n_0_1_503;
wire n_0_637;
wire n_0_1_504;
wire n_0_638;
wire n_0_1_505;
wire n_0_639;
wire n_0_1_506;
wire n_0_640;
wire n_0_1_507;
wire n_0_641;
wire n_0_1_508;
wire n_0_642;
wire n_0_1_509;
wire n_0_643;
wire n_0_1_510;
wire n_0_644;
wire n_0_1_511;
wire n_0_645;
wire n_0_1_512;
wire n_0_1_513;
wire n_0_1_514;
wire sph__n7810;
wire n_0_1_516;
wire n_0_1_517;
wire n_0_646;
wire n_0_1_518;
wire n_0_1_519;
wire n_0_1_520;
wire n_0_1_521;
wire n_0_1_522;
wire n_0_1_523;
wire n_0_647;
wire n_0_648;
wire n_0_1_524;
wire n_0_1_525;
wire n_0_649;
wire n_0_1_526;
wire n_0_650;
wire n_0_1_527;
wire n_0_651;
wire n_0_1_528;
wire n_0_652;
wire n_0_1_529;
wire n_0_653;
wire n_0_1_530;
wire n_0_654;
wire n_0_1_531;
wire n_0_655;
wire opt_ipo_n5703;
wire n_0_656;
wire n_0_1_533;
wire n_0_657;
wire n_0_1_534;
wire n_0_658;
wire n_0_1_535;
wire n_0_659;
wire n_0_1_536;
wire n_0_660;
wire n_0_1_537;
wire n_0_661;
wire n_0_1_538;
wire n_0_662;
wire n_0_1_539;
wire n_0_663;
wire n_0_1_540;
wire n_0_664;
wire n_0_1_541;
wire n_0_665;
wire n_0_1_542;
wire n_0_666;
wire n_0_1_543;
wire n_0_667;
wire n_0_1_544;
wire n_0_668;
wire n_0_1_545;
wire n_0_669;
wire n_0_1_546;
wire n_0_670;
wire n_0_1_547;
wire n_0_671;
wire n_0_1_548;
wire n_0_672;
wire n_0_1_549;
wire n_0_673;
wire slo__n3026;
wire n_0_674;
wire n_0_1_551;
wire n_0_675;
wire n_0_1_552;
wire n_0_676;
wire n_0_1_553;
wire n_0_1_560;
wire n_0_679;
wire n_0_1_561;
wire n_0_1_562;
wire n_0_1_563;
wire slo___n3078;
wire n_0_1_565;
wire n_0_1_566;
wire n_0_680;
wire n_0_681;
wire n_0_1_567;
wire n_0_1_568;
wire n_0_682;
wire n_0_1_569;
wire n_0_683;
wire n_0_1_570;
wire n_0_684;
wire n_0_1_571;
wire n_0_685;
wire slo__sro_n3368;
wire n_0_686;
wire n_0_1_573;
wire n_0_687;
wire n_0_1_574;
wire n_0_688;
wire n_0_1_575;
wire n_0_689;
wire n_0_1_576;
wire slo__n1615;
wire n_0_1_577;
wire n_0_691;
wire n_0_1_578;
wire n_0_692;
wire n_0_1_579;
wire n_0_693;
wire n_0_1_580;
wire n_0_694;
wire n_0_1_581;
wire n_0_695;
wire n_0_1_582;
wire n_0_696;
wire n_0_1_583;
wire n_0_697;
wire n_0_1_584;
wire n_0_698;
wire n_0_1_585;
wire n_0_699;
wire n_0_1_586;
wire n_0_700;
wire n_0_1_587;
wire n_0_701;
wire n_0_1_588;
wire n_0_703;
wire n_0_1_590;
wire n_0_704;
wire n_0_1_591;
wire n_0_705;
wire n_0_1_592;
wire n_0_706;
wire n_0_1_593;
wire n_0_707;
wire n_0_1_594;
wire n_0_708;
wire slo__n3281;
wire n_0_709;
wire n_0_1_596;
wire n_0_711;
wire n_0_1_598;
wire n_0_1_603;
wire n_0_712;
wire n_0_1_604;
wire n_0_1_605;
wire n_0_1_607;
wire n_0_1_608;
wire n_0_1_609;
wire n_0_713;
wire n_0_714;
wire n_0_1_610;
wire n_0_1_611;
wire n_0_715;
wire n_0_1_612;
wire n_0_716;
wire n_0_1_613;
wire n_0_717;
wire n_0_1_614;
wire n_0_718;
wire n_0_1_615;
wire n_0_719;
wire n_0_1_616;
wire n_0_720;
wire n_0_1_617;
wire n_0_721;
wire n_0_1_618;
wire n_0_722;
wire n_0_1_619;
wire n_0_723;
wire n_0_1_620;
wire n_0_724;
wire n_0_1_621;
wire n_0_725;
wire n_0_1_622;
wire n_0_726;
wire n_0_1_623;
wire n_0_727;
wire n_0_1_624;
wire n_0_728;
wire n_0_1_625;
wire n_0_729;
wire n_0_1_626;
wire n_0_730;
wire n_0_1_627;
wire n_0_731;
wire n_0_1_628;
wire n_0_732;
wire n_0_1_629;
wire n_0_733;
wire n_0_1_630;
wire n_0_734;
wire n_0_1_631;
wire n_0_735;
wire n_0_1_632;
wire n_0_736;
wire n_0_1_633;
wire n_0_737;
wire n_0_1_634;
wire n_0_738;
wire n_0_1_635;
wire n_0_740;
wire n_0_1_637;
wire n_0_741;
wire n_0_1_638;
wire n_0_742;
wire n_0_1_639;
wire n_0_744;
wire n_0_1_641;
wire n_0_1_646;
wire n_0_745;
wire n_0_1_647;
wire n_0_1_648;
wire n_0_1_649;
wire n_0_1_650;
wire n_0_1_651;
wire n_0_746;
wire n_0_747;
wire n_0_1_653;
wire n_0_1_654;
wire n_0_748;
wire n_0_1_655;
wire n_0_749;
wire n_0_1_656;
wire n_0_750;
wire slo__sro_n2477;
wire n_0_751;
wire n_0_1_658;
wire n_0_752;
wire n_0_1_659;
wire n_0_753;
wire n_0_1_660;
wire n_0_754;
wire n_0_1_661;
wire n_0_755;
wire n_0_1_662;
wire n_0_756;
wire n_0_1_663;
wire n_0_757;
wire n_0_1_664;
wire n_0_758;
wire n_0_1_665;
wire n_0_759;
wire n_0_1_666;
wire n_0_760;
wire n_0_1_667;
wire n_0_761;
wire n_0_1_668;
wire n_0_762;
wire CLOCK_slh__n7169;
wire n_0_763;
wire n_0_1_670;
wire CLOCK_slo__mro_n6798;
wire n_0_1_671;
wire n_0_765;
wire n_0_1_672;
wire n_0_766;
wire n_0_1_673;
wire n_0_767;
wire n_0_1_674;
wire n_0_768;
wire n_0_1_675;
wire n_0_769;
wire n_0_1_676;
wire n_0_770;
wire n_0_1_677;
wire n_0_771;
wire n_0_1_678;
wire n_0_773;
wire n_0_1_680;
wire n_0_774;
wire n_0_1_681;
wire n_0_775;
wire n_0_1_682;
wire n_0_776;
wire n_0_1_683;
wire n_0_777;
wire n_0_1_684;
wire n_0_1_689;
wire n_0_778;
wire n_0_1_690;
wire n_0_1_691;
wire CLOCK_slo__sro_n6742;
wire n_0_1_693;
wire n_0_1_694;
wire n_0_1_695;
wire n_0_779;
wire n_0_780;
wire n_0_1_696;
wire n_0_1_697;
wire n_0_781;
wire n_0_1_698;
wire n_0_782;
wire n_0_1_699;
wire n_0_783;
wire n_0_1_700;
wire n_0_784;
wire n_0_1_701;
wire n_0_786;
wire n_0_1_703;
wire n_0_787;
wire n_0_1_704;
wire n_0_788;
wire n_0_1_705;
wire n_0_789;
wire n_0_1_706;
wire n_0_790;
wire n_0_1_707;
wire n_0_791;
wire n_0_1_708;
wire n_0_792;
wire n_0_1_709;
wire n_0_793;
wire n_0_1_710;
wire n_0_794;
wire n_0_1_711;
wire n_0_795;
wire n_0_1_712;
wire n_0_796;
wire n_0_1_713;
wire n_0_798;
wire n_0_1_715;
wire n_0_799;
wire n_0_1_716;
wire n_0_800;
wire n_0_1_717;
wire n_0_802;
wire n_0_1_719;
wire n_0_803;
wire n_0_1_720;
wire n_0_804;
wire n_0_1_721;
wire n_0_805;
wire n_0_1_722;
wire n_0_808;
wire n_0_1_725;
wire n_0_1_732;
wire n_0_811;
wire n_0_1_733;
wire n_0_1_734;
wire n_0_1_735;
wire n_0_1_736;
wire n_0_1_737;
wire n_0_1_738;
wire n_0_812;
wire n_0_1_739;
wire n_0_814;
wire n_0_1_740;
wire n_0_815;
wire n_0_1_741;
wire n_0_816;
wire n_0_1_742;
wire n_0_817;
wire n_0_1_743;
wire n_0_818;
wire n_0_1_744;
wire n_0_819;
wire n_0_1_745;
wire n_0_820;
wire n_0_1_746;
wire n_0_821;
wire n_0_1_747;
wire n_0_822;
wire n_0_1_748;
wire n_0_824;
wire n_0_1_750;
wire n_0_825;
wire n_0_1_751;
wire n_0_830;
wire n_0_1_756;
wire n_0_831;
wire n_0_1_757;
wire n_0_832;
wire n_0_1_758;
wire n_0_833;
wire n_0_1_759;
wire n_0_834;
wire n_0_1_760;
wire slo___n3416;
wire n_0_1_761;
wire n_0_836;
wire n_0_1_762;
wire n_0_837;
wire n_0_1_763;
wire n_0_838;
wire n_0_1_764;
wire n_0_839;
wire n_0_1_765;
wire n_0_840;
wire n_0_1_766;
wire n_0_842;
wire n_0_1_768;
wire n_0_1_774;
wire \A_imm[31] ;
wire \A_imm[30] ;
wire \A_imm[29] ;
wire \A_imm[28] ;
wire \A_imm[27] ;
wire \A_imm[24] ;
wire \A_imm[23] ;
wire \A_imm[22] ;
wire opt_ipo_n5683;
wire opt_ipo_n5720;
wire \A_imm[18] ;
wire sph__n7808;
wire \A_imm[16] ;
wire \A_imm[14] ;
wire \A_imm[13] ;
wire \A_imm[12] ;
wire CLOCK_slh__n7189;
wire opt_ipo_n5794;
wire \A_imm[9] ;
wire spw__n7740;
wire \A_imm[7] ;
wire \A_imm[6] ;
wire opt_ipo_n5146;
wire \A_imm[4] ;
wire \A_imm[3] ;
wire \A_imm[2] ;
wire \A_imm[1] ;
wire opt_ipo_n5679;
wire n_0_1_781;
wire n_0_1_782;
wire n_0_1_783;
wire n_0_1_787;
wire n_0_1_788;
wire n_0_1_789;
wire n_0_1_790;
wire n_0_1_791;
wire n_0_1_792;
wire n_0_1_793;
wire n_0_1_794;
wire n_0_1_795;
wire n_0_1_797;
wire n_0_1_798;
wire n_0_1_799;
wire n_0_1_800;
wire n_0_1_801;
wire n_0_1_803;
wire n_0_1_805;
wire n_0_1_807;
wire n_0_1_809;
wire n_0_1_811;
wire n_0_1_812;
wire n_0_1_813;
wire n_0_1_814;
wire n_0_1_815;
wire CLOCK_slo__sro_n6743;
wire n_0_1_817;
wire n_0_1_819;
wire n_0_1_820;
wire n_0_1_821;
wire n_0_1_822;
wire n_0_1_823;
wire n_0_1_825;
wire n_0_1_827;
wire n_0_1_829;
wire n_0_1_831;
wire n_0_1_833;
wire n_0_1_835;
wire n_0_1_839;
wire n_0_1_840;
wire n_0_1_841;
wire n_0_1_842;
wire n_0_1_843;
wire n_0_1_844;
wire n_0_1_845;
wire n_0_1_846;
wire n_0_1_847;
wire n_0_1_848;
wire n_0_1_849;
wire n_0_1_850;
wire n_0_1_851;
wire n_0_1_852;
wire n_0_1_853;
wire n_0_1_854;
wire n_0_1_855;
wire n_0_1_856;
wire n_0_1_857;
wire n_0_1_858;
wire n_0_1_859;
wire n_0_1_860;
wire n_0_1_861;
wire n_0_1_862;
wire n_0_1_863;
wire n_0_1_864;
wire n_0_1_865;
wire n_0_1_866;
wire n_0_1_867;
wire n_0_1_868;
wire n_0_1_784;
wire n_0_1_776;
wire n_0_188;
wire n_0_1_0;
wire n_0_189;
wire n_0_1_1;
wire n_0_1_2;
wire n_0_190;
wire n_0_1_3;
wire n_0_191;
wire n_0_1_4;
wire n_0_192;
wire n_0_1_5;
wire n_0_193;
wire n_0_1_6;
wire n_0_194;
wire n_0_1_7;
wire n_0_195;
wire n_0_1_8;
wire n_0_196;
wire n_0_1_9;
wire n_0_197;
wire n_0_1_10;
wire n_0_198;
wire n_0_1_11;
wire n_0_199;
wire n_0_1_12;
wire n_0_200;
wire n_0_1_13;
wire n_0_201;
wire n_0_1_14;
wire n_0_202;
wire n_0_1_15;
wire n_0_203;
wire n_0_1_16;
wire n_0_1_17;
wire n_0_204;
wire n_0_1_18;
wire n_0_1_19;
wire n_0_205;
wire n_0_1_20;
wire n_0_1_21;
wire n_0_206;
wire n_0_1_22;
wire n_0_1_23;
wire n_0_207;
wire n_0_1_24;
wire n_0_1_25;
wire n_0_208;
wire n_0_1_26;
wire n_0_1_27;
wire n_0_209;
wire n_0_1_28;
wire n_0_1_29;
wire n_0_210;
wire n_0_1_30;
wire n_0_1_31;
wire n_0_211;
wire n_0_1_32;
wire n_0_1_33;
wire n_0_212;
wire n_0_1_34;
wire n_0_1_35;
wire n_0_213;
wire n_0_1_36;
wire n_0_1_37;
wire n_0_214;
wire n_0_1_38;
wire n_0_1_39;
wire n_0_215;
wire n_0_1_40;
wire n_0_1_41;
wire n_0_216;
wire n_0_1_42;
wire n_0_1_43;
wire n_0_217;
wire n_0_1_44;
wire n_0_1_45;
wire n_0_218;
wire n_0_1_46;
wire n_0_219;
wire n_0_1_47;
wire n_0_220;
wire n_0_1_48;
wire n_0_1_49;
wire n_0_221;
wire n_0_1_50;
wire n_0_1_51;
wire n_0_222;
wire n_0_1_52;
wire n_0_1_53;
wire n_0_223;
wire n_0_1_54;
wire n_0_1_55;
wire n_0_224;
wire n_0_1_56;
wire n_0_1_57;
wire n_0_225;
wire n_0_1_58;
wire n_0_1_59;
wire n_0_226;
wire n_0_1_60;
wire n_0_1_61;
wire n_0_227;
wire n_0_1_62;
wire n_0_1_63;
wire n_0_228;
wire n_0_1_64;
wire n_0_1_65;
wire n_0_229;
wire n_0_1_66;
wire n_0_1_67;
wire n_0_230;
wire n_0_1_68;
wire n_0_1_69;
wire n_0_231;
wire n_0_1_70;
wire n_0_1_71;
wire n_0_232;
wire n_0_1_72;
wire n_0_1_73;
wire n_0_233;
wire n_0_1_78;
wire n_0_1_83;
wire n_0_234;
wire n_0_1_84;
wire n_0_235;
wire n_0_1_85;
wire n_0_236;
wire n_0_1_86;
wire n_0_237;
wire n_0_1_87;
wire n_0_238;
wire n_0_1_88;
wire n_0_1_89;
wire n_0_239;
wire n_0_1_554;
wire n_0_1_555;
wire n_0_240;
wire n_0_1_589;
wire n_0_1_597;
wire n_0_241;
wire n_0_1_636;
wire n_0_1_640;
wire n_0_242;
wire n_0_1_679;
wire n_0_1_702;
wire n_0_243;
wire n_0_1_714;
wire n_0_244;
wire sgo__sro_n1290;
wire n_0_245;
wire n_0_1_723;
wire n_0_246;
wire n_0_1_724;
wire sgo__sro_n1194;
wire n_0_247;
wire n_0_1_727;
wire n_0_248;
wire n_0_1_749;
wire n_0_249;
wire n_0_1_752;
wire n_0_1_753;
wire n_0_250;
wire n_0_1_754;
wire n_0_1_755;
wire n_0_1_767;
wire n_0_1_769;
wire sgo__n779;
wire spw__n7739;
wire sgo__sro_n770;
wire slo__n3230;
wire n_0_1_838;
wire n_0_1_869;
wire n_0_1_870;
wire n_0_1_871;
wire n_0_1_872;
wire n_0_1_873;
wire n_0_1_874;
wire n_0_1_875;
wire n_0_1_876;
wire n_0_1_877;
wire n_0_1_878;
wire n_0_1_879;
wire n_0_1_880;
wire n_0_1_881;
wire n_0_1_882;
wire n_0_1_883;
wire n_0_1_884;
wire n_0_1_885;
wire n_0_1_886;
wire n_0_1_887;
wire n_0_1_888;
wire n_0_1_889;
wire n_0_1_890;
wire n_0_1_891;
wire n_0_1_892;
wire sgo__n874;
wire n_0_1_894;
wire sgo__sro_n741;
wire sgo__n850;
wire n_0_1_897;
wire n_0_1_898;
wire n_0_1_899;
wire n_0_1_900;
wire n_0_1_901;
wire n_0_1_902;
wire n_0_1_903;
wire n_0_1_904;
wire n_0_1_905;
wire n_0_1_906;
wire n_0_1_907;
wire n_0_1_908;
wire n_0_1_909;
wire n_0_283;
wire n_0_1_910;
wire n_0_677;
wire n_0_1_911;
wire n_0_1_912;
wire n_0_678;
wire n_0_1_913;
wire n_0_1_559;
wire n_0_1_914;
wire n_0_1_558;
wire n_0_1_557;
wire n_0_1_915;
wire slo__n3617;
wire n_0_702;
wire n_0_1_916;
wire n_0_1_917;
wire n_0_710;
wire n_0_1_918;
wire n_0_1_600;
wire n_0_1_919;
wire spw__n7776;
wire n_0_1_920;
wire n_0_1_599;
wire slo__n1550;
wire n_0_739;
wire n_0_1_922;
wire n_0_1_923;
wire n_0_743;
wire n_0_1_924;
wire n_0_1_642;
wire n_0_1_643;
wire n_0_1_925;
wire n_0_1_645;
wire n_0_1_926;
wire n_0_1_644;
wire n_0_772;
wire n_0_1_927;
wire n_0_1_688;
wire n_0_1_928;
wire n_0_1_687;
wire n_0_1_686;
wire n_0_1_929;
wire n_0_1_930;
wire n_0_785;
wire n_0_1_931;
wire n_0_1_786;
wire n_0_1_932;
wire n_0_797;
wire n_0_1_933;
wire n_0_1_810;
wire n_0_1_934;
wire n_0_801;
wire n_0_1_935;
wire n_0_1_818;
wire n_0_1_936;
wire n_0_806;
wire n_0_1_937;
wire n_0_1_938;
wire sgo__n1325;
wire n_0_1_939;
wire n_0_1_830;
wire n_0_1_940;
wire n_0_809;
wire slo__n1788;
wire n_0_1_942;
wire n_0_810;
wire n_0_1_943;
wire n_0_1_731;
wire n_0_1_944;
wire n_0_1_945;
wire n_0_1_729;
wire n_0_1_836;
wire n_0_1_946;
wire n_0_1_730;
wire n_0_1_947;
wire n_0_1_728;
wire n_0_1_948;
wire n_0_813;
wire n_0_1_949;
wire n_0_823;
wire n_0_1_950;
wire n_0_1_796;
wire n_0_826;
wire n_0_1_951;
wire opt_ipo_n5151;
wire n_0_827;
wire n_0_1_952;
wire n_0_1_804;
wire spw__n7729;
wire n_0_1_953;
wire n_0_1_806;
wire n_0_829;
wire n_0_1_954;
wire n_0_841;
wire n_0_1_955;
wire n_0_1_770;
wire n_0_843;
wire n_0_1_956;
wire n_0_1_771;
wire n_0_1_957;
wire n_0_844;
wire n_0_1_958;
wire n_0_1_959;
wire n_0_1_772;
wire sgo__n681;
wire n_0_1_775;
wire n_0_1_961;
wire n_0_1_962;
wire n_0_1_963;
wire n_0_1_964;
wire n_0_1_965;
wire n_0_1_966;
wire n_0_1_778;
wire n_0_1_967;
wire n_0_1_968;
wire n_0_1_969;
wire n_0_1_808;
wire n_0_1_826;
wire n_0_1_828;
wire n_0_1_832;
wire slo__n4931;
wire n_0_1_970;
wire n_0_251;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_255;
wire n_0_256;
wire n_0_257;
wire n_0_258;
wire n_0_259;
wire n_0_260;
wire n_0_261;
wire n_0_262;
wire n_0_263;
wire n_0_264;
wire n_0_265;
wire n_0_266;
wire n_0_267;
wire n_0_268;
wire n_0_269;
wire n_0_270;
wire n_0_271;
wire n_0_272;
wire n_0_273;
wire n_0_274;
wire n_0_275;
wire n_0_276;
wire n_0_277;
wire n_0_278;
wire n_0_279;
wire n_0_280;
wire n_0_281;
wire n_0_282;
wire n_0_284;
wire n_0_285;
wire n_0_286;
wire n_0_287;
wire n_0_288;
wire n_0_289;
wire n_0_290;
wire n_0_291;
wire n_0_292;
wire n_0_293;
wire n_0_294;
wire n_0_295;
wire n_0_296;
wire n_0_297;
wire n_0_298;
wire n_0_299;
wire n_0_300;
wire n_0_301;
wire n_0_302;
wire n_0_303;
wire n_0_304;
wire n_0_305;
wire n_0_306;
wire n_0_307;
wire n_0_308;
wire n_0_309;
wire n_0_310;
wire n_0_311;
wire n_0_312;
wire n_0_313;
wire n_0_314;
wire n_0_315;
wire n_0_316;
wire hfn_ipo_n43;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire uc_28;
wire uc_29;
wire uc_30;
wire uc_31;
wire uc_32;
wire uc_33;
wire uc_34;
wire uc_35;
wire uc_36;
wire uc_37;
wire uc_38;
wire uc_39;
wire uc_40;
wire uc_41;
wire uc_42;
wire uc_43;
wire uc_44;
wire uc_45;
wire uc_46;
wire uc_47;
wire uc_48;
wire uc_49;
wire uc_50;
wire uc_51;
wire uc_52;
wire uc_53;
wire uc_54;
wire uc_55;
wire uc_56;
wire uc_57;
wire uc_58;
wire uc_59;
wire uc_60;
wire uc_61;
wire uc_62;
wire uc_63;
wire uc_64;
wire uc_65;
wire uc_66;
wire uc_67;
wire uc_68;
wire uc_69;
wire uc_70;
wire uc_71;
wire uc_72;
wire uc_73;
wire uc_74;
wire uc_75;
wire uc_76;
wire uc_77;
wire uc_78;
wire uc_79;
wire uc_80;
wire uc_81;
wire uc_82;
wire uc_83;
wire uc_84;
wire uc_85;
wire uc_86;
wire uc_87;
wire uc_88;
wire uc_89;
wire uc_90;
wire uc_91;
wire uc_92;
wire uc_93;
wire uc_94;
wire uc_95;
wire uc_96;
wire uc_97;
wire uc_98;
wire uc_99;
wire uc_100;
wire uc_101;
wire uc_102;
wire uc_103;
wire uc_104;
wire uc_105;
wire uc_106;
wire uc_107;
wire uc_108;
wire uc_109;
wire uc_110;
wire uc_111;
wire uc_112;
wire uc_113;
wire uc_114;
wire uc_115;
wire uc_116;
wire uc_117;
wire uc_118;
wire uc_119;
wire uc_120;
wire uc_121;
wire uc_122;
wire uc_123;
wire uc_124;
wire uc_125;
wire uc_126;
wire uc_127;
wire uc_128;
wire uc_129;
wire uc_130;
wire uc_131;
wire uc_132;
wire uc_133;
wire uc_134;
wire uc_135;
wire uc_136;
wire uc_137;
wire uc_138;
wire uc_139;
wire uc_140;
wire uc_141;
wire uc_142;
wire uc_143;
wire uc_144;
wire uc_145;
wire uc_146;
wire uc_147;
wire uc_148;
wire uc_149;
wire uc_150;
wire uc_151;
wire uc_152;
wire uc_153;
wire uc_154;
wire uc_155;
wire uc_156;
wire uc_157;
wire uc_158;
wire uc_159;
wire uc_160;
wire uc_161;
wire uc_162;
wire uc_163;
wire uc_164;
wire uc_165;
wire uc_166;
wire uc_167;
wire uc_168;
wire uc_169;
wire uc_170;
wire uc_171;
wire uc_172;
wire uc_173;
wire uc_174;
wire uc_175;
wire uc_176;
wire uc_177;
wire uc_178;
wire uc_179;
wire uc_180;
wire uc_181;
wire uc_182;
wire uc_183;
wire uc_184;
wire uc_185;
wire uc_186;
wire uc_187;
wire uc_188;
wire uc_189;
wire uc_190;
wire uc_191;
wire uc_192;
wire uc_193;
wire uc_194;
wire uc_195;
wire uc_196;
wire uc_197;
wire uc_198;
wire uc_199;
wire uc_200;
wire uc_201;
wire uc_202;
wire uc_203;
wire uc_204;
wire uc_205;
wire uc_206;
wire uc_207;
wire uc_208;
wire uc_209;
wire uc_210;
wire uc_211;
wire uc_212;
wire uc_213;
wire uc_214;
wire uc_215;
wire uc_216;
wire uc_217;
wire uc_218;
wire uc_219;
wire uc_220;
wire uc_221;
wire uc_222;
wire uc_223;
wire uc_224;
wire uc_225;
wire uc_226;
wire uc_227;
wire uc_228;
wire uc_229;
wire uc_230;
wire uc_231;
wire uc_232;
wire uc_233;
wire uc_234;
wire uc_235;
wire uc_236;
wire uc_237;
wire uc_238;
wire uc_239;
wire uc_240;
wire uc_241;
wire uc_242;
wire uc_243;
wire uc_244;
wire uc_245;
wire uc_246;
wire uc_247;
wire uc_248;
wire uc_249;
wire uc_250;
wire uc_251;
wire uc_252;
wire uc_253;
wire uc_254;
wire uc_255;
wire uc_256;
wire uc_257;
wire uc_258;
wire uc_259;
wire uc_260;
wire uc_261;
wire uc_262;
wire uc_263;
wire uc_264;
wire uc_265;
wire uc_266;
wire uc_267;
wire uc_268;
wire uc_269;
wire uc_270;
wire uc_271;
wire uc_272;
wire uc_273;
wire uc_274;
wire uc_275;
wire uc_276;
wire uc_277;
wire uc_278;
wire uc_279;
wire uc_280;
wire uc_281;
wire uc_282;
wire uc_283;
wire uc_284;
wire uc_285;
wire uc_286;
wire uc_287;
wire uc_288;
wire uc_289;
wire uc_290;
wire uc_291;
wire uc_292;
wire uc_293;
wire uc_294;
wire uc_295;
wire uc_296;
wire uc_297;
wire uc_298;
wire uc_299;
wire uc_300;
wire uc_301;
wire uc_302;
wire uc_303;
wire uc_304;
wire uc_305;
wire uc_306;
wire uc_307;
wire uc_308;
wire uc_309;
wire uc_310;
wire uc_311;
wire uc_312;
wire uc_313;
wire uc_314;
wire uc_315;
wire uc_316;
wire uc_317;
wire uc_318;
wire uc_319;
wire uc_320;
wire uc_321;
wire uc_322;
wire uc_323;
wire uc_324;
wire uc_325;
wire uc_326;
wire uc_327;
wire uc_328;
wire uc_329;
wire uc_330;
wire uc_331;
wire uc_332;
wire uc_333;
wire uc_334;
wire uc_335;
wire uc_336;
wire uc_337;
wire uc_338;
wire uc_339;
wire uc_340;
wire uc_341;
wire uc_342;
wire uc_343;
wire uc_344;
wire uc_345;
wire uc_346;
wire uc_347;
wire uc_348;
wire uc_349;
wire uc_350;
wire uc_351;
wire uc_352;
wire uc_353;
wire uc_354;
wire uc_355;
wire uc_356;
wire uc_357;
wire uc_358;
wire uc_359;
wire uc_360;
wire uc_361;
wire uc_362;
wire uc_363;
wire uc_364;
wire uc_365;
wire uc_366;
wire uc_367;
wire uc_368;
wire uc_369;
wire uc_370;
wire uc_371;
wire uc_372;
wire uc_373;
wire uc_374;
wire uc_375;
wire uc_376;
wire uc_377;
wire uc_378;
wire uc_379;
wire uc_380;
wire uc_381;
wire uc_382;
wire uc_383;
wire uc_384;
wire uc_385;
wire uc_386;
wire uc_387;
wire uc_388;
wire uc_389;
wire uc_390;
wire uc_391;
wire uc_392;
wire uc_393;
wire uc_394;
wire uc_395;
wire uc_396;
wire uc_397;
wire uc_398;
wire uc_399;
wire uc_400;
wire uc_401;
wire uc_402;
wire uc_403;
wire uc_404;
wire uc_405;
wire uc_406;
wire uc_407;
wire uc_408;
wire uc_409;
wire uc_410;
wire uc_411;
wire uc_412;
wire uc_413;
wire uc_414;
wire uc_415;
wire uc_416;
wire uc_417;
wire uc_418;
wire uc_419;
wire uc_420;
wire uc_421;
wire uc_422;
wire uc_423;
wire uc_424;
wire uc_425;
wire uc_426;
wire uc_427;
wire uc_428;
wire uc_429;
wire uc_430;
wire uc_431;
wire uc_432;
wire uc_433;
wire uc_434;
wire uc_435;
wire uc_436;
wire uc_437;
wire uc_438;
wire uc_439;
wire uc_440;
wire uc_441;
wire uc_442;
wire uc_443;
wire uc_444;
wire uc_445;
wire uc_446;
wire uc_447;
wire uc_448;
wire uc_449;
wire uc_450;
wire uc_451;
wire uc_452;
wire uc_453;
wire uc_454;
wire uc_455;
wire uc_456;
wire uc_457;
wire uc_458;
wire uc_459;
wire uc_460;
wire uc_461;
wire uc_462;
wire uc_463;
wire uc_464;
wire uc_465;
wire uc_466;
wire uc_467;
wire uc_468;
wire uc_469;
wire uc_470;
wire uc_471;
wire uc_472;
wire uc_473;
wire uc_474;
wire uc_475;
wire uc_476;
wire uc_477;
wire uc_478;
wire uc_479;
wire uc_480;
wire uc_481;
wire uc_482;
wire uc_483;
wire uc_484;
wire uc_485;
wire uc_486;
wire uc_487;
wire uc_488;
wire uc_489;
wire uc_490;
wire uc_491;
wire uc_492;
wire uc_493;
wire uc_494;
wire uc_495;
wire uc_496;
wire uc_497;
wire uc_498;
wire uc_499;
wire uc_500;
wire uc_501;
wire uc_502;
wire uc_503;
wire drc_ipo_n58;
wire hfn_ipo_n41;
wire opt_ipo_n5135;
wire drc_ipo_n52;
wire slo__xsl_n4224;
wire drc_ipo_n50;
wire drc_ipo_n59;
wire drc_ipo_n56;
wire sph__n7809;
wire drc_ipo_n54;
wire drc_ipo_n53;
wire drc_ipo_n48;
wire sgo__n678;
wire hfn_ipo_n46;
wire sgo__n731;
wire sgo__n734;
wire sgo__sro_n769;
wire CLOCK_slo__sro_n6809;
wire sgo__sro_n697;
wire sgo__n895;
wire sgo__sro_n702;
wire sgo__sro_n703;
wire sgo__sro_n704;
wire sgo__sro_n705;
wire sgo__sro_n739;
wire CLOCK_slh__n7179;
wire sgo__sro_n719;
wire sgo__sro_n720;
wire CLOCK_slh__n7200;
wire sgo__sro_n722;
wire sgo__sro_n771;
wire sgo__sro_n772;
wire sgo__n759;
wire sgo__n847;
wire opt_ipo_n5506;
wire sgo__sro_n799;
wire sgo__sro_n800;
wire sgo__sro_n801;
wire sgo__n839;
wire sgo__sro_n809;
wire sgo__n962;
wire sgo__sro_n811;
wire sgo__n877;
wire sgo__n880;
wire sgo__n943;
wire spw__n7777;
wire opt_ipo_n5145;
wire sgo__sro_n905;
wire sgo__sro_n906;
wire sgo__sro_n907;
wire sgo__sro_n908;
wire sgo__sro_n909;
wire opt_ipo_n5165;
wire sgo__n959;
wire sgo__n1009;
wire sgo__sro_n1195;
wire sgo__n1043;
wire CLOCK_slh__n7195;
wire sgo__n1053;
wire sgo__n1056;
wire sgo__sro_n1197;
wire sgo__n1116;
wire opt_ipo_n5682;
wire sgo__sro_n1208;
wire sgo__sro_n1209;
wire sgo__sro_n1210;
wire sgo__n1238;
wire sgo__n1241;
wire sgo__n1251;
wire sgo__n1223;
wire sgo__n1324;
wire spw__n7730;
wire sgo__sro_n1289;
wire CLOCK_slo__mro_n6730;
wire sgo__sro_n1270;
wire sgo__sro_n1272;
wire sgo__sro_n1273;
wire slo___n2464;
wire sgo__n1339;
wire CLOCK_slh__n7202;
wire opt_ipo_n5795;
wire opt_ipo_n5785;
wire slo__xsl_n1366;
wire slo__xsl_n1367;
wire slo__n1376;
wire slo__n1475;
wire slo__n3378;
wire slo__sro_n1458;
wire slo__xsl_n1425;
wire slo__xsl_n1426;
wire slo__n1402;
wire slo__sro_n1459;
wire slo__n1493;
wire slo__n1559;
wire slo__n1580;
wire slo__n1581;
wire slo__n1588;
wire slo__sro_n1594;
wire slo__sro_n1595;
wire slo__sro_n1596;
wire slo__sro_n1605;
wire slo__sro_n1606;
wire slo__sro_n1607;
wire slo__sro_n1608;
wire slo__sro_n1622;
wire slo__sro_n1623;
wire slo__n1627;
wire slo__n1649;
wire slo__xsl_n1694;
wire slo__xsl_n1641;
wire slo__xsl_n1642;
wire slo__xsl_n1695;
wire slo__n1702;
wire slo__xsl_n1669;
wire slo__xsl_n1670;
wire slo__sro_n1746;
wire slo__sro_n1747;
wire CLOCK_slh__n7160;
wire slo__sro_n1748;
wire slo__xsl_n1736;
wire slo__xsl_n1737;
wire slo__sro_n1749;
wire slo__n1762;
wire slo__n1801;
wire slo__xsl_n1889;
wire slo__xsl_n1890;
wire slo__n1812;
wire slo__n1828;
wire slo__n1897;
wire slo__mro_n1860;
wire slo__mro_n1861;
wire slo__sro_n1908;
wire slo__n1936;
wire slo__xsl_n1963;
wire slo__xsl_n1964;
wire CLOCK_slh__n7206;
wire CLOCK_slh__n7207;
wire opt_ipo_n5774;
wire slo__xsl_n2010;
wire slo__xsl_n2011;
wire slo__n2069;
wire slo__mro_n2075;
wire slo__sro_n2080;
wire CLOCK_slh__n7196;
wire opt_ipo_n5164;
wire spw__n7778;
wire slo__sro_n2149;
wire slo__sro_n2150;
wire CLOCK_slo__mro_n6799;
wire slo__n2216;
wire slo__n2235;
wire slo___n2244;
wire slo___n2245;
wire slo__n2232;
wire CLOCK_slo__sro_n6735;
wire slo___n2247;
wire slo___n2248;
wire slo__sro_n2333;
wire opt_ipo_n5191;
wire slo__n2517;
wire opt_ipo_n5672;
wire slo__n2528;
wire slo__n2400;
wire slo__n2915;
wire slo__n2805;
wire CLOCK_slo__sro_n6740;
wire slo__n2762;
wire slo__sro_n2570;
wire CLOCK_slh__n7168;
wire slo__n2712;
wire slo__n2871;
wire CLOCK_slh__n7190;
wire slo__n2969;
wire slo__sro_n2992;
wire slo__n2885;
wire slo__n3030;
wire slo__sro_n2959;
wire CLOCK_slh__n7158;
wire opt_ipo_n5710;
wire opt_ipo_n5712;
wire spw__n7741;
wire slo___n3116;
wire slo__n3016;
wire slo__sro_n3170;
wire slo__sro_n3243;
wire slo__sro_n3317;
wire slo__n3307;
wire slo__n3134;
wire slo__n3345;
wire slo__n3204;
wire slo__sro_n3369;
wire slo__sro_n3370;
wire CLOCK_slh__n7159;
wire slo__n3399;
wire slo__n3402;
wire slo__sro_n3406;
wire slo__sro_n3407;
wire opt_ipo_n5664;
wire CLOCK_slo__sro_n6736;
wire CLOCK_slo__sro_n6734;
wire slo___n3458;
wire opt_ipo_n5711;
wire slo___n3489;
wire opt_ipo_n5686;
wire opt_ipo_n5103;
wire CTS_n_tid1_5915;
wire opt_ipo_n5107;
wire opt_ipo_n5108;
wire slo___n3496;
wire CLOCK_sgo__n6410;
wire slo__n3547;
wire slo__n3614;
wire slo__n3522;
wire slo__sro_n3675;
wire slo__n3595;
wire slo__sro_n3584;
wire slo__n3691;
wire opt_ipo_n5195;
wire slo__n3640;
wire slo__sro_n3685;
wire slo__n3760;
wire opt_ipo_n5719;
wire opt_ipo_n5702;
wire slo__sro_n3808;
wire opt_ipo_n5125;
wire CLOCK_slh__n7194;
wire slo__sro_n3734;
wire slo__sro_n3735;
wire slo__sro_n3736;
wire slo__n3799;
wire CLOCK_sgo__n6468;
wire slo__n3910;
wire slo__sro_n4174;
wire CLOCK_spw__n7299;
wire slo__n3840;
wire slo__xsl_n3900;
wire slo__xsl_n3901;
wire slo__sro_n4175;
wire slo__sro_n4176;
wire CLOCK_slh__n7201;
wire slo__xsl_n4223;
wire slo__n4197;
wire opt_ipo_n5196;
wire slo__xsl_n4322;
wire spw__n7686;
wire slo__xsl_n4323;
wire CLOCK_spw__n7322;
wire opt_ipo_n5152;
wire CLOCK_spw__n7329;
wire slo__xsl_n4785;
wire slo__xsl_n4487;
wire slo__xsl_n4488;
wire slo__xsl_n4786;
wire opt_ipo_n5197;
wire slo__n4849;
wire opt_ipo_n5198;
wire CLOCK_opt_ipo_n5880;
wire opt_ipo_n5204;
wire opt_ipo_n5205;
wire CLOCK_spw__n7344;
wire opt_ipo_n5208;
wire opt_ipo_n5209;
wire CLOCK_slh__n7180;
wire opt_ipo_n5223;
wire opt_ipo_n5224;
wire opt_ipo_n5230;
wire CLOCK_spw__n7303;
wire opt_ipo_n5258;
wire opt_ipo_n5278;
wire opt_ipo_n5280;
wire opt_ipo_n5285;
wire CLOCK_spw__n7320;
wire CLOCK_slo__sro_n6741;
wire CLOCK_slh__n7170;
wire opt_ipo_n5297;
wire CLOCK_slh__n7188;
wire CLOCK_spw__n7291;
wire opt_ipo_n5303;
wire opt_ipo_n5307;
wire opt_ipo_n5311;
wire opt_ipo_n5312;
wire opt_ipo_n5314;
wire opt_ipo_n5315;
wire CLOCK_spw__n7321;
wire opt_ipo_n5332;
wire opt_ipo_n5339;
wire opt_ipo_n5358;
wire opt_ipo_n5362;
wire CLOCK_spw__n7292;
wire opt_ipo_n5373;
wire opt_ipo_n5374;
wire opt_ipo_n5385;
wire opt_ipo_n5393;
wire opt_ipo_n5395;
wire opt_ipo_n5398;
wire opt_ipo_n5411;
wire opt_ipo_n5415;
wire opt_ipo_n5416;
wire opt_ipo_n5417;
wire opt_ipo_n5419;
wire opt_ipo_n5423;
wire opt_ipo_n5433;
wire opt_ipo_n5438;
wire CLOCK_slh__n7178;
wire opt_ipo_n5459;
wire opt_ipo_n5465;
wire opt_ipo_n5466;


BUF_X16 hfn_ipo_c43 (.Z (hfn_ipo_n43), .A (n_0_1_752));
BUF_X4 sgo__c894 (.Z (sgo__n895), .A (\A_imm_2s_complement[15] ));
NAND2_X4 i_0_1_1658 (.ZN (n_0_316), .A1 (CTS_n_tid1_5915), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1657 (.ZN (n_0_315), .A1 (A[31]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1656 (.ZN (n_0_314), .A1 (A[30]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1655 (.ZN (n_0_313), .A1 (A[29]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1654 (.ZN (n_0_312), .A1 (A[28]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1653 (.ZN (n_0_311), .A1 (A[27]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1652 (.ZN (n_0_310), .A1 (A[26]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1651 (.ZN (n_0_309), .A1 (A[25]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1650 (.ZN (n_0_308), .A1 (A[24]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1649 (.ZN (n_0_307), .A1 (A[23]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1648 (.ZN (n_0_306), .A1 (A[22]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1647 (.ZN (n_0_305), .A1 (A[21]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1646 (.ZN (n_0_304), .A1 (A[20]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1645 (.ZN (n_0_303), .A1 (A[19]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1644 (.ZN (n_0_302), .A1 (A[18]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1643 (.ZN (n_0_301), .A1 (A[17]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1642 (.ZN (n_0_300), .A1 (A[16]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1641 (.ZN (n_0_299), .A1 (A[15]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1640 (.ZN (n_0_298), .A1 (A[14]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1639 (.ZN (n_0_297), .A1 (A[13]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1638 (.ZN (n_0_296), .A1 (A[12]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1637 (.ZN (n_0_295), .A1 (A[11]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1636 (.ZN (n_0_294), .A1 (A[10]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1635 (.ZN (n_0_293), .A1 (A[9]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1634 (.ZN (n_0_292), .A1 (A[8]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1633 (.ZN (n_0_291), .A1 (A[7]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1632 (.ZN (n_0_290), .A1 (A[6]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1631 (.ZN (n_0_289), .A1 (A[5]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1630 (.ZN (n_0_288), .A1 (A[4]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1629 (.ZN (n_0_287), .A1 (A[3]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1628 (.ZN (n_0_286), .A1 (A[2]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1627 (.ZN (n_0_285), .A1 (A[1]), .A2 (hfn_ipo_n45));
AND2_X1 i_0_1_1626 (.ZN (n_0_284), .A1 (A[0]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1625 (.ZN (n_0_282), .A1 (B[31]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1624 (.ZN (n_0_281), .A1 (B[30]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1623 (.ZN (n_0_280), .A1 (B[29]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1622 (.ZN (n_0_279), .A1 (B[28]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1621 (.ZN (n_0_278), .A1 (B[27]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1620 (.ZN (n_0_277), .A1 (B[26]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1619 (.ZN (n_0_276), .A1 (B[25]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1618 (.ZN (n_0_275), .A1 (B[24]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1617 (.ZN (n_0_274), .A1 (B[23]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1616 (.ZN (n_0_273), .A1 (B[22]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1615 (.ZN (n_0_272), .A1 (B[21]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1614 (.ZN (n_0_271), .A1 (B[20]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1613 (.ZN (n_0_270), .A1 (B[19]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1612 (.ZN (n_0_269), .A1 (B[18]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1611 (.ZN (n_0_268), .A1 (B[17]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1610 (.ZN (n_0_267), .A1 (B[16]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1609 (.ZN (n_0_266), .A1 (B[15]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1608 (.ZN (n_0_265), .A1 (B[14]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1607 (.ZN (n_0_264), .A1 (B[13]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1606 (.ZN (n_0_263), .A1 (B[12]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1605 (.ZN (n_0_262), .A1 (B[11]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1604 (.ZN (n_0_261), .A1 (B[10]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1603 (.ZN (n_0_260), .A1 (B[9]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1602 (.ZN (n_0_259), .A1 (B[8]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1601 (.ZN (n_0_258), .A1 (B[7]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1600 (.ZN (n_0_257), .A1 (B[6]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1599 (.ZN (n_0_256), .A1 (B[5]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1598 (.ZN (n_0_255), .A1 (B[4]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1597 (.ZN (n_0_254), .A1 (B[3]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1596 (.ZN (n_0_253), .A1 (B[2]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1595 (.ZN (n_0_252), .A1 (B[1]), .A2 (hfn_ipo_n46));
AND2_X1 i_0_1_1594 (.ZN (n_0_251), .A1 (B[0]), .A2 (hfn_ipo_n46));
INV_X1 i_0_1_1593 (.ZN (n_0_1_970), .A (reset));
AOI21_X4 i_0_1_1592 (.ZN (slo__n4849), .A (n_0_1_835), .B1 (n_0_29), .B2 (A_in));
INV_X8 i_0_1_1591 (.ZN (\A_imm[30] ), .A (sgo__n734));
AOI21_X2 i_0_1_1590 (.ZN (n_0_1_832), .A (n_0_1_833), .B1 (n_0_28), .B2 (A_in));
INV_X8 i_0_1_1589 (.ZN (\A_imm[29] ), .A (n_0_1_832));
AOI21_X2 i_0_1_1588 (.ZN (n_0_1_828), .A (n_0_1_829), .B1 (n_0_26), .B2 (hfn_ipo_n41));
INV_X8 i_0_1_1587 (.ZN (\A_imm[27] ), .A (n_0_1_828));
AOI21_X2 i_0_1_1586 (.ZN (n_0_1_826), .A (n_0_1_827), .B1 (n_0_25), .B2 (hfn_ipo_n41));
INV_X4 opt_ipo_c6238 (.ZN (opt_ipo_n5683), .A (n_0_1_693));
AOI21_X1 i_0_1_1582 (.ZN (n_0_1_808), .A (n_0_1_809), .B1 (n_0_16), .B2 (hfn_ipo_n41));
CLKBUF_X1 sph__c8607 (.Z (sph__n7809), .A (sph__n7808));
INV_X2 i_0_1_1580 (.ZN (n_0_1_969), .A (A_in));
NOR2_X1 i_0_1_1579 (.ZN (n_0_1_968), .A1 (n_0_4), .A2 (n_0_1_969));
CLKBUF_X2 slo__c3697 (.Z (slo__n3378), .A (slo__sro_n3368));
NOR2_X1 i_0_1_1577 (.ZN (n_0_1_967), .A1 (A_in), .A2 (n_0_1_839));
AOI21_X4 i_0_1_1576 (.ZN (n_0_1_778), .A (n_0_1_967), .B1 (n_0_1), .B2 (A_in));
INV_X4 i_0_1_1575 (.ZN (\A_imm[2] ), .A (n_0_1_778));
INV_X1 i_0_1_1574 (.ZN (n_0_1_966), .A (n_0_0));
NAND2_X1 i_0_1_1573 (.ZN (n_0_1_965), .A1 (n_0_1_969), .A2 (n_0_154));
OAI21_X2 i_0_1_1572 (.ZN (\A_imm[1] ), .A (n_0_1_965), .B1 (n_0_1_966), .B2 (n_0_1_969));
INV_X1 i_0_1_1571 (.ZN (n_0_1_964), .A (\A_imm_2s_complement[31] ));
INV_X1 i_0_1_1570 (.ZN (n_0_1_963), .A (drc_ipo_n58));
INV_X1 i_0_1_1569 (.ZN (n_0_1_962), .A (n_0_31));
NAND2_X1 i_0_1_1568 (.ZN (n_0_1_961), .A1 (n_0_1_963), .A2 (n_0_185));
OAI21_X1 i_0_1_1567 (.ZN (n_0_1_775), .A (n_0_1_961), .B1 (n_0_1_962), .B2 (n_0_1_963));
BUF_X4 opt_ipo_c5735 (.Z (opt_ipo_n5151), .A (n_0_1_920));
NAND2_X4 i_0_1_1565 (.ZN (n_0_1_772), .A1 (n_0_1_774), .A2 (n_0_186));
INV_X1 i_0_1_1564 (.ZN (n_0_1_959), .A (n_0_1_772));
NAND3_X1 i_0_1_1563 (.ZN (n_0_1_958), .A1 (n_0_30), .A2 (A_in), .A3 (n_0_1_959));
OAI21_X1 i_0_1_1562 (.ZN (n_0_844), .A (n_0_1_958), .B1 (n_0_1_964), .B2 (n_0_1_774));
NAND2_X1 i_0_1_1561 (.ZN (n_0_1_957), .A1 (n_0_1_775), .A2 (n_0_186));
NOR2_X4 i_0_1_1560 (.ZN (n_0_1_771), .A1 (n_0_1_774), .A2 (n_0_186));
NAND2_X1 i_0_1_1559 (.ZN (n_0_1_956), .A1 (\A_imm_2s_complement[30] ), .A2 (n_0_1_771));
OAI211_X1 i_0_1_1528 (.ZN (n_0_843), .A (n_0_1_958), .B (n_0_1_956), .C1 (n_0_1_964), .C2 (n_0_1_957));
INV_X2 i_0_1_1527 (.ZN (n_0_1_770), .A (n_0_1_957));
AOI22_X2 i_0_1_1526 (.ZN (n_0_1_955), .A1 (\A_imm_2s_complement[29] ), .A2 (n_0_1_770)
    , .B1 (\A_imm_2s_complement[28] ), .B2 (n_0_1_771));
OAI21_X2 i_0_1_1523 (.ZN (n_0_841), .A (n_0_1_955), .B1 (slo__xsl_n1736), .B2 (n_0_1_772));
AOI22_X1 i_0_1_1522 (.ZN (n_0_1_954), .A1 (opt_ipo_n5411), .A2 (n_0_1_770), .B1 (opt_ipo_n5162), .B2 (n_0_1_771));
OAI21_X1 i_0_1_1520 (.ZN (n_0_829), .A (n_0_1_954), .B1 (slo__xsl_n1366), .B2 (n_0_1_772));
AOI21_X2 i_0_1_1519 (.ZN (n_0_1_806), .A (n_0_1_807), .B1 (n_0_15), .B2 (hfn_ipo_n41));
AOI22_X1 i_0_1_1517 (.ZN (n_0_1_953), .A1 (opt_ipo_n5162), .A2 (n_0_1_770), .B1 (sgo__n895), .B2 (n_0_1_771));
BUF_X2 spw__L1_c8528 (.Z (spw__n7729), .A (opt_ipo_n5285));
AOI21_X1 i_0_1_1513 (.ZN (n_0_1_804), .A (n_0_1_805), .B1 (n_0_14), .B2 (hfn_ipo_n41));
AOI22_X1 i_0_1_1511 (.ZN (n_0_1_952), .A1 (sgo__n895), .A2 (n_0_1_770), .B1 (slo__n2107), .B2 (n_0_1_771));
OAI21_X1 i_0_1_1510 (.ZN (n_0_827), .A (n_0_1_952), .B1 (n_0_1_772), .B2 (slo__n1828));
AOI21_X4 i_0_1_1507 (.ZN (sgo__n681), .A (n_0_1_803), .B1 (n_0_13), .B2 (hfn_ipo_n41));
AOI22_X1 i_0_1_1499 (.ZN (n_0_1_951), .A1 (slo__n2107), .A2 (n_0_1_770), .B1 (opt_ipo_n5710), .B2 (n_0_1_771));
OAI21_X1 i_0_1_1495 (.ZN (n_0_826), .A (n_0_1_951), .B1 (n_0_1_772), .B2 (slo__xsl_n4487));
AOI21_X2 i_0_1_1487 (.ZN (n_0_1_796), .A (n_0_1_797), .B1 (n_0_10), .B2 (hfn_ipo_n41));
AOI22_X2 i_0_1_1484 (.ZN (n_0_1_950), .A1 (slo__n3026), .A2 (n_0_1_770), .B1 (opt_ipo_n5466), .B2 (n_0_1_771));
OAI21_X1 i_0_1_1483 (.ZN (n_0_823), .A (n_0_1_950), .B1 (n_0_1_772), .B2 (slo___n3458));
NAND2_X1 i_0_1_1481 (.ZN (n_0_1_949), .A1 (n_0_1_959), .A2 (opt_ipo_n5459));
NAND2_X1 i_0_1_1478 (.ZN (n_0_813), .A1 (n_0_1_739), .A2 (n_0_1_949));
OR3_X1 i_0_1_1475 (.ZN (n_0_1_948), .A1 (n_0_1_735), .A2 (n_0_1_738), .A3 (n_0_1_775));
INV_X4 i_0_1_1466 (.ZN (n_0_1_728), .A (n_0_1_948));
NAND2_X1 i_0_1_1451 (.ZN (n_0_1_947), .A1 (opt_ipo_n5358), .A2 (n_0_1_728));
NOR2_X4 i_0_1_1449 (.ZN (n_0_1_730), .A1 (n_0_1_737), .A2 (n_0_1_736));
NAND2_X1 i_0_1_1448 (.ZN (n_0_1_946), .A1 (\A_imm[30] ), .A2 (n_0_1_730));
NAND2_X4 i_0_1_1447 (.ZN (n_0_1_836), .A1 (n_0_30), .A2 (A_in));
NAND2_X4 i_0_1_1440 (.ZN (n_0_1_729), .A1 (n_0_1_732), .A2 (n_0_1_735));
OR2_X1 i_0_1_1439 (.ZN (n_0_1_945), .A1 (n_0_1_836), .A2 (n_0_1_729));
NAND2_X1 i_0_1_1438 (.ZN (n_0_1_944), .A1 (n_0_1_732), .A2 (n_0_1_736));
INV_X4 i_0_1_1437 (.ZN (n_0_1_731), .A (n_0_1_944));
NAND2_X1 i_0_1_1436 (.ZN (n_0_1_943), .A1 (sgo__n731), .A2 (n_0_1_731));
NAND4_X1 i_0_1_1435 (.ZN (n_0_810), .A1 (n_0_1_947), .A2 (n_0_1_943), .A3 (n_0_1_946), .A4 (n_0_1_945));
NAND2_X1 i_0_1_1434 (.ZN (n_0_1_942), .A1 (\A_imm_2s_complement[29] ), .A2 (n_0_1_728));
CLKBUF_X2 slo__c1989 (.Z (slo__n1788), .A (\A_imm[7] ));
OAI211_X1 i_0_1_1431 (.ZN (n_0_809), .A (slo__sro_n1746), .B (n_0_1_942), .C1 (sgo__n734), .C2 (n_0_1_729));
NAND2_X1 i_0_1_1430 (.ZN (n_0_1_940), .A1 (\A_imm_2s_complement[27] ), .A2 (n_0_1_728));
AOI21_X4 i_0_1_1429 (.ZN (n_0_1_830), .A (n_0_1_831), .B1 (n_0_27), .B2 (A_in));
AOI22_X1 i_0_1_1428 (.ZN (n_0_1_939), .A1 (\A_imm_2s_complement[28] ), .A2 (n_0_1_731)
    , .B1 (\A_imm[27] ), .B2 (n_0_1_730));
INV_X16 sgo__c1448 (.ZN (n_0_1_792), .A (sgo__n1325));
NAND2_X1 i_0_1_1426 (.ZN (n_0_1_938), .A1 (\A_imm_2s_complement[26] ), .A2 (n_0_1_728));
AOI22_X1 i_0_1_1423 (.ZN (n_0_1_937), .A1 (\A_imm_2s_complement[27] ), .A2 (n_0_1_731)
    , .B1 (slo__n1897), .B2 (n_0_1_730));
OAI211_X1 i_0_1_1422 (.ZN (n_0_806), .A (n_0_1_937), .B (n_0_1_938), .C1 (slo__n2762), .C2 (n_0_1_729));
NAND2_X1 i_0_1_1399 (.ZN (n_0_1_936), .A1 (\A_imm_2s_complement[21] ), .A2 (n_0_1_728));
AOI21_X4 i_0_1_1398 (.ZN (n_0_1_818), .A (n_0_1_819), .B1 (n_0_21), .B2 (hfn_ipo_n41));
AOI22_X1 i_0_1_1397 (.ZN (n_0_1_935), .A1 (\A_imm_2s_complement[22] ), .A2 (n_0_1_731)
    , .B1 (opt_ipo_n5135), .B2 (n_0_1_730));
OAI211_X1 i_0_1_1396 (.ZN (n_0_801), .A (n_0_1_935), .B (n_0_1_936), .C1 (n_0_1_729), .C2 (slo__xsl_n1641));
NAND2_X1 i_0_1_1395 (.ZN (n_0_1_934), .A1 (opt_ipo_n5411), .A2 (n_0_1_728));
AOI21_X4 i_0_1_1394 (.ZN (n_0_1_810), .A (n_0_1_811), .B1 (n_0_17), .B2 (hfn_ipo_n41));
AOI22_X1 i_0_1_1393 (.ZN (n_0_1_933), .A1 (\A_imm_2s_complement[18] ), .A2 (n_0_1_731)
    , .B1 (slo__n3402), .B2 (n_0_1_730));
OAI211_X1 i_0_1_1392 (.ZN (n_0_797), .A (n_0_1_933), .B (n_0_1_934), .C1 (n_0_1_729), .C2 (slo__xsl_n1425));
NAND2_X1 i_0_1_1387 (.ZN (n_0_1_932), .A1 (\A_imm_2s_complement[5] ), .A2 (n_0_1_728));
AOI21_X4 i_0_1_1386 (.ZN (n_0_1_786), .A (n_0_1_787), .B1 (n_0_5), .B2 (A_in));
AOI22_X1 i_0_1_1366 (.ZN (n_0_1_931), .A1 (opt_ipo_n5205), .A2 (n_0_1_731), .B1 (slo__n3378), .B2 (n_0_1_730));
OAI211_X1 i_0_1_1364 (.ZN (n_0_785), .A (n_0_1_931), .B (n_0_1_932), .C1 (n_0_1_729), .C2 (slo__xsl_n1694));
OR3_X2 i_0_1_1355 (.ZN (n_0_1_930), .A1 (opt_ipo_n5683), .A2 (n_0_1_695), .A3 (n_0_1_736));
NAND2_X1 i_0_1_1353 (.ZN (n_0_1_929), .A1 (\A_imm_2s_complement[25] ), .A2 (opt_ipo_n5278));
NAND2_X4 i_0_1_1352 (.ZN (n_0_1_686), .A1 (opt_ipo_n5683), .A2 (n_0_1_689));
NOR2_X4 i_0_1_1351 (.ZN (n_0_1_687), .A1 (n_0_1_693), .A2 (n_0_1_694));
NAND2_X1 i_0_1_1350 (.ZN (n_0_1_928), .A1 (n_0_1_693), .A2 (n_0_1_689));
INV_X2 i_0_1_1349 (.ZN (n_0_1_688), .A (n_0_1_928));
AOI22_X1 i_0_1_1348 (.ZN (n_0_1_927), .A1 (\A_imm_2s_complement[26] ), .A2 (opt_ipo_n5679)
    , .B1 (opt_ipo_n5362), .B2 (n_0_1_687));
OAI211_X1 i_0_1_1345 (.ZN (n_0_772), .A (n_0_1_927), .B (n_0_1_929), .C1 (slo__xsl_n1889), .C2 (n_0_1_686));
NOR2_X4 i_0_1_1344 (.ZN (n_0_1_644), .A1 (n_0_1_648), .A2 (opt_ipo_n5152));
NAND2_X4 i_0_1_1343 (.ZN (n_0_1_926), .A1 (n_0_1_646), .A2 (opt_ipo_n5152));
INV_X8 i_0_1_1342 (.ZN (n_0_1_645), .A (n_0_1_926));
AOI22_X1 i_0_1_1333 (.ZN (n_0_1_925), .A1 (\A_imm_2s_complement[30] ), .A2 (CLOCK_spw__n7344)
    , .B1 (\A_imm[29] ), .B2 (opt_ipo_n5395));
NAND2_X4 i_0_1_1332 (.ZN (n_0_1_643), .A1 (n_0_1_646), .A2 (n_0_1_651));
NOR3_X4 i_0_1_1325 (.ZN (n_0_1_642), .A1 (opt_ipo_n5682), .A2 (opt_ipo_n5398), .A3 (n_0_1_651));
NAND2_X1 i_0_1_1324 (.ZN (n_0_1_924), .A1 (\A_imm_2s_complement[29] ), .A2 (opt_ipo_n5393));
OAI211_X1 i_0_1_1301 (.ZN (n_0_743), .A (n_0_1_925), .B (n_0_1_924), .C1 (sgo__n734), .C2 (n_0_1_643));
NAND2_X1 i_0_1_1300 (.ZN (n_0_1_923), .A1 (\A_imm_2s_complement[25] ), .A2 (opt_ipo_n5393));
AOI22_X1 i_0_1_1279 (.ZN (n_0_1_922), .A1 (\A_imm_2s_complement[26] ), .A2 (CLOCK_spw__n7344)
    , .B1 (opt_ipo_n5362), .B2 (opt_ipo_n5395));
OAI211_X1 i_0_1_1278 (.ZN (n_0_739), .A (n_0_1_922), .B (n_0_1_923), .C1 (slo__xsl_n1889), .C2 (n_0_1_643));
INV_X4 opt_ipo_c5730 (.ZN (opt_ipo_n5146), .A (sgo__n847));
INV_X4 i_0_1_1276 (.ZN (n_0_1_599), .A (slo__sro_n1458));
AOI222_X1 slo__sro_c4279 (.ZN (n_0_1_401), .A1 (n_0_1_430), .A2 (opt_ipo_n5205), .B1 (opt_ipo_n5419)
    , .B2 (\A_imm_2s_complement[5] ), .C1 (opt_ipo_n5686), .C2 (slo__n3378));
INV_X1 slo__sro_c4554 (.ZN (slo__sro_n4176), .A (drc_ipo_n58));
AOI22_X1 i_0_1_1203 (.ZN (n_0_1_919), .A1 (\A_imm_2s_complement[30] ), .A2 (slo__n4931)
    , .B1 (\A_imm_2s_complement[29] ), .B2 (spw__n7778));
NAND2_X1 i_0_1_1202 (.ZN (slo__n1580), .A1 (opt_ipo_n5315), .A2 (n_0_1_603));
CLKBUF_X1 slo__c3664 (.Z (slo__n3345), .A (CLOCK_spw__n7299));
NAND2_X1 i_0_1_1200 (.ZN (n_0_1_918), .A1 (\A_imm[29] ), .A2 (opt_ipo_n5311));
OAI211_X1 i_0_1_1197 (.ZN (n_0_710), .A (n_0_1_919), .B (n_0_1_918), .C1 (sgo__n734), .C2 (n_0_1_600));
NAND2_X1 i_0_1_1196 (.ZN (n_0_1_917), .A1 (\A_imm_2s_complement[21] ), .A2 (spw__n7777));
AOI22_X1 i_0_1_1189 (.ZN (n_0_1_916), .A1 (\A_imm_2s_complement[22] ), .A2 (slo__n4931)
    , .B1 (opt_ipo_n5135), .B2 (opt_ipo_n5312));
OAI211_X1 i_0_1_1188 (.ZN (n_0_702), .A (n_0_1_916), .B (n_0_1_917), .C1 (slo__xsl_n1641), .C2 (n_0_1_600));
OAI21_X1 slo__sro_c4012 (.ZN (slo__sro_n3675), .A (sgo__n759), .B1 (drc_ipo_n48), .B2 (opt_ipo_n5224));
NAND2_X1 i_0_1_1126 (.ZN (n_0_1_915), .A1 (\A_imm_2s_complement[30] ), .A2 (opt_ipo_n5258));
NAND2_X4 i_0_1_1125 (.ZN (n_0_1_557), .A1 (n_0_1_560), .A2 (n_0_1_565));
NOR2_X4 i_0_1_1124 (.ZN (n_0_1_558), .A1 (n_0_1_562), .A2 (slo___n3489));
NAND2_X4 i_0_1_1121 (.ZN (n_0_1_914), .A1 (slo__n3691), .A2 (slo___n3496));
INV_X4 i_0_1_1120 (.ZN (n_0_1_559), .A (n_0_1_914));
AOI22_X1 i_0_1_1105 (.ZN (n_0_1_913), .A1 (\A_imm_2s_complement[31] ), .A2 (slo___n2464)
    , .B1 (\A_imm[30] ), .B2 (opt_ipo_n5774));
OAI211_X1 i_0_1_1104 (.ZN (n_0_678), .A (n_0_1_913), .B (n_0_1_915), .C1 (n_0_1_836), .C2 (n_0_1_557));
AOI22_X1 i_0_1_1051 (.ZN (n_0_1_912), .A1 (opt_ipo_n5358), .A2 (slo___n2464), .B1 (sgo__n1241), .B2 (opt_ipo_n5258));
NAND2_X1 i_0_1_1050 (.ZN (n_0_1_911), .A1 (\A_imm[29] ), .A2 (opt_ipo_n5774));
OAI211_X1 i_0_1_1049 (.ZN (n_0_677), .A (n_0_1_912), .B (n_0_1_911), .C1 (sgo__n734), .C2 (n_0_1_557));
NAND2_X1 i_0_1_1048 (.ZN (n_0_1_910), .A1 (CLOCK_slh_n7157), .A2 (clk));
NAND2_X4 i_0_1_1047 (.ZN (n_0_283), .A1 (n_0_1_910), .A2 (hfn_ipo_n46));
INV_X1 i_0_1_1046 (.ZN (n_0_1_909), .A (n_0_124));
XNOR2_X2 i_0_1_1045 (.ZN (n_0_1_908), .A (A_in), .B (drc_ipo_n58));
INV_X1 i_0_1_1044 (.ZN (n_0_1_907), .A (n_0_813));
INV_X1 i_0_1_219 (.ZN (n_0_1_906), .A (\aggregated_res[14][5] ));
INV_X1 i_0_1_218 (.ZN (n_0_1_905), .A (\aggregated_res[14][4] ));
INV_X1 i_0_1_217 (.ZN (n_0_1_904), .A (\aggregated_res[14][3] ));
INV_X1 i_0_1_216 (.ZN (n_0_1_903), .A (\aggregated_res[14][2] ));
NAND4_X1 i_0_1_215 (.ZN (n_0_1_902), .A1 (n_0_1_906), .A2 (n_0_1_905), .A3 (n_0_1_904), .A4 (n_0_1_903));
INV_X1 i_0_1_214 (.ZN (n_0_1_901), .A (\aggregated_res[14][9] ));
INV_X1 i_0_1_213 (.ZN (n_0_1_900), .A (\aggregated_res[14][8] ));
INV_X1 i_0_1_212 (.ZN (n_0_1_899), .A (\aggregated_res[14][7] ));
INV_X1 i_0_1_211 (.ZN (n_0_1_898), .A (\aggregated_res[14][6] ));
NAND4_X1 i_0_1_210 (.ZN (n_0_1_897), .A1 (n_0_1_901), .A2 (n_0_1_900), .A3 (n_0_1_899), .A4 (n_0_1_898));
BUF_X4 sgo__c817 (.Z (sgo__n839), .A (\A_imm_2s_complement[23] ));
BUF_X8 sgo__c710 (.Z (sgo__n759), .A (drc_ipo_n59));
BUF_X4 sgo__c875 (.Z (sgo__n877), .A (\A_imm_2s_complement[27] ));
INV_X1 i_0_1_205 (.ZN (n_0_1_892), .A (\aggregated_res[14][50] ));
INV_X4 i_0_1_204 (.ZN (n_0_1_891), .A (\aggregated_res[14][49] ));
INV_X4 i_0_1_203 (.ZN (n_0_1_890), .A (\aggregated_res[14][48] ));
INV_X4 i_0_1_202 (.ZN (n_0_1_889), .A (\aggregated_res[14][47] ));
INV_X1 i_0_1_200 (.ZN (n_0_1_887), .A (\aggregated_res[14][32] ));
INV_X1 i_0_1_199 (.ZN (n_0_1_886), .A (\aggregated_res[14][31] ));
INV_X1 i_0_1_198 (.ZN (n_0_1_885), .A (\aggregated_res[14][15] ));
INV_X1 i_0_1_197 (.ZN (n_0_1_884), .A (\aggregated_res[14][14] ));
NAND4_X1 i_0_1_196 (.ZN (n_0_1_883), .A1 (n_0_1_887), .A2 (n_0_1_886), .A3 (n_0_1_885), .A4 (n_0_1_884));
NOR3_X4 i_0_1_195 (.ZN (n_0_1_882), .A1 (n_0_1_888), .A2 (\aggregated_res[14][59] ), .A3 (n_0_1_883));
INV_X2 i_0_1_194 (.ZN (n_0_1_881), .A (\aggregated_res[14][58] ));
INV_X2 i_0_1_193 (.ZN (n_0_1_880), .A (\aggregated_res[14][57] ));
INV_X1 i_0_1_192 (.ZN (n_0_1_879), .A (\aggregated_res[14][56] ));
INV_X2 i_0_1_191 (.ZN (n_0_1_878), .A (\aggregated_res[14][55] ));
NAND4_X4 i_0_1_190 (.ZN (n_0_1_877), .A1 (n_0_1_880), .A2 (n_0_1_881), .A3 (slo__n2528), .A4 (n_0_1_878));
INV_X1 i_0_1_188 (.ZN (n_0_1_875), .A (\aggregated_res[14][13] ));
INV_X1 i_0_1_187 (.ZN (n_0_1_874), .A (\aggregated_res[14][12] ));
INV_X1 i_0_1_186 (.ZN (n_0_1_873), .A (\aggregated_res[14][11] ));
INV_X1 i_0_1_185 (.ZN (n_0_1_872), .A (\aggregated_res[14][10] ));
NAND4_X1 i_0_1_184 (.ZN (n_0_1_871), .A1 (n_0_1_875), .A2 (n_0_1_874), .A3 (n_0_1_873), .A4 (n_0_1_872));
INV_X1 i_0_1_183 (.ZN (n_0_1_870), .A (\aggregated_res[14][62] ));
INV_X2 i_0_1_182 (.ZN (n_0_1_869), .A (\aggregated_res[14][61] ));
INV_X1 i_0_1_181 (.ZN (n_0_1_838), .A (\aggregated_res[14][60] ));
CLKBUF_X2 slo__c3544 (.Z (slo__n3230), .A (\A_imm[12] ));
NAND2_X4 sgo__sro_c726 (.ZN (sgo__sro_n770), .A1 (sgo__sro_n771), .A2 (sgo__sro_n772));
NOR2_X2 CLOCK_slo__mro_c7543 (.ZN (CLOCK_slo__mro_n6799), .A1 (\aggregated_res[14][44] ), .A2 (\aggregated_res[14][43] ));
NOR2_X2 sgo__c862 (.ZN (opt_ipo_n5506), .A1 (opt_ipo_n5239), .A2 (A_in));
NOR2_X2 i_0_1_176 (.ZN (n_0_1_769), .A1 (sgo__sro_n1272), .A2 (n_0_1_908));
NAND2_X2 i_0_1_175 (.ZN (n_0_1_767), .A1 (slo__n2232), .A2 (hfn_ipo_n46));
NOR2_X4 i_0_1_174 (.ZN (n_0_1_755), .A1 (n_0_1_769), .A2 (reset));
NAND2_X1 i_0_1_173 (.ZN (n_0_1_754), .A1 (n_0_1_755), .A2 (\aggregated_res[14][63] ));
OAI21_X1 i_0_1_172 (.ZN (n_0_250), .A (n_0_1_754), .B1 (sgo__n1223), .B2 (n_0_1_909));
INV_X1 i_0_1_171 (.ZN (n_0_1_753), .A (n_0_123));
INV_X8 i_0_1_170 (.ZN (n_0_1_752), .A (n_0_1_755));
OAI22_X1 i_0_1_169 (.ZN (n_0_249), .A1 (n_0_1_753), .A2 (sgo__n1223), .B1 (hfn_ipo_n43), .B2 (n_0_1_870));
INV_X1 i_0_1_168 (.ZN (n_0_1_749), .A (n_0_122));
OAI22_X1 i_0_1_167 (.ZN (n_0_248), .A1 (n_0_1_749), .A2 (sgo__n1223), .B1 (hfn_ipo_n43), .B2 (n_0_1_869));
INV_X1 i_0_1_166 (.ZN (n_0_1_727), .A (n_0_121));
OAI22_X1 i_0_1_165 (.ZN (n_0_247), .A1 (n_0_1_727), .A2 (sgo__n1223), .B1 (hfn_ipo_n43), .B2 (n_0_1_838));
INV_X1 sgo__sro_c1281 (.ZN (sgo__sro_n1197), .A (opt_ipo_n5258));
NAND2_X1 i_0_1_163 (.ZN (n_0_1_724), .A1 (n_0_1_755), .A2 (\aggregated_res[14][59] ));
OAI21_X1 i_0_1_162 (.ZN (n_0_246), .A (n_0_1_724), .B1 (sgo__n1223), .B2 (n_0_120));
INV_X1 i_0_1_161 (.ZN (n_0_1_723), .A (n_0_119));
OAI22_X1 i_0_1_160 (.ZN (n_0_245), .A1 (n_0_1_723), .A2 (sgo__n1223), .B1 (hfn_ipo_n43), .B2 (n_0_1_881));
INV_X1 CLOCK_slo__sro_c7469 (.ZN (CLOCK_slo__sro_n6742), .A (slo__xsl_n1425));
OAI22_X1 i_0_1_158 (.ZN (n_0_244), .A1 (n_0_118), .A2 (sgo__n1223), .B1 (hfn_ipo_n43), .B2 (n_0_1_880));
INV_X1 i_0_1_157 (.ZN (n_0_1_714), .A (n_0_117));
OAI22_X1 i_0_1_156 (.ZN (n_0_243), .A1 (n_0_1_714), .A2 (sgo__n1223), .B1 (hfn_ipo_n43), .B2 (n_0_1_879));
INV_X16 i_0_1_155 (.ZN (n_0_1_702), .A (slo__n2400));
NAND2_X4 i_0_1_154 (.ZN (n_0_1_679), .A1 (n_0_1_702), .A2 (n_0_116));
OAI21_X2 i_0_1_153 (.ZN (n_0_242), .A (n_0_1_679), .B1 (hfn_ipo_n43), .B2 (n_0_1_878));
INV_X1 i_0_1_152 (.ZN (n_0_1_640), .A (n_0_115));
NAND2_X1 i_0_1_151 (.ZN (n_0_1_636), .A1 (n_0_1_755), .A2 (\aggregated_res[14][54] ));
OAI21_X1 i_0_1_150 (.ZN (n_0_241), .A (n_0_1_636), .B1 (sgo__n1223), .B2 (n_0_1_640));
INV_X1 i_0_1_149 (.ZN (n_0_1_597), .A (n_0_114));
NAND2_X1 i_0_1_148 (.ZN (n_0_1_589), .A1 (n_0_1_755), .A2 (\aggregated_res[14][53] ));
OAI21_X1 i_0_1_147 (.ZN (n_0_240), .A (n_0_1_589), .B1 (sgo__n1223), .B2 (n_0_1_597));
INV_X1 i_0_1_142 (.ZN (n_0_1_555), .A (n_0_113));
NAND2_X1 i_0_1_137 (.ZN (n_0_1_554), .A1 (n_0_1_755), .A2 (\aggregated_res[14][52] ));
OAI21_X1 i_0_1_136 (.ZN (n_0_239), .A (n_0_1_554), .B1 (sgo__n1223), .B2 (n_0_1_555));
NAND2_X1 i_0_1_135 (.ZN (n_0_1_89), .A1 (n_0_1_702), .A2 (n_0_112));
NAND2_X1 i_0_1_134 (.ZN (n_0_1_88), .A1 (n_0_1_755), .A2 (\aggregated_res[14][51] ));
NAND2_X1 i_0_1_133 (.ZN (n_0_238), .A1 (n_0_1_89), .A2 (n_0_1_88));
INV_X2 i_0_1_132 (.ZN (n_0_1_87), .A (n_0_111));
OAI22_X1 i_0_1_131 (.ZN (n_0_237), .A1 (n_0_1_87), .A2 (sgo__n1223), .B1 (hfn_ipo_n43), .B2 (n_0_1_892));
INV_X1 i_0_1_130 (.ZN (n_0_1_86), .A (n_0_110));
OAI22_X2 i_0_1_129 (.ZN (n_0_236), .A1 (n_0_1_86), .A2 (sgo__n1223), .B1 (hfn_ipo_n43), .B2 (n_0_1_891));
NAND2_X1 i_0_1_128 (.ZN (n_0_1_85), .A1 (n_0_1_702), .A2 (n_0_109));
OAI21_X1 i_0_1_127 (.ZN (n_0_235), .A (n_0_1_85), .B1 (hfn_ipo_n43), .B2 (n_0_1_890));
NAND2_X1 i_0_1_126 (.ZN (n_0_1_84), .A1 (slo__n2517), .A2 (n_0_108));
OAI21_X2 i_0_1_125 (.ZN (n_0_234), .A (n_0_1_84), .B1 (hfn_ipo_n43), .B2 (n_0_1_889));
INV_X1 i_0_1_124 (.ZN (n_0_1_83), .A (\aggregated_res[14][46] ));
NAND2_X1 i_0_1_123 (.ZN (n_0_1_78), .A1 (n_0_1_702), .A2 (n_0_107));
OAI21_X1 i_0_1_122 (.ZN (n_0_233), .A (n_0_1_78), .B1 (hfn_ipo_n43), .B2 (n_0_1_83));
INV_X1 i_0_1_121 (.ZN (n_0_1_73), .A (\aggregated_res[14][45] ));
NAND2_X1 i_0_1_120 (.ZN (n_0_1_72), .A1 (n_0_1_702), .A2 (n_0_106));
OAI21_X1 i_0_1_119 (.ZN (n_0_232), .A (n_0_1_72), .B1 (hfn_ipo_n43), .B2 (n_0_1_73));
INV_X1 i_0_1_118 (.ZN (n_0_1_71), .A (\aggregated_res[14][44] ));
NAND2_X1 i_0_1_117 (.ZN (n_0_1_70), .A1 (slo__n1376), .A2 (n_0_105));
OAI21_X1 i_0_1_116 (.ZN (n_0_231), .A (n_0_1_70), .B1 (hfn_ipo_n43), .B2 (n_0_1_71));
INV_X1 i_0_1_115 (.ZN (n_0_1_69), .A (\aggregated_res[14][43] ));
NAND2_X1 i_0_1_114 (.ZN (n_0_1_68), .A1 (n_0_1_702), .A2 (n_0_104));
OAI21_X1 i_0_1_113 (.ZN (n_0_230), .A (n_0_1_68), .B1 (hfn_ipo_n43), .B2 (n_0_1_69));
INV_X1 i_0_1_112 (.ZN (n_0_1_67), .A (\aggregated_res[14][42] ));
NAND2_X1 i_0_1_111 (.ZN (n_0_1_66), .A1 (slo__n2517), .A2 (n_0_103));
OAI21_X2 i_0_1_110 (.ZN (n_0_229), .A (n_0_1_66), .B1 (hfn_ipo_n43), .B2 (n_0_1_67));
INV_X1 i_0_1_109 (.ZN (n_0_1_65), .A (\aggregated_res[14][41] ));
NAND2_X4 i_0_1_108 (.ZN (n_0_1_64), .A1 (n_0_1_702), .A2 (n_0_102));
OAI21_X1 i_0_1_107 (.ZN (n_0_228), .A (n_0_1_64), .B1 (hfn_ipo_n43), .B2 (n_0_1_65));
INV_X1 i_0_1_106 (.ZN (n_0_1_63), .A (\aggregated_res[14][40] ));
NAND2_X1 i_0_1_105 (.ZN (n_0_1_62), .A1 (n_0_1_702), .A2 (n_0_101));
OAI21_X1 i_0_1_104 (.ZN (n_0_227), .A (n_0_1_62), .B1 (hfn_ipo_n43), .B2 (n_0_1_63));
INV_X1 i_0_1_103 (.ZN (n_0_1_61), .A (\aggregated_res[14][39] ));
NAND2_X1 i_0_1_102 (.ZN (n_0_1_60), .A1 (n_0_1_702), .A2 (n_0_100));
OAI21_X1 i_0_1_101 (.ZN (n_0_226), .A (n_0_1_60), .B1 (hfn_ipo_n43), .B2 (n_0_1_61));
INV_X1 i_0_1_100 (.ZN (n_0_1_59), .A (\aggregated_res[14][38] ));
NAND2_X1 i_0_1_99 (.ZN (n_0_1_58), .A1 (n_0_1_702), .A2 (n_0_99));
OAI21_X1 i_0_1_98 (.ZN (n_0_225), .A (n_0_1_58), .B1 (hfn_ipo_n43), .B2 (n_0_1_59));
INV_X1 i_0_1_97 (.ZN (n_0_1_57), .A (\aggregated_res[14][37] ));
NAND2_X1 i_0_1_96 (.ZN (n_0_1_56), .A1 (n_0_1_702), .A2 (n_0_98));
OAI21_X1 i_0_1_95 (.ZN (n_0_224), .A (n_0_1_56), .B1 (hfn_ipo_n43), .B2 (n_0_1_57));
INV_X1 i_0_1_94 (.ZN (n_0_1_55), .A (\aggregated_res[14][36] ));
NAND2_X1 i_0_1_93 (.ZN (n_0_1_54), .A1 (n_0_1_702), .A2 (n_0_97));
OAI21_X1 i_0_1_92 (.ZN (n_0_223), .A (n_0_1_54), .B1 (hfn_ipo_n43), .B2 (n_0_1_55));
INV_X1 i_0_1_91 (.ZN (n_0_1_53), .A (\aggregated_res[14][35] ));
NAND2_X1 i_0_1_90 (.ZN (n_0_1_52), .A1 (n_0_1_702), .A2 (n_0_96));
OAI21_X1 i_0_1_89 (.ZN (n_0_222), .A (n_0_1_52), .B1 (hfn_ipo_n44), .B2 (n_0_1_53));
INV_X1 i_0_1_88 (.ZN (n_0_1_51), .A (\aggregated_res[14][34] ));
NAND2_X2 i_0_1_87 (.ZN (n_0_1_50), .A1 (n_0_1_702), .A2 (n_0_95));
OAI21_X1 i_0_1_86 (.ZN (n_0_221), .A (n_0_1_50), .B1 (hfn_ipo_n44), .B2 (n_0_1_51));
INV_X1 i_0_1_85 (.ZN (n_0_1_49), .A (\aggregated_res[14][33] ));
NAND2_X1 i_0_1_84 (.ZN (n_0_1_48), .A1 (n_0_1_702), .A2 (n_0_94));
OAI21_X1 i_0_1_83 (.ZN (n_0_220), .A (n_0_1_48), .B1 (hfn_ipo_n44), .B2 (n_0_1_49));
NAND2_X2 i_0_1_82 (.ZN (n_0_1_47), .A1 (n_0_1_702), .A2 (n_0_93));
OAI21_X1 i_0_1_81 (.ZN (n_0_219), .A (n_0_1_47), .B1 (hfn_ipo_n44), .B2 (n_0_1_887));
NAND2_X4 i_0_1_80 (.ZN (n_0_1_46), .A1 (n_0_1_702), .A2 (n_0_92));
OAI21_X1 i_0_1_79 (.ZN (n_0_218), .A (n_0_1_46), .B1 (hfn_ipo_n44), .B2 (n_0_1_886));
INV_X1 i_0_1_78 (.ZN (n_0_1_45), .A (\aggregated_res[14][30] ));
NAND2_X4 i_0_1_77 (.ZN (n_0_1_44), .A1 (n_0_1_702), .A2 (n_0_91));
OAI21_X1 i_0_1_76 (.ZN (n_0_217), .A (n_0_1_44), .B1 (hfn_ipo_n44), .B2 (n_0_1_45));
INV_X1 i_0_1_75 (.ZN (n_0_1_43), .A (\aggregated_res[14][29] ));
NAND2_X4 i_0_1_74 (.ZN (n_0_1_42), .A1 (n_0_1_702), .A2 (n_0_90));
OAI21_X2 i_0_1_73 (.ZN (n_0_216), .A (n_0_1_42), .B1 (hfn_ipo_n44), .B2 (n_0_1_43));
INV_X1 i_0_1_72 (.ZN (n_0_1_41), .A (\aggregated_res[14][28] ));
NAND2_X2 i_0_1_71 (.ZN (n_0_1_40), .A1 (slo__n2235), .A2 (n_0_89));
OAI21_X2 i_0_1_70 (.ZN (n_0_215), .A (n_0_1_40), .B1 (hfn_ipo_n44), .B2 (n_0_1_41));
INV_X1 i_0_1_69 (.ZN (n_0_1_39), .A (\aggregated_res[14][27] ));
NAND2_X1 i_0_1_68 (.ZN (n_0_1_38), .A1 (slo__n2235), .A2 (n_0_88));
OAI21_X1 i_0_1_67 (.ZN (n_0_214), .A (n_0_1_38), .B1 (hfn_ipo_n44), .B2 (n_0_1_39));
INV_X1 i_0_1_66 (.ZN (n_0_1_37), .A (\aggregated_res[14][26] ));
NAND2_X1 i_0_1_65 (.ZN (n_0_1_36), .A1 (slo__n2235), .A2 (n_0_87));
OAI21_X1 i_0_1_64 (.ZN (n_0_213), .A (n_0_1_36), .B1 (hfn_ipo_n44), .B2 (n_0_1_37));
INV_X1 i_0_1_63 (.ZN (n_0_1_35), .A (\aggregated_res[14][25] ));
NAND2_X1 i_0_1_62 (.ZN (n_0_1_34), .A1 (slo__n2235), .A2 (n_0_86));
OAI21_X1 i_0_1_61 (.ZN (n_0_212), .A (n_0_1_34), .B1 (hfn_ipo_n44), .B2 (n_0_1_35));
INV_X1 i_0_1_60 (.ZN (n_0_1_33), .A (\aggregated_res[14][24] ));
NAND2_X1 i_0_1_59 (.ZN (n_0_1_32), .A1 (slo__n2235), .A2 (n_0_85));
OAI21_X1 i_0_1_58 (.ZN (n_0_211), .A (n_0_1_32), .B1 (hfn_ipo_n44), .B2 (n_0_1_33));
INV_X1 i_0_1_57 (.ZN (n_0_1_31), .A (\aggregated_res[14][23] ));
NAND2_X2 i_0_1_56 (.ZN (n_0_1_30), .A1 (slo__n1376), .A2 (n_0_84));
OAI21_X2 i_0_1_55 (.ZN (n_0_210), .A (n_0_1_30), .B1 (hfn_ipo_n44), .B2 (n_0_1_31));
INV_X1 i_0_1_54 (.ZN (n_0_1_29), .A (\aggregated_res[14][22] ));
NAND2_X2 i_0_1_53 (.ZN (n_0_1_28), .A1 (slo__n1376), .A2 (n_0_83));
OAI21_X1 i_0_1_52 (.ZN (n_0_209), .A (n_0_1_28), .B1 (hfn_ipo_n44), .B2 (n_0_1_29));
INV_X1 i_0_1_51 (.ZN (n_0_1_27), .A (\aggregated_res[14][21] ));
NAND2_X1 i_0_1_50 (.ZN (n_0_1_26), .A1 (slo__n1376), .A2 (n_0_82));
OAI21_X1 i_0_1_49 (.ZN (n_0_208), .A (n_0_1_26), .B1 (hfn_ipo_n44), .B2 (n_0_1_27));
INV_X1 i_0_1_48 (.ZN (n_0_1_25), .A (\aggregated_res[14][20] ));
NAND2_X1 i_0_1_47 (.ZN (n_0_1_24), .A1 (slo__n1376), .A2 (n_0_81));
OAI21_X1 i_0_1_46 (.ZN (n_0_207), .A (n_0_1_24), .B1 (hfn_ipo_n44), .B2 (n_0_1_25));
INV_X1 i_0_1_45 (.ZN (n_0_1_23), .A (\aggregated_res[14][19] ));
NAND2_X1 i_0_1_44 (.ZN (n_0_1_22), .A1 (slo__n1376), .A2 (n_0_80));
OAI21_X1 i_0_1_43 (.ZN (n_0_206), .A (n_0_1_22), .B1 (hfn_ipo_n44), .B2 (n_0_1_23));
INV_X1 i_0_1_42 (.ZN (n_0_1_21), .A (\aggregated_res[14][18] ));
NAND2_X1 i_0_1_41 (.ZN (n_0_1_20), .A1 (slo__n1376), .A2 (n_0_79));
OAI21_X1 i_0_1_40 (.ZN (n_0_205), .A (n_0_1_20), .B1 (hfn_ipo_n44), .B2 (n_0_1_21));
INV_X1 i_0_1_39 (.ZN (n_0_1_19), .A (\aggregated_res[14][17] ));
NAND2_X1 i_0_1_38 (.ZN (n_0_1_18), .A1 (slo__n1376), .A2 (n_0_78));
OAI21_X1 i_0_1_37 (.ZN (n_0_204), .A (n_0_1_18), .B1 (hfn_ipo_n44), .B2 (n_0_1_19));
INV_X1 i_0_1_36 (.ZN (n_0_1_17), .A (\aggregated_res[14][16] ));
NAND2_X1 i_0_1_35 (.ZN (n_0_1_16), .A1 (slo__n2235), .A2 (n_0_77));
OAI21_X1 i_0_1_34 (.ZN (n_0_203), .A (n_0_1_16), .B1 (hfn_ipo_n44), .B2 (n_0_1_17));
NAND2_X4 i_0_1_33 (.ZN (n_0_1_15), .A1 (n_0_1_702), .A2 (n_0_76));
OAI21_X2 i_0_1_32 (.ZN (n_0_202), .A (n_0_1_15), .B1 (hfn_ipo_n44), .B2 (n_0_1_885));
NAND2_X4 i_0_1_31 (.ZN (n_0_1_14), .A1 (n_0_1_702), .A2 (n_0_75));
OAI21_X2 i_0_1_30 (.ZN (n_0_201), .A (n_0_1_14), .B1 (hfn_ipo_n44), .B2 (n_0_1_884));
NAND2_X4 i_0_1_29 (.ZN (n_0_1_13), .A1 (n_0_1_702), .A2 (n_0_74));
OAI21_X1 i_0_1_28 (.ZN (n_0_200), .A (n_0_1_13), .B1 (hfn_ipo_n44), .B2 (n_0_1_875));
NAND2_X4 i_0_1_27 (.ZN (n_0_1_12), .A1 (n_0_1_702), .A2 (n_0_73));
OAI21_X1 i_0_1_26 (.ZN (n_0_199), .A (n_0_1_12), .B1 (hfn_ipo_n44), .B2 (n_0_1_874));
NAND2_X4 i_0_1_25 (.ZN (n_0_1_11), .A1 (n_0_1_702), .A2 (n_0_72));
OAI21_X1 i_0_1_24 (.ZN (n_0_198), .A (n_0_1_11), .B1 (hfn_ipo_n44), .B2 (n_0_1_873));
NAND2_X4 i_0_1_23 (.ZN (n_0_1_10), .A1 (n_0_1_702), .A2 (n_0_71));
OAI21_X1 i_0_1_22 (.ZN (n_0_197), .A (n_0_1_10), .B1 (hfn_ipo_n44), .B2 (n_0_1_872));
NAND2_X4 i_0_1_21 (.ZN (n_0_1_9), .A1 (n_0_1_702), .A2 (n_0_70));
OAI21_X1 i_0_1_20 (.ZN (n_0_196), .A (n_0_1_9), .B1 (hfn_ipo_n44), .B2 (n_0_1_901));
NAND2_X4 i_0_1_19 (.ZN (n_0_1_8), .A1 (n_0_1_702), .A2 (n_0_69));
OAI21_X1 i_0_1_18 (.ZN (n_0_195), .A (n_0_1_8), .B1 (hfn_ipo_n44), .B2 (n_0_1_900));
NAND2_X4 i_0_1_17 (.ZN (n_0_1_7), .A1 (n_0_1_702), .A2 (n_0_68));
OAI21_X1 i_0_1_16 (.ZN (n_0_194), .A (n_0_1_7), .B1 (hfn_ipo_n44), .B2 (n_0_1_899));
NAND2_X4 i_0_1_15 (.ZN (n_0_1_6), .A1 (n_0_1_702), .A2 (n_0_67));
OAI21_X1 i_0_1_14 (.ZN (n_0_193), .A (n_0_1_6), .B1 (hfn_ipo_n44), .B2 (n_0_1_898));
NAND2_X4 i_0_1_13 (.ZN (n_0_1_5), .A1 (n_0_1_702), .A2 (n_0_66));
OAI21_X1 i_0_1_12 (.ZN (n_0_192), .A (n_0_1_5), .B1 (hfn_ipo_n44), .B2 (n_0_1_906));
NAND2_X4 i_0_1_11 (.ZN (n_0_1_4), .A1 (n_0_1_702), .A2 (n_0_65));
OAI21_X1 i_0_1_10 (.ZN (n_0_191), .A (n_0_1_4), .B1 (hfn_ipo_n44), .B2 (n_0_1_905));
NAND2_X4 i_0_1_9 (.ZN (n_0_1_3), .A1 (n_0_1_702), .A2 (n_0_64));
OAI21_X1 i_0_1_8 (.ZN (n_0_190), .A (n_0_1_3), .B1 (hfn_ipo_n44), .B2 (n_0_1_904));
INV_X1 i_0_1_7 (.ZN (n_0_1_2), .A (n_0_63));
NAND2_X1 i_0_1_6 (.ZN (n_0_1_1), .A1 (n_0_1_908), .A2 (hfn_ipo_n46));
OAI22_X1 i_0_1_5 (.ZN (n_0_189), .A1 (sgo__n1223), .A2 (n_0_1_2), .B1 (n_0_1_903), .B2 (n_0_1_1));
INV_X1 i_0_1_4 (.ZN (n_0_1_0), .A (n_0_62));
OAI22_X1 i_0_1_3 (.ZN (n_0_188), .A1 (sgo__n1223), .A2 (n_0_1_0), .B1 (n_0_1_907), .B2 (n_0_1_1));
INV_X2 i_0_1_2 (.ZN (n_0_1_776), .A (opt_ipo_n5459));
INV_X2 i_0_1_1 (.ZN (n_0_1_784), .A (slo__n3378));
INV_X1 i_0_1_1558 (.ZN (n_0_1_868), .A (n_0_157));
INV_X1 i_0_1_1557 (.ZN (n_0_1_867), .A (n_0_125));
INV_X1 i_0_1_1556 (.ZN (n_0_1_866), .A (n_0_126));
INV_X1 i_0_1_1555 (.ZN (n_0_1_865), .A (n_0_127));
INV_X1 i_0_1_1554 (.ZN (n_0_1_864), .A (n_0_128));
INV_X1 i_0_1_1553 (.ZN (n_0_1_863), .A (n_0_129));
INV_X1 i_0_1_1552 (.ZN (n_0_1_862), .A (n_0_130));
INV_X1 i_0_1_1551 (.ZN (n_0_1_861), .A (n_0_131));
INV_X1 i_0_1_1550 (.ZN (n_0_1_860), .A (n_0_132));
INV_X1 i_0_1_1549 (.ZN (n_0_1_859), .A (n_0_133));
INV_X1 i_0_1_1548 (.ZN (n_0_1_858), .A (n_0_134));
INV_X1 i_0_1_1547 (.ZN (n_0_1_857), .A (n_0_135));
INV_X1 i_0_1_1546 (.ZN (n_0_1_856), .A (n_0_136));
INV_X1 i_0_1_1545 (.ZN (n_0_1_855), .A (n_0_137));
INV_X1 i_0_1_1544 (.ZN (n_0_1_854), .A (n_0_138));
INV_X1 i_0_1_1543 (.ZN (n_0_1_853), .A (n_0_139));
INV_X1 i_0_1_1542 (.ZN (n_0_1_852), .A (n_0_140));
INV_X1 i_0_1_1541 (.ZN (n_0_1_851), .A (opt_ipo_n5711));
INV_X1 i_0_1_1540 (.ZN (n_0_1_850), .A (n_0_142));
INV_X1 i_0_1_1539 (.ZN (n_0_1_849), .A (n_0_143));
INV_X1 i_0_1_1538 (.ZN (n_0_1_848), .A (n_0_144));
INV_X1 i_0_1_1537 (.ZN (n_0_1_847), .A (n_0_145));
INV_X1 i_0_1_1536 (.ZN (n_0_1_846), .A (n_0_146));
INV_X1 i_0_1_1535 (.ZN (n_0_1_845), .A (n_0_147));
INV_X1 i_0_1_1534 (.ZN (n_0_1_844), .A (n_0_148));
INV_X1 i_0_1_1533 (.ZN (n_0_1_843), .A (opt_ipo_n5702));
INV_X1 i_0_1_1532 (.ZN (n_0_1_842), .A (n_0_150));
INV_X1 i_0_1_1531 (.ZN (n_0_1_841), .A (n_0_151));
INV_X1 i_0_1_1530 (.ZN (n_0_1_840), .A (n_0_152));
INV_X1 i_0_1_1529 (.ZN (n_0_1_839), .A (n_0_153));
INV_X4 i_0_1_1525 (.ZN (\A_imm[31] ), .A (n_0_1_836));
NOR2_X1 i_0_1_1524 (.ZN (n_0_1_835), .A1 (n_0_1_867), .A2 (A_in));
NOR2_X1 i_0_1_1521 (.ZN (n_0_1_833), .A1 (n_0_1_866), .A2 (A_in));
NOR2_X1 i_0_1_1518 (.ZN (n_0_1_831), .A1 (n_0_1_865), .A2 (A_in));
INV_X8 i_0_1_1516 (.ZN (\A_imm[28] ), .A (n_0_1_830));
NOR2_X1 i_0_1_1515 (.ZN (n_0_1_829), .A1 (n_0_1_864), .A2 (hfn_ipo_n41));
NOR2_X1 i_0_1_1512 (.ZN (n_0_1_827), .A1 (n_0_1_863), .A2 (hfn_ipo_n41));
NOR2_X1 i_0_1_1509 (.ZN (n_0_1_825), .A1 (n_0_1_862), .A2 (hfn_ipo_n41));
AOI21_X4 i_0_1_1508 (.ZN (sgo__n880), .A (n_0_1_825), .B1 (n_0_24), .B2 (hfn_ipo_n41));
NOR2_X1 i_0_1_1506 (.ZN (n_0_1_823), .A1 (n_0_1_861), .A2 (hfn_ipo_n41));
AOI21_X4 i_0_1_1505 (.ZN (n_0_1_822), .A (n_0_1_823), .B1 (n_0_23), .B2 (hfn_ipo_n41));
INV_X4 i_0_1_1504 (.ZN (\A_imm[24] ), .A (n_0_1_822));
NOR2_X1 i_0_1_1503 (.ZN (n_0_1_821), .A1 (n_0_1_860), .A2 (hfn_ipo_n41));
AOI21_X2 i_0_1_1502 (.ZN (n_0_1_820), .A (n_0_1_821), .B1 (n_0_22), .B2 (hfn_ipo_n41));
INV_X4 i_0_1_1501 (.ZN (\A_imm[23] ), .A (n_0_1_820));
NOR2_X1 i_0_1_1500 (.ZN (n_0_1_819), .A1 (n_0_1_859), .A2 (hfn_ipo_n41));
INV_X4 i_0_1_1498 (.ZN (\A_imm[22] ), .A (n_0_1_818));
NOR2_X1 i_0_1_1497 (.ZN (n_0_1_817), .A1 (n_0_1_858), .A2 (hfn_ipo_n41));
AOI21_X4 i_0_1_1496 (.ZN (sgo__n847), .A (n_0_1_817), .B1 (n_0_20), .B2 (hfn_ipo_n41));
NOR2_X1 i_0_1_1494 (.ZN (n_0_1_815), .A1 (n_0_1_857), .A2 (hfn_ipo_n41));
AOI21_X4 i_0_1_1493 (.ZN (n_0_1_814), .A (n_0_1_815), .B1 (n_0_19), .B2 (hfn_ipo_n41));
CLKBUF_X2 opt_ipo_c6275 (.Z (opt_ipo_n5720), .A (n_0_1_392));
NOR2_X1 i_0_1_1491 (.ZN (n_0_1_813), .A1 (n_0_1_856), .A2 (hfn_ipo_n41));
AOI21_X2 i_0_1_1490 (.ZN (n_0_1_812), .A (n_0_1_813), .B1 (n_0_18), .B2 (hfn_ipo_n41));
NOR2_X1 i_0_1_1488 (.ZN (n_0_1_811), .A1 (n_0_1_855), .A2 (hfn_ipo_n41));
INV_X4 i_0_1_1486 (.ZN (\A_imm[18] ), .A (n_0_1_810));
NOR2_X1 i_0_1_1485 (.ZN (n_0_1_809), .A1 (n_0_1_854), .A2 (hfn_ipo_n41));
NOR2_X1 i_0_1_1482 (.ZN (n_0_1_807), .A1 (n_0_1_853), .A2 (hfn_ipo_n41));
INV_X2 i_0_1_1480 (.ZN (\A_imm[16] ), .A (n_0_1_806));
NOR2_X1 i_0_1_1479 (.ZN (n_0_1_805), .A1 (n_0_1_852), .A2 (hfn_ipo_n41));
NOR2_X1 i_0_1_1476 (.ZN (n_0_1_803), .A1 (n_0_1_851), .A2 (hfn_ipo_n41));
INV_X8 i_0_1_1474 (.ZN (\A_imm[14] ), .A (sgo__n681));
NOR2_X1 i_0_1_1473 (.ZN (n_0_1_801), .A1 (n_0_1_850), .A2 (hfn_ipo_n41));
AOI21_X4 i_0_1_1472 (.ZN (n_0_1_800), .A (n_0_1_801), .B1 (n_0_12), .B2 (hfn_ipo_n41));
INV_X4 i_0_1_1471 (.ZN (\A_imm[13] ), .A (n_0_1_800));
NOR2_X1 i_0_1_1470 (.ZN (n_0_1_799), .A1 (n_0_1_849), .A2 (hfn_ipo_n41));
AOI21_X2 i_0_1_1469 (.ZN (n_0_1_798), .A (n_0_1_799), .B1 (n_0_11), .B2 (hfn_ipo_n41));
INV_X2 i_0_1_1468 (.ZN (\A_imm[12] ), .A (n_0_1_798));
NOR2_X1 i_0_1_1467 (.ZN (n_0_1_797), .A1 (n_0_1_848), .A2 (hfn_ipo_n41));
CLKBUF_X1 CLOCK_slh__c7900 (.Z (CLOCK_slh__n7190), .A (CLOCK_slh__n7189));
NOR2_X1 i_0_1_1464 (.ZN (n_0_1_795), .A1 (n_0_1_847), .A2 (hfn_ipo_n41));
AOI21_X4 i_0_1_1463 (.ZN (n_0_1_794), .A (n_0_1_795), .B1 (n_0_9), .B2 (A_in));
INV_X4 opt_ipo_c6349 (.ZN (opt_ipo_n5794), .A (opt_ipo_n5795));
NOR2_X1 i_0_1_1461 (.ZN (n_0_1_793), .A1 (n_0_1_846), .A2 (A_in));
AOI21_X2 i_0_1_1460 (.ZN (sgo__n1324), .A (n_0_1_793), .B1 (n_0_8), .B2 (A_in));
INV_X16 i_0_1_1459 (.ZN (\A_imm[9] ), .A (n_0_1_792));
NOR2_X1 i_0_1_1458 (.ZN (n_0_1_791), .A1 (n_0_1_845), .A2 (A_in));
AOI21_X4 i_0_1_1457 (.ZN (n_0_1_790), .A (n_0_1_791), .B1 (n_0_7), .B2 (A_in));
BUF_X1 spw__L2_c3_c8539 (.Z (spw__n7739), .A (spw__n7740));
NOR2_X1 i_0_1_1455 (.ZN (n_0_1_789), .A1 (n_0_1_844), .A2 (A_in));
AOI21_X4 i_0_1_1454 (.ZN (n_0_1_788), .A (n_0_1_789), .B1 (n_0_6), .B2 (A_in));
INV_X4 i_0_1_1453 (.ZN (\A_imm[7] ), .A (n_0_1_788));
NOR2_X1 i_0_1_1452 (.ZN (n_0_1_787), .A1 (n_0_1_843), .A2 (A_in));
INV_X8 i_0_1_1450 (.ZN (spw__n7741), .A (n_0_1_786));
NOR2_X1 i_0_1_1446 (.ZN (n_0_1_783), .A1 (n_0_1_841), .A2 (A_in));
AOI21_X4 i_0_1_1445 (.ZN (n_0_1_782), .A (n_0_1_783), .B1 (n_0_3), .B2 (A_in));
INV_X4 i_0_1_1444 (.ZN (\A_imm[4] ), .A (n_0_1_782));
NOR2_X1 i_0_1_1443 (.ZN (n_0_1_781), .A1 (n_0_1_840), .A2 (A_in));
AOI21_X4 i_0_1_1442 (.ZN (sgo__n1116), .A (n_0_1_781), .B1 (n_0_2), .B2 (A_in));
INV_X4 i_0_1_1441 (.ZN (\A_imm[3] ), .A (sgo__n1116));
INV_X2 i_0_1_1433 (.ZN (n_0_1_774), .A (n_0_1_775));
AOI22_X1 i_0_1_1425 (.ZN (n_0_1_768), .A1 (sgo__n1241), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (sgo__n844));
OAI21_X1 i_0_1_1424 (.ZN (n_0_842), .A (n_0_1_768), .B1 (n_0_1_772), .B2 (sgo__n734));
AOI22_X2 i_0_1_1421 (.ZN (n_0_1_766), .A1 (sgo__n877), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (\A_imm_2s_complement[28] ));
OAI21_X2 i_0_1_1420 (.ZN (n_0_840), .A (n_0_1_766), .B1 (n_0_1_772), .B2 (slo__xsl_n1669));
AOI22_X1 i_0_1_1419 (.ZN (n_0_1_765), .A1 (sgo__n943), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (sgo__n877));
OAI21_X1 i_0_1_1418 (.ZN (n_0_839), .A (n_0_1_765), .B1 (n_0_1_772), .B2 (slo__n2762));
AOI22_X1 i_0_1_1417 (.ZN (n_0_1_764), .A1 (\A_imm_2s_complement[25] ), .A2 (n_0_1_771)
    , .B1 (n_0_1_770), .B2 (\A_imm_2s_complement[26] ));
OAI21_X1 i_0_1_1416 (.ZN (n_0_838), .A (n_0_1_764), .B1 (n_0_1_772), .B2 (slo__xsl_n1889));
AOI22_X1 i_0_1_1415 (.ZN (n_0_1_763), .A1 (slo__n1550), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (\A_imm_2s_complement[25] ));
OAI21_X1 i_0_1_1414 (.ZN (n_0_837), .A (n_0_1_763), .B1 (n_0_1_772), .B2 (slo__xsl_n2010));
AOI22_X1 i_0_1_1413 (.ZN (n_0_1_762), .A1 (\A_imm_2s_complement[23] ), .A2 (n_0_1_771)
    , .B1 (n_0_1_770), .B2 (\A_imm_2s_complement[24] ));
OAI21_X1 i_0_1_1412 (.ZN (n_0_836), .A (n_0_1_762), .B1 (n_0_1_772), .B2 (sgo__n1238));
AOI22_X1 i_0_1_1411 (.ZN (n_0_1_761), .A1 (\A_imm_2s_complement[22] ), .A2 (n_0_1_771)
    , .B1 (\A_imm_2s_complement[23] ), .B2 (n_0_1_770));
BUF_X2 slo___L1_c3733 (.Z (slo___n3416), .A (opt_ipo_n5159));
AOI22_X1 i_0_1_1409 (.ZN (n_0_1_760), .A1 (\A_imm_2s_complement[21] ), .A2 (n_0_1_771)
    , .B1 (\A_imm_2s_complement[22] ), .B2 (n_0_1_770));
OAI21_X1 i_0_1_1408 (.ZN (n_0_834), .A (n_0_1_760), .B1 (n_0_1_772), .B2 (slo__xsl_n1641));
AOI22_X1 i_0_1_1407 (.ZN (n_0_1_759), .A1 (opt_ipo_n5339), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (\A_imm_2s_complement[21] ));
OAI21_X1 i_0_1_1406 (.ZN (n_0_833), .A (n_0_1_759), .B1 (n_0_1_772), .B2 (opt_ipo_n5145));
AOI22_X1 i_0_1_1405 (.ZN (n_0_1_758), .A1 (\A_imm_2s_complement[19] ), .A2 (n_0_1_771)
    , .B1 (n_0_1_770), .B2 (opt_ipo_n5785));
OAI21_X1 i_0_1_1404 (.ZN (n_0_832), .A (n_0_1_758), .B1 (n_0_1_772), .B2 (opt_ipo_n5195));
AOI22_X1 i_0_1_1403 (.ZN (n_0_1_757), .A1 (\A_imm_2s_complement[18] ), .A2 (n_0_1_771)
    , .B1 (n_0_1_770), .B2 (opt_ipo_n5373));
OAI21_X1 i_0_1_1402 (.ZN (n_0_831), .A (n_0_1_757), .B1 (n_0_1_772), .B2 (opt_ipo_n5307));
AOI22_X1 i_0_1_1401 (.ZN (n_0_1_756), .A1 (opt_ipo_n5411), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (\A_imm_2s_complement[18] ));
OAI21_X1 i_0_1_1400 (.ZN (n_0_830), .A (n_0_1_756), .B1 (n_0_1_772), .B2 (slo__xsl_n1425));
AOI22_X1 i_0_1_1391 (.ZN (n_0_1_751), .A1 (slo__n1702), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (opt_ipo_n5710));
OAI21_X1 i_0_1_1390 (.ZN (n_0_825), .A (n_0_1_751), .B1 (n_0_1_772), .B2 (slo__n1559));
AOI22_X1 i_0_1_1389 (.ZN (n_0_1_750), .A1 (slo__n3026), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (slo__n1702));
OAI21_X1 i_0_1_1388 (.ZN (n_0_824), .A (n_0_1_750), .B1 (n_0_1_772), .B2 (slo__n1402));
AOI22_X1 i_0_1_1385 (.ZN (n_0_1_748), .A1 (opt_ipo_n5197), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (opt_ipo_n5465));
OAI21_X1 i_0_1_1384 (.ZN (n_0_822), .A (n_0_1_748), .B1 (n_0_1_772), .B2 (opt_ipo_n5165));
AOI22_X1 i_0_1_1383 (.ZN (n_0_1_747), .A1 (slo__n2969), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (opt_ipo_n5197));
OAI21_X1 i_0_1_1382 (.ZN (n_0_821), .A (n_0_1_747), .B1 (n_0_1_772), .B2 (n_0_1_792));
AOI22_X1 i_0_1_1381 (.ZN (n_0_1_746), .A1 (CLOCK_spw__n7292), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (slo__n2969));
OAI21_X1 i_0_1_1380 (.ZN (n_0_820), .A (n_0_1_746), .B1 (n_0_1_772), .B2 (opt_ipo_n5794));
AOI22_X1 i_0_1_1379 (.ZN (n_0_1_745), .A1 (opt_ipo_n5204), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (CLOCK_spw__n7292));
OAI21_X1 i_0_1_1378 (.ZN (n_0_819), .A (n_0_1_745), .B1 (n_0_1_772), .B2 (sgo__n874));
AOI22_X1 i_0_1_1377 (.ZN (n_0_1_744), .A1 (slo__n3910), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (opt_ipo_n5204));
OAI21_X1 i_0_1_1376 (.ZN (n_0_818), .A (n_0_1_744), .B1 (n_0_1_772), .B2 (slo__xsl_n1694));
AOI22_X1 i_0_1_1375 (.ZN (n_0_1_743), .A1 (slo__n2805), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (slo__n3910));
OAI21_X1 i_0_1_1374 (.ZN (n_0_817), .A (n_0_1_743), .B1 (n_0_1_772), .B2 (n_0_1_784));
AOI22_X1 i_0_1_1373 (.ZN (n_0_1_742), .A1 (\A_imm_2s_complement[3] ), .A2 (n_0_1_771)
    , .B1 (n_0_1_770), .B2 (slo__n2805));
OAI21_X1 i_0_1_1372 (.ZN (n_0_816), .A (n_0_1_742), .B1 (n_0_1_772), .B2 (sgo__n959));
AOI22_X1 i_0_1_1371 (.ZN (n_0_1_741), .A1 (\A_imm_2s_complement[2] ), .A2 (n_0_1_771)
    , .B1 (n_0_1_770), .B2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_1370 (.ZN (n_0_815), .A (n_0_1_741), .B1 (n_0_1_772), .B2 (slo__xsl_n3900));
AOI22_X1 i_0_1_1369 (.ZN (n_0_1_740), .A1 (\A_imm_2s_complement[1] ), .A2 (n_0_1_771)
    , .B1 (n_0_1_770), .B2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_1368 (.ZN (n_0_814), .A (n_0_1_740), .B1 (n_0_1_772), .B2 (sgo__n1043));
AOI22_X1 i_0_1_1367 (.ZN (n_0_1_739), .A1 (sgo__n759), .A2 (n_0_1_771), .B1 (n_0_1_770), .B2 (\A_imm_2s_complement[1] ));
AND2_X1 i_0_1_1365 (.ZN (n_0_812), .A1 (n_0_186), .A2 (sgo__n759));
MUX2_X1 i_0_1_1363 (.Z (n_0_1_738), .A (n_0_184), .B (n_0_32), .S (drc_ipo_n58));
NAND2_X1 i_0_1_1362 (.ZN (n_0_1_737), .A1 (n_0_1_775), .A2 (n_0_1_738));
MUX2_X2 i_0_1_1361 (.Z (n_0_1_736), .A (n_0_183), .B (n_0_33), .S (drc_ipo_n58));
INV_X1 i_0_1_1360 (.ZN (n_0_1_735), .A (n_0_1_736));
NAND3_X1 i_0_1_1359 (.ZN (n_0_1_734), .A1 (n_0_1_737), .A2 (n_0_1_736), .A3 (\A_imm_2s_complement[31] ));
OAI21_X1 i_0_1_1358 (.ZN (n_0_1_733), .A (\A_imm[31] ), .B1 (n_0_1_775), .B2 (n_0_1_738));
OAI21_X1 i_0_1_1357 (.ZN (n_0_811), .A (n_0_1_734), .B1 (n_0_1_733), .B2 (n_0_1_736));
XNOR2_X1 i_0_1_1356 (.ZN (n_0_1_732), .A (n_0_1_774), .B (n_0_1_738));
AOI222_X1 i_0_1_1347 (.ZN (n_0_1_725), .A1 (\A_imm_2s_complement[29] ), .A2 (n_0_1_731)
    , .B1 (n_0_1_730), .B2 (\A_imm[28] ), .C1 (n_0_1_728), .C2 (\A_imm_2s_complement[28] ));
OAI21_X1 i_0_1_1346 (.ZN (n_0_808), .A (n_0_1_725), .B1 (n_0_1_729), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_1341 (.ZN (n_0_1_722), .A1 (\A_imm_2s_complement[26] ), .A2 (n_0_1_731)
    , .B1 (n_0_1_730), .B2 (opt_ipo_n5362), .C1 (n_0_1_728), .C2 (\A_imm_2s_complement[25] ));
OAI21_X1 i_0_1_1340 (.ZN (n_0_805), .A (n_0_1_722), .B1 (n_0_1_729), .B2 (slo__xsl_n1889));
AOI222_X1 i_0_1_1339 (.ZN (n_0_1_721), .A1 (\A_imm_2s_complement[25] ), .A2 (n_0_1_731)
    , .B1 (n_0_1_730), .B2 (slo__n2216), .C1 (n_0_1_728), .C2 (\A_imm_2s_complement[24] ));
OAI21_X1 i_0_1_1338 (.ZN (n_0_804), .A (n_0_1_721), .B1 (n_0_1_729), .B2 (slo__xsl_n2010));
AOI222_X2 i_0_1_1337 (.ZN (n_0_1_720), .A1 (\A_imm_2s_complement[24] ), .A2 (n_0_1_731)
    , .B1 (n_0_1_730), .B2 (slo__n3760), .C1 (\A_imm_2s_complement[23] ), .C2 (n_0_1_728));
OAI21_X1 i_0_1_1336 (.ZN (n_0_803), .A (n_0_1_720), .B1 (n_0_1_729), .B2 (sgo__n1238));
AOI222_X2 i_0_1_1335 (.ZN (n_0_1_719), .A1 (sgo__n839), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (slo__n1649), .C1 (n_0_1_728), .C2 (\A_imm_2s_complement[22] ));
OAI21_X1 i_0_1_1334 (.ZN (n_0_802), .A (n_0_1_719), .B1 (n_0_1_729), .B2 (slo__n1812));
AOI222_X1 i_0_1_1331 (.ZN (n_0_1_717), .A1 (\A_imm_2s_complement[21] ), .A2 (n_0_1_731)
    , .B1 (n_0_1_730), .B2 (opt_ipo_n5196), .C1 (n_0_1_728), .C2 (opt_ipo_n5785));
OAI21_X1 i_0_1_1330 (.ZN (n_0_800), .A (n_0_1_717), .B1 (n_0_1_729), .B2 (opt_ipo_n5145));
AOI222_X2 i_0_1_1329 (.ZN (n_0_1_716), .A1 (opt_ipo_n5785), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (opt_ipo_n5303), .C1 (n_0_1_728), .C2 (\A_imm_2s_complement[19] ));
OAI21_X2 i_0_1_1328 (.ZN (n_0_799), .A (n_0_1_716), .B1 (n_0_1_729), .B2 (opt_ipo_n5195));
AOI222_X2 i_0_1_1327 (.ZN (n_0_1_715), .A1 (opt_ipo_n5373), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (slo__n2915), .C1 (n_0_1_728), .C2 (\A_imm_2s_complement[18] ));
OAI21_X1 i_0_1_1326 (.ZN (n_0_798), .A (n_0_1_715), .B1 (n_0_1_729), .B2 (opt_ipo_n5307));
AOI222_X1 i_0_1_1323 (.ZN (n_0_1_713), .A1 (opt_ipo_n5411), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (slo__n3547), .C1 (n_0_1_728), .C2 (opt_ipo_n5162));
OAI21_X1 i_0_1_1322 (.ZN (n_0_796), .A (n_0_1_713), .B1 (n_0_1_729), .B2 (slo__xsl_n1366));
AOI222_X1 i_0_1_1321 (.ZN (n_0_1_712), .A1 (sgo__n1056), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (opt_ipo_n5415), .C1 (n_0_1_728), .C2 (opt_ipo_n5653));
OAI21_X1 i_0_1_1320 (.ZN (n_0_795), .A (n_0_1_712), .B1 (n_0_1_729), .B2 (slo__n1493));
AOI222_X1 i_0_1_1319 (.ZN (n_0_1_711), .A1 (sgo__n895), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (\A_imm[14] ), .C1 (n_0_1_728), .C2 (opt_ipo_n5672));
OAI21_X1 i_0_1_1318 (.ZN (n_0_794), .A (n_0_1_711), .B1 (n_0_1_729), .B2 (slo__n1828));
AOI222_X2 i_0_1_1317 (.ZN (n_0_1_710), .A1 (opt_ipo_n5672), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (\A_imm[13] ), .C1 (n_0_1_728), .C2 (\A_imm_2s_complement[13] ));
OAI21_X2 i_0_1_1316 (.ZN (n_0_793), .A (n_0_1_710), .B1 (n_0_1_729), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_1315 (.ZN (n_0_1_709), .A1 (opt_ipo_n5710), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (slo__n3230), .C1 (n_0_1_728), .C2 (\A_imm_2s_complement[12] ));
OAI21_X1 i_0_1_1314 (.ZN (n_0_792), .A (n_0_1_709), .B1 (n_0_1_729), .B2 (slo__n1559));
AOI222_X1 i_0_1_1313 (.ZN (n_0_1_708), .A1 (slo__n1702), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (opt_ipo_n5297), .C1 (n_0_1_728), .C2 (slo__n3026));
OAI21_X1 i_0_1_1312 (.ZN (n_0_791), .A (n_0_1_708), .B1 (n_0_1_729), .B2 (slo__n1402));
AOI222_X1 i_0_1_1311 (.ZN (n_0_1_707), .A1 (slo__n3026), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (opt_ipo_n5164), .C1 (n_0_1_728), .C2 (opt_ipo_n5466));
OAI21_X1 i_0_1_1310 (.ZN (n_0_790), .A (n_0_1_707), .B1 (n_0_1_729), .B2 (slo___n3458));
AOI222_X2 i_0_1_1309 (.ZN (n_0_1_706), .A1 (opt_ipo_n5466), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (\A_imm[9] ), .C1 (n_0_1_728), .C2 (opt_ipo_n5198));
OAI21_X1 i_0_1_1308 (.ZN (n_0_789), .A (n_0_1_706), .B1 (n_0_1_729), .B2 (opt_ipo_n5165));
AOI222_X2 i_0_1_1307 (.ZN (n_0_1_705), .A1 (opt_ipo_n5198), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (slo__n3281), .C1 (n_0_1_728), .C2 (\A_imm_2s_complement[8] ));
OAI21_X1 i_0_1_1306 (.ZN (n_0_788), .A (n_0_1_705), .B1 (n_0_1_729), .B2 (n_0_1_792));
AOI222_X1 i_0_1_1305 (.ZN (n_0_1_704), .A1 (slo__n2969), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (slo__n1788), .C1 (CLOCK_spw__n7292), .C2 (n_0_1_728));
OAI21_X1 i_0_1_1304 (.ZN (n_0_787), .A (n_0_1_704), .B1 (n_0_1_729), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_1303 (.ZN (n_0_1_703), .A1 (\A_imm_2s_complement[7] ), .A2 (n_0_1_731)
    , .B1 (n_0_1_730), .B2 (spw__n7740), .C1 (n_0_1_728), .C2 (opt_ipo_n5205));
OAI21_X1 i_0_1_1302 (.ZN (n_0_786), .A (n_0_1_703), .B1 (n_0_1_729), .B2 (sgo__n874));
AOI222_X1 i_0_1_1299 (.ZN (n_0_1_701), .A1 (\A_imm_2s_complement[5] ), .A2 (n_0_1_731)
    , .B1 (n_0_1_730), .B2 (sgo__n962), .C1 (\A_imm_2s_complement[4] ), .C2 (n_0_1_728));
OAI21_X1 i_0_1_1298 (.ZN (n_0_784), .A (n_0_1_701), .B1 (n_0_1_729), .B2 (n_0_1_784));
AOI222_X1 i_0_1_1297 (.ZN (n_0_1_700), .A1 (slo__n2805), .A2 (n_0_1_731), .B1 (n_0_1_730)
    , .B2 (slo__n1801), .C1 (n_0_1_728), .C2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_1296 (.ZN (n_0_783), .A (n_0_1_700), .B1 (n_0_1_729), .B2 (sgo__n959));
AOI222_X1 i_0_1_1295 (.ZN (n_0_1_699), .A1 (\A_imm_2s_complement[3] ), .A2 (n_0_1_731)
    , .B1 (n_0_1_730), .B2 (sgo__n1053), .C1 (n_0_1_728), .C2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_1294 (.ZN (n_0_782), .A (n_0_1_699), .B1 (n_0_1_729), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_1293 (.ZN (n_0_1_698), .A1 (\A_imm_2s_complement[2] ), .A2 (n_0_1_731)
    , .B1 (n_0_1_730), .B2 (opt_ipo_n5459), .C1 (n_0_1_728), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_1292 (.ZN (n_0_781), .A (n_0_1_698), .B1 (n_0_1_729), .B2 (sgo__n1043));
NAND2_X1 i_0_1_1291 (.ZN (n_0_1_697), .A1 (\A_imm_2s_complement[1] ), .A2 (n_0_1_731));
OAI21_X1 i_0_1_1290 (.ZN (n_0_1_696), .A (sgo__n759), .B1 (n_0_1_730), .B2 (n_0_1_728));
OAI211_X1 i_0_1_1289 (.ZN (n_0_780), .A (n_0_1_697), .B (n_0_1_696), .C1 (n_0_1_776), .C2 (n_0_1_729));
AND2_X1 i_0_1_1288 (.ZN (n_0_779), .A1 (n_0_1_732), .A2 (sgo__n759));
MUX2_X2 i_0_1_1287 (.Z (n_0_1_695), .A (n_0_182), .B (n_0_34), .S (drc_ipo_n58));
NAND2_X1 i_0_1_1286 (.ZN (n_0_1_694), .A1 (n_0_1_736), .A2 (n_0_1_695));
MUX2_X2 i_0_1_1285 (.Z (n_0_1_693), .A (n_0_181), .B (n_0_35), .S (drc_ipo_n58));
NAND2_X1 CLOCK_slo__sro_c7471 (.ZN (CLOCK_slo__sro_n6740), .A1 (n_0_1_671), .A2 (CLOCK_slo__sro_n6741));
NAND3_X1 i_0_1_1283 (.ZN (n_0_1_691), .A1 (n_0_1_694), .A2 (opt_ipo_n5682), .A3 (\A_imm_2s_complement[31] ));
OAI21_X1 i_0_1_1282 (.ZN (n_0_1_690), .A (\A_imm[31] ), .B1 (n_0_1_736), .B2 (n_0_1_695));
OAI21_X2 i_0_1_1281 (.ZN (n_0_778), .A (n_0_1_691), .B1 (n_0_1_690), .B2 (opt_ipo_n5682));
XNOR2_X2 i_0_1_1280 (.ZN (n_0_1_689), .A (n_0_1_735), .B (n_0_1_695));
AOI222_X1 i_0_1_1275 (.ZN (n_0_1_684), .A1 (sgo__n731), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (\A_imm[30] ), .C1 (opt_ipo_n5278), .C2 (sgo__n844));
OAI21_X1 i_0_1_1274 (.ZN (n_0_777), .A (n_0_1_684), .B1 (n_0_1_686), .B2 (n_0_1_836));
AOI222_X1 i_0_1_1273 (.ZN (n_0_1_683), .A1 (\A_imm_2s_complement[30] ), .A2 (opt_ipo_n5679)
    , .B1 (n_0_1_687), .B2 (\A_imm[29] ), .C1 (opt_ipo_n5278), .C2 (\A_imm_2s_complement[29] ));
OAI21_X1 i_0_1_1272 (.ZN (n_0_776), .A (n_0_1_683), .B1 (n_0_1_686), .B2 (sgo__n734));
AOI222_X1 i_0_1_1271 (.ZN (n_0_1_682), .A1 (\A_imm_2s_complement[29] ), .A2 (opt_ipo_n5679)
    , .B1 (n_0_1_687), .B2 (\A_imm[28] ), .C1 (opt_ipo_n5278), .C2 (\A_imm_2s_complement[28] ));
OAI21_X1 i_0_1_1270 (.ZN (n_0_775), .A (n_0_1_682), .B1 (n_0_1_686), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_1269 (.ZN (n_0_1_681), .A1 (\A_imm_2s_complement[28] ), .A2 (opt_ipo_n5679)
    , .B1 (n_0_1_687), .B2 (\A_imm[27] ), .C1 (\A_imm_2s_complement[27] ), .C2 (opt_ipo_n5278));
OAI21_X1 i_0_1_1268 (.ZN (n_0_774), .A (n_0_1_681), .B1 (n_0_1_686), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_1267 (.ZN (n_0_1_680), .A1 (\A_imm_2s_complement[27] ), .A2 (opt_ipo_n5679)
    , .B1 (n_0_1_687), .B2 (slo__n1897), .C1 (opt_ipo_n5278), .C2 (\A_imm_2s_complement[26] ));
OAI21_X1 i_0_1_1266 (.ZN (n_0_773), .A (n_0_1_680), .B1 (n_0_1_686), .B2 (slo__n2762));
AOI222_X2 i_0_1_1263 (.ZN (n_0_1_678), .A1 (\A_imm_2s_complement[25] ), .A2 (opt_ipo_n5679)
    , .B1 (n_0_1_687), .B2 (slo__n2216), .C1 (opt_ipo_n5278), .C2 (\A_imm_2s_complement[24] ));
OAI21_X1 i_0_1_1262 (.ZN (n_0_771), .A (n_0_1_678), .B1 (n_0_1_686), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_1261 (.ZN (n_0_1_677), .A1 (\A_imm_2s_complement[24] ), .A2 (opt_ipo_n5679)
    , .B1 (n_0_1_687), .B2 (slo__n3760), .C1 (opt_ipo_n5278), .C2 (\A_imm_2s_complement[23] ));
OAI21_X1 i_0_1_1260 (.ZN (n_0_770), .A (n_0_1_677), .B1 (n_0_1_686), .B2 (sgo__n1238));
AOI222_X2 i_0_1_1259 (.ZN (n_0_1_676), .A1 (sgo__n839), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (slo__n1649), .C1 (opt_ipo_n5278), .C2 (sgo__n836));
OAI21_X1 i_0_1_1258 (.ZN (n_0_769), .A (n_0_1_676), .B1 (n_0_1_686), .B2 (slo__n1812));
AOI222_X2 i_0_1_1257 (.ZN (n_0_1_675), .A1 (\A_imm_2s_complement[22] ), .A2 (opt_ipo_n5679)
    , .B1 (n_0_1_687), .B2 (opt_ipo_n5135), .C1 (\A_imm_2s_complement[21] ), .C2 (opt_ipo_n5278));
OAI21_X1 i_0_1_1256 (.ZN (n_0_768), .A (n_0_1_675), .B1 (n_0_1_686), .B2 (slo__xsl_n1641));
AOI222_X1 i_0_1_1255 (.ZN (n_0_1_674), .A1 (sgo__n1009), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (opt_ipo_n5196), .C1 (opt_ipo_n5278), .C2 (opt_ipo_n5785));
OAI21_X1 i_0_1_1254 (.ZN (n_0_767), .A (n_0_1_674), .B1 (n_0_1_686), .B2 (opt_ipo_n5145));
AOI222_X1 i_0_1_1253 (.ZN (n_0_1_673), .A1 (opt_ipo_n5339), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (opt_ipo_n5303), .C1 (opt_ipo_n5278), .C2 (\A_imm_2s_complement[19] ));
OAI21_X1 i_0_1_1252 (.ZN (n_0_766), .A (n_0_1_673), .B1 (n_0_1_686), .B2 (opt_ipo_n5195));
AOI222_X1 i_0_1_1251 (.ZN (n_0_1_672), .A1 (opt_ipo_n5373), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (slo__n2915), .C1 (opt_ipo_n5278), .C2 (\A_imm_2s_complement[18] ));
OAI21_X1 i_0_1_1250 (.ZN (n_0_765), .A (n_0_1_672), .B1 (n_0_1_686), .B2 (opt_ipo_n5307));
AOI222_X1 i_0_1_1249 (.ZN (n_0_1_671), .A1 (\A_imm_2s_complement[18] ), .A2 (opt_ipo_n5679)
    , .B1 (n_0_1_687), .B2 (slo__n3402), .C1 (opt_ipo_n5278), .C2 (CLOCK_opt_ipo_n5880));
OR2_X1 CLOCK_slo__sro_c7553 (.ZN (CLOCK_slo__sro_n6809), .A1 (n_0_1_772), .A2 (slo__n1493));
AOI222_X1 i_0_1_1247 (.ZN (n_0_1_670), .A1 (opt_ipo_n5411), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (slo__n3547), .C1 (\A_imm_2s_complement[16] ), .C2 (opt_ipo_n5278));
OAI21_X1 i_0_1_1246 (.ZN (n_0_763), .A (n_0_1_670), .B1 (n_0_1_686), .B2 (slo__xsl_n1366));
CLKBUF_X1 CLOCK_slh__c7880 (.Z (CLOCK_slh__n7170), .A (CLOCK_slh__n7169));
OAI21_X1 i_0_1_1244 (.ZN (n_0_762), .A (sgo__sro_n905), .B1 (n_0_1_686), .B2 (slo__n1493));
AOI222_X1 i_0_1_1243 (.ZN (n_0_1_668), .A1 (opt_ipo_n5653), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (\A_imm[14] ), .C1 (opt_ipo_n5278), .C2 (opt_ipo_n5672));
OAI21_X1 i_0_1_1242 (.ZN (n_0_761), .A (n_0_1_668), .B1 (n_0_1_686), .B2 (slo__n1828));
AOI222_X1 i_0_1_1241 (.ZN (n_0_1_667), .A1 (slo__n2107), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (\A_imm[13] ), .C1 (opt_ipo_n5278), .C2 (opt_ipo_n5710));
OAI21_X1 i_0_1_1240 (.ZN (n_0_760), .A (n_0_1_667), .B1 (n_0_1_686), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_1239 (.ZN (n_0_1_666), .A1 (opt_ipo_n5710), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (slo__n3230), .C1 (opt_ipo_n5278), .C2 (slo__n1702));
OAI21_X1 i_0_1_1238 (.ZN (n_0_759), .A (n_0_1_666), .B1 (n_0_1_686), .B2 (slo__n1559));
AOI222_X1 i_0_1_1237 (.ZN (n_0_1_665), .A1 (\A_imm_2s_complement[12] ), .A2 (opt_ipo_n5679)
    , .B1 (n_0_1_687), .B2 (opt_ipo_n5297), .C1 (opt_ipo_n5278), .C2 (\A_imm_2s_complement[11] ));
OAI21_X1 i_0_1_1236 (.ZN (n_0_758), .A (n_0_1_665), .B1 (n_0_1_686), .B2 (slo__n1402));
AOI222_X1 i_0_1_1235 (.ZN (n_0_1_664), .A1 (slo__n3026), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (opt_ipo_n5164), .C1 (opt_ipo_n5278), .C2 (opt_ipo_n5466));
OAI21_X1 i_0_1_1234 (.ZN (n_0_757), .A (n_0_1_664), .B1 (n_0_1_686), .B2 (slo___n3458));
AOI222_X1 i_0_1_1233 (.ZN (n_0_1_663), .A1 (opt_ipo_n5465), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (\A_imm[9] ), .C1 (opt_ipo_n5278), .C2 (opt_ipo_n5197));
OAI21_X1 i_0_1_1232 (.ZN (n_0_756), .A (n_0_1_663), .B1 (n_0_1_686), .B2 (opt_ipo_n5165));
AOI222_X2 i_0_1_1231 (.ZN (n_0_1_662), .A1 (opt_ipo_n5197), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (slo__n3281), .C1 (opt_ipo_n5278), .C2 (slo__n2969));
OAI21_X1 i_0_1_1230 (.ZN (n_0_755), .A (n_0_1_662), .B1 (n_0_1_686), .B2 (n_0_1_792));
AOI222_X2 i_0_1_1229 (.ZN (n_0_1_661), .A1 (\A_imm_2s_complement[8] ), .A2 (n_0_1_688)
    , .B1 (n_0_1_687), .B2 (slo__n1788), .C1 (\A_imm_2s_complement[7] ), .C2 (opt_ipo_n5280));
OAI21_X1 i_0_1_1228 (.ZN (n_0_754), .A (n_0_1_661), .B1 (n_0_1_686), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_1227 (.ZN (n_0_1_660), .A1 (\A_imm_2s_complement[7] ), .A2 (opt_ipo_n5679)
    , .B1 (n_0_1_687), .B2 (spw__n7740), .C1 (opt_ipo_n5280), .C2 (opt_ipo_n5205));
OAI21_X1 i_0_1_1226 (.ZN (n_0_753), .A (n_0_1_660), .B1 (n_0_1_686), .B2 (sgo__n874));
AOI222_X1 i_0_1_1225 (.ZN (n_0_1_659), .A1 (opt_ipo_n5204), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (slo__n3378), .C1 (opt_ipo_n5278), .C2 (slo__n3910));
OAI21_X1 i_0_1_1224 (.ZN (n_0_752), .A (n_0_1_659), .B1 (n_0_1_686), .B2 (slo__xsl_n1694));
AOI222_X1 i_0_1_1223 (.ZN (n_0_1_658), .A1 (slo__n3910), .A2 (opt_ipo_n5679), .B1 (n_0_1_687)
    , .B2 (sgo__n962), .C1 (opt_ipo_n5278), .C2 (slo__n2805));
OAI21_X1 i_0_1_1222 (.ZN (n_0_751), .A (n_0_1_658), .B1 (n_0_1_686), .B2 (n_0_1_784));
OAI21_X1 i_0_1_1220 (.ZN (n_0_750), .A (slo__sro_n2333), .B1 (n_0_1_686), .B2 (sgo__n959));
AOI222_X1 i_0_1_1219 (.ZN (n_0_1_656), .A1 (\A_imm_2s_complement[3] ), .A2 (opt_ipo_n5679)
    , .B1 (n_0_1_687), .B2 (sgo__n1053), .C1 (opt_ipo_n5280), .C2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_1218 (.ZN (n_0_749), .A (n_0_1_656), .B1 (n_0_1_686), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_1217 (.ZN (n_0_1_655), .A1 (\A_imm_2s_complement[2] ), .A2 (opt_ipo_n5679)
    , .B1 (n_0_1_687), .B2 (opt_ipo_n5459), .C1 (opt_ipo_n5280), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_1216 (.ZN (n_0_748), .A (n_0_1_655), .B1 (n_0_1_686), .B2 (sgo__n1043));
NAND2_X1 i_0_1_1215 (.ZN (n_0_1_654), .A1 (\A_imm_2s_complement[1] ), .A2 (opt_ipo_n5679));
OAI21_X1 i_0_1_1214 (.ZN (n_0_1_653), .A (sgo__n759), .B1 (n_0_1_687), .B2 (opt_ipo_n5280));
OAI211_X1 i_0_1_1213 (.ZN (n_0_747), .A (n_0_1_654), .B (n_0_1_653), .C1 (n_0_1_776), .C2 (n_0_1_686));
AND2_X1 i_0_1_1212 (.ZN (n_0_746), .A1 (n_0_1_689), .A2 (sgo__n759));
MUX2_X2 i_0_1_1211 (.Z (slo__n1588), .A (n_0_179), .B (n_0_37), .S (drc_ipo_n58));
INV_X2 i_0_1_1210 (.ZN (n_0_1_651), .A (slo__n1588));
MUX2_X2 i_0_1_1209 (.Z (n_0_1_650), .A (n_0_180), .B (n_0_36), .S (drc_ipo_n58));
OAI21_X1 i_0_1_1208 (.ZN (n_0_1_649), .A (\A_imm[31] ), .B1 (opt_ipo_n5682), .B2 (opt_ipo_n5398));
NAND2_X4 i_0_1_1207 (.ZN (n_0_1_648), .A1 (n_0_1_693), .A2 (n_0_1_650));
NAND3_X1 i_0_1_1206 (.ZN (n_0_1_647), .A1 (n_0_1_648), .A2 (\A_imm_2s_complement[31] ), .A3 (opt_ipo_n5152));
OAI21_X1 i_0_1_1205 (.ZN (n_0_745), .A (n_0_1_647), .B1 (n_0_1_649), .B2 (opt_ipo_n5152));
XNOR2_X2 i_0_1_1204 (.ZN (n_0_1_646), .A (opt_ipo_n5683), .B (n_0_1_650));
AOI222_X1 i_0_1_1199 (.ZN (n_0_1_641), .A1 (\A_imm_2s_complement[31] ), .A2 (CLOCK_spw__n7344)
    , .B1 (opt_ipo_n5395), .B2 (\A_imm[30] ), .C1 (opt_ipo_n5393), .C2 (sgo__n844));
OAI21_X1 i_0_1_1198 (.ZN (n_0_744), .A (n_0_1_641), .B1 (n_0_1_643), .B2 (n_0_1_836));
AOI222_X1 i_0_1_1195 (.ZN (n_0_1_639), .A1 (sgo__n1241), .A2 (CLOCK_spw__n7344), .B1 (opt_ipo_n5395)
    , .B2 (\A_imm[28] ), .C1 (opt_ipo_n5393), .C2 (sgo__n678));
OAI21_X1 i_0_1_1194 (.ZN (n_0_742), .A (n_0_1_639), .B1 (n_0_1_643), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_1193 (.ZN (n_0_1_638), .A1 (sgo__n678), .A2 (CLOCK_spw__n7344), .B1 (opt_ipo_n5395)
    , .B2 (\A_imm[27] ), .C1 (opt_ipo_n5393), .C2 (\A_imm_2s_complement[27] ));
OAI21_X1 i_0_1_1192 (.ZN (n_0_741), .A (n_0_1_638), .B1 (n_0_1_643), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_1191 (.ZN (n_0_1_637), .A1 (\A_imm_2s_complement[27] ), .A2 (CLOCK_spw__n7344)
    , .B1 (opt_ipo_n5395), .B2 (slo__n1897), .C1 (opt_ipo_n5393), .C2 (\A_imm_2s_complement[26] ));
OAI21_X1 i_0_1_1190 (.ZN (n_0_740), .A (n_0_1_637), .B1 (n_0_1_643), .B2 (slo__n2762));
AOI222_X1 i_0_1_1187 (.ZN (n_0_1_635), .A1 (sgo__n1339), .A2 (CLOCK_spw__n7344), .B1 (opt_ipo_n5395)
    , .B2 (slo__n2216), .C1 (opt_ipo_n5393), .C2 (\A_imm_2s_complement[24] ));
OAI21_X1 i_0_1_1186 (.ZN (n_0_738), .A (n_0_1_635), .B1 (n_0_1_643), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_1185 (.ZN (n_0_1_634), .A1 (\A_imm_2s_complement[24] ), .A2 (CLOCK_spw__n7344)
    , .B1 (opt_ipo_n5395), .B2 (slo__n3760), .C1 (\A_imm_2s_complement[23] ), .C2 (opt_ipo_n5393));
OAI21_X1 i_0_1_1184 (.ZN (n_0_737), .A (n_0_1_634), .B1 (n_0_1_643), .B2 (sgo__n1238));
AOI222_X2 i_0_1_1183 (.ZN (n_0_1_633), .A1 (sgo__n839), .A2 (CLOCK_spw__n7344), .B1 (opt_ipo_n5395)
    , .B2 (slo__n1649), .C1 (opt_ipo_n5393), .C2 (\A_imm_2s_complement[22] ));
OAI21_X1 i_0_1_1182 (.ZN (n_0_736), .A (n_0_1_633), .B1 (n_0_1_643), .B2 (slo__n1812));
AOI222_X1 i_0_1_1181 (.ZN (n_0_1_632), .A1 (sgo__n836), .A2 (CLOCK_spw__n7344), .B1 (opt_ipo_n5395)
    , .B2 (opt_ipo_n5135), .C1 (opt_ipo_n5393), .C2 (\A_imm_2s_complement[21] ));
OAI21_X1 i_0_1_1180 (.ZN (n_0_735), .A (n_0_1_632), .B1 (n_0_1_643), .B2 (slo__xsl_n1641));
AOI222_X1 i_0_1_1179 (.ZN (n_0_1_631), .A1 (sgo__n1009), .A2 (CLOCK_spw__n7344), .B1 (opt_ipo_n5395)
    , .B2 (opt_ipo_n5196), .C1 (opt_ipo_n5393), .C2 (opt_ipo_n5339));
OAI21_X1 i_0_1_1178 (.ZN (n_0_734), .A (n_0_1_631), .B1 (n_0_1_643), .B2 (opt_ipo_n5145));
AOI222_X2 i_0_1_1177 (.ZN (n_0_1_630), .A1 (opt_ipo_n5785), .A2 (CLOCK_spw__n7344)
    , .B1 (opt_ipo_n5395), .B2 (opt_ipo_n5303), .C1 (opt_ipo_n5393), .C2 (\A_imm_2s_complement[19] ));
OAI21_X1 i_0_1_1176 (.ZN (n_0_733), .A (n_0_1_630), .B1 (n_0_1_643), .B2 (opt_ipo_n5195));
AOI222_X1 i_0_1_1175 (.ZN (n_0_1_629), .A1 (opt_ipo_n5373), .A2 (CLOCK_spw__n7344)
    , .B1 (opt_ipo_n5395), .B2 (slo__n2915), .C1 (opt_ipo_n5393), .C2 (\A_imm_2s_complement[18] ));
OAI21_X1 i_0_1_1174 (.ZN (n_0_732), .A (n_0_1_629), .B1 (n_0_1_643), .B2 (opt_ipo_n5307));
AOI222_X1 i_0_1_1173 (.ZN (n_0_1_628), .A1 (\A_imm_2s_complement[18] ), .A2 (CLOCK_spw__n7344)
    , .B1 (opt_ipo_n5395), .B2 (slo__n3402), .C1 (opt_ipo_n5393), .C2 (CLOCK_opt_ipo_n5880));
OAI21_X1 i_0_1_1172 (.ZN (n_0_731), .A (n_0_1_628), .B1 (n_0_1_643), .B2 (slo__xsl_n1425));
AOI222_X1 i_0_1_1171 (.ZN (n_0_1_627), .A1 (opt_ipo_n5411), .A2 (CLOCK_spw__n7344)
    , .B1 (opt_ipo_n5395), .B2 (slo__n3547), .C1 (opt_ipo_n5393), .C2 (opt_ipo_n5162));
OAI21_X1 i_0_1_1170 (.ZN (n_0_730), .A (n_0_1_627), .B1 (n_0_1_643), .B2 (slo__xsl_n1366));
AOI222_X2 i_0_1_1169 (.ZN (n_0_1_626), .A1 (opt_ipo_n5162), .A2 (n_0_1_645), .B1 (opt_ipo_n5395)
    , .B2 (opt_ipo_n5415), .C1 (opt_ipo_n5393), .C2 (opt_ipo_n5653));
OAI21_X1 i_0_1_1168 (.ZN (n_0_729), .A (n_0_1_626), .B1 (n_0_1_643), .B2 (slo__n1493));
AOI222_X1 i_0_1_1167 (.ZN (n_0_1_625), .A1 (sgo__n895), .A2 (n_0_1_645), .B1 (opt_ipo_n5395)
    , .B2 (\A_imm[14] ), .C1 (opt_ipo_n5393), .C2 (\A_imm_2s_complement[14] ));
OAI21_X1 i_0_1_1166 (.ZN (n_0_728), .A (n_0_1_625), .B1 (n_0_1_643), .B2 (slo__n1828));
AOI222_X1 i_0_1_1165 (.ZN (n_0_1_624), .A1 (\A_imm_2s_complement[14] ), .A2 (n_0_1_645)
    , .B1 (opt_ipo_n5395), .B2 (\A_imm[13] ), .C1 (\A_imm_2s_complement[13] ), .C2 (n_0_1_642));
OAI21_X1 i_0_1_1164 (.ZN (n_0_727), .A (n_0_1_624), .B1 (n_0_1_643), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_1163 (.ZN (n_0_1_623), .A1 (opt_ipo_n5710), .A2 (n_0_1_645), .B1 (opt_ipo_n5395)
    , .B2 (slo__n3230), .C1 (opt_ipo_n5393), .C2 (\A_imm_2s_complement[12] ));
OAI21_X1 i_0_1_1162 (.ZN (n_0_726), .A (n_0_1_623), .B1 (n_0_1_643), .B2 (slo__n1559));
AOI222_X1 i_0_1_1161 (.ZN (n_0_1_622), .A1 (slo__n1702), .A2 (n_0_1_645), .B1 (opt_ipo_n5395)
    , .B2 (opt_ipo_n5297), .C1 (opt_ipo_n5393), .C2 (slo__n3026));
OAI21_X1 i_0_1_1160 (.ZN (n_0_725), .A (n_0_1_622), .B1 (n_0_1_643), .B2 (slo__n1402));
AOI222_X1 i_0_1_1159 (.ZN (n_0_1_621), .A1 (slo__n3026), .A2 (n_0_1_645), .B1 (opt_ipo_n5395)
    , .B2 (opt_ipo_n5164), .C1 (opt_ipo_n5393), .C2 (opt_ipo_n5465));
OAI21_X1 i_0_1_1158 (.ZN (n_0_724), .A (n_0_1_621), .B1 (n_0_1_643), .B2 (slo___n3458));
AOI222_X1 i_0_1_1157 (.ZN (n_0_1_620), .A1 (opt_ipo_n5466), .A2 (n_0_1_645), .B1 (opt_ipo_n5395)
    , .B2 (\A_imm[9] ), .C1 (opt_ipo_n5393), .C2 (opt_ipo_n5198));
OAI21_X1 i_0_1_1156 (.ZN (n_0_723), .A (n_0_1_620), .B1 (n_0_1_643), .B2 (opt_ipo_n5165));
AOI222_X1 i_0_1_1155 (.ZN (n_0_1_619), .A1 (opt_ipo_n5197), .A2 (n_0_1_645), .B1 (opt_ipo_n5395)
    , .B2 (slo__n3281), .C1 (opt_ipo_n5393), .C2 (slo__n2969));
OAI21_X1 i_0_1_1154 (.ZN (n_0_722), .A (n_0_1_619), .B1 (n_0_1_643), .B2 (n_0_1_792));
AOI222_X1 i_0_1_1153 (.ZN (n_0_1_618), .A1 (slo__n2969), .A2 (n_0_1_645), .B1 (opt_ipo_n5395)
    , .B2 (slo__n1788), .C1 (opt_ipo_n5393), .C2 (CLOCK_spw__n7291));
OAI21_X1 i_0_1_1152 (.ZN (n_0_721), .A (n_0_1_618), .B1 (n_0_1_643), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_1151 (.ZN (n_0_1_617), .A1 (CLOCK_spw__n7291), .A2 (n_0_1_645), .B1 (opt_ipo_n5395)
    , .B2 (\A_imm[6] ), .C1 (opt_ipo_n5393), .C2 (opt_ipo_n5205));
OAI21_X1 i_0_1_1150 (.ZN (n_0_720), .A (n_0_1_617), .B1 (n_0_1_643), .B2 (sgo__n874));
AOI222_X1 i_0_1_1149 (.ZN (n_0_1_616), .A1 (n_0_1_645), .A2 (opt_ipo_n5205), .B1 (opt_ipo_n5395)
    , .B2 (slo__n3378), .C1 (n_0_1_642), .C2 (\A_imm_2s_complement[5] ));
OAI21_X1 i_0_1_1148 (.ZN (n_0_719), .A (n_0_1_616), .B1 (n_0_1_643), .B2 (slo__xsl_n1694));
AOI222_X1 i_0_1_1147 (.ZN (n_0_1_615), .A1 (slo__n3910), .A2 (n_0_1_645), .B1 (opt_ipo_n5395)
    , .B2 (sgo__n962), .C1 (n_0_1_642), .C2 (\A_imm_2s_complement[4] ));
OAI21_X1 i_0_1_1146 (.ZN (n_0_718), .A (n_0_1_615), .B1 (n_0_1_643), .B2 (n_0_1_784));
AOI222_X1 i_0_1_1145 (.ZN (n_0_1_614), .A1 (slo__n2805), .A2 (n_0_1_645), .B1 (opt_ipo_n5395)
    , .B2 (slo__n1801), .C1 (opt_ipo_n5393), .C2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_1144 (.ZN (n_0_717), .A (n_0_1_614), .B1 (n_0_1_643), .B2 (sgo__n959));
AOI222_X1 i_0_1_1143 (.ZN (n_0_1_613), .A1 (\A_imm_2s_complement[3] ), .A2 (n_0_1_645)
    , .B1 (opt_ipo_n5395), .B2 (sgo__n1053), .C1 (opt_ipo_n5393), .C2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_1142 (.ZN (n_0_716), .A (n_0_1_613), .B1 (n_0_1_643), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_1141 (.ZN (n_0_1_612), .A1 (\A_imm_2s_complement[2] ), .A2 (n_0_1_645)
    , .B1 (opt_ipo_n5395), .B2 (opt_ipo_n5459), .C1 (n_0_1_642), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_1140 (.ZN (n_0_715), .A (n_0_1_612), .B1 (n_0_1_643), .B2 (sgo__n1043));
NAND2_X1 i_0_1_1139 (.ZN (n_0_1_611), .A1 (\A_imm_2s_complement[1] ), .A2 (n_0_1_645));
OAI21_X1 i_0_1_1138 (.ZN (n_0_1_610), .A (sgo__n759), .B1 (opt_ipo_n5395), .B2 (opt_ipo_n5393));
OAI211_X1 i_0_1_1137 (.ZN (n_0_714), .A (n_0_1_611), .B (n_0_1_610), .C1 (n_0_1_776), .C2 (n_0_1_643));
AND2_X1 i_0_1_1136 (.ZN (n_0_713), .A1 (n_0_1_646), .A2 (sgo__n759));
MUX2_X2 i_0_1_1135 (.Z (n_0_1_609), .A (n_0_178), .B (n_0_38), .S (drc_ipo_n58));
NAND2_X1 i_0_1_1134 (.ZN (n_0_1_608), .A1 (n_0_1_609), .A2 (slo__n1588));
CLKBUF_X1 CLOCK_slh__c7912 (.Z (CLOCK_slh__n7202), .A (CLOCK_slh__n7201));
NAND3_X1 i_0_1_1131 (.ZN (n_0_1_605), .A1 (n_0_1_608), .A2 (opt_ipo_n5314), .A3 (\A_imm_2s_complement[31] ));
OAI21_X1 i_0_1_1130 (.ZN (n_0_1_604), .A (\A_imm[31] ), .B1 (opt_ipo_n5152), .B2 (n_0_1_609));
OAI21_X1 i_0_1_1129 (.ZN (n_0_712), .A (n_0_1_605), .B1 (n_0_1_604), .B2 (opt_ipo_n5314));
XNOR2_X1 i_0_1_1128 (.ZN (n_0_1_603), .A (n_0_1_651), .B (n_0_1_609));
AOI222_X1 i_0_1_1123 (.ZN (n_0_1_598), .A1 (sgo__n731), .A2 (slo__n4931), .B1 (opt_ipo_n5311)
    , .B2 (\A_imm[30] ), .C1 (spw__n7778), .C2 (sgo__n844));
OAI21_X1 i_0_1_1122 (.ZN (n_0_711), .A (n_0_1_598), .B1 (n_0_1_600), .B2 (n_0_1_836));
AOI222_X1 i_0_1_1119 (.ZN (n_0_1_596), .A1 (sgo__n1241), .A2 (slo__n4931), .B1 (opt_ipo_n5311)
    , .B2 (\A_imm[28] ), .C1 (spw__n7778), .C2 (sgo__n678));
OAI21_X1 i_0_1_1118 (.ZN (n_0_709), .A (n_0_1_596), .B1 (n_0_1_600), .B2 (slo__xsl_n1736));
CLKBUF_X2 slo__c3594 (.Z (slo__n3281), .A (opt_ipo_n5795));
OAI21_X1 i_0_1_1116 (.ZN (n_0_708), .A (slo__sro_n3243), .B1 (n_0_1_600), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_1115 (.ZN (n_0_1_594), .A1 (\A_imm_2s_complement[27] ), .A2 (slo__n4931)
    , .B1 (opt_ipo_n5311), .B2 (slo__n1897), .C1 (\A_imm_2s_complement[26] ), .C2 (spw__n7777));
OAI21_X1 i_0_1_1114 (.ZN (n_0_707), .A (n_0_1_594), .B1 (n_0_1_600), .B2 (slo__n2762));
AOI222_X1 i_0_1_1113 (.ZN (n_0_1_593), .A1 (sgo__n943), .A2 (slo__n4931), .B1 (opt_ipo_n5311)
    , .B2 (opt_ipo_n5362), .C1 (slo__n3614), .C2 (\A_imm_2s_complement[25] ));
OAI21_X1 i_0_1_1112 (.ZN (n_0_706), .A (n_0_1_593), .B1 (n_0_1_600), .B2 (slo__xsl_n1889));
AOI222_X1 i_0_1_1111 (.ZN (n_0_1_592), .A1 (sgo__n1339), .A2 (slo__n4931), .B1 (opt_ipo_n5311)
    , .B2 (slo__n2216), .C1 (spw__n7777), .C2 (\A_imm_2s_complement[24] ));
OAI21_X1 i_0_1_1110 (.ZN (n_0_705), .A (n_0_1_592), .B1 (n_0_1_600), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_1109 (.ZN (n_0_1_591), .A1 (\A_imm_2s_complement[24] ), .A2 (slo__n4931)
    , .B1 (opt_ipo_n5311), .B2 (slo__n3760), .C1 (\A_imm_2s_complement[23] ), .C2 (spw__n7777));
OAI21_X1 i_0_1_1108 (.ZN (n_0_704), .A (n_0_1_591), .B1 (n_0_1_600), .B2 (sgo__n1238));
AOI222_X1 i_0_1_1107 (.ZN (n_0_1_590), .A1 (sgo__n839), .A2 (slo__n4931), .B1 (opt_ipo_n5311)
    , .B2 (slo__n1649), .C1 (n_0_1_599), .C2 (\A_imm_2s_complement[22] ));
OAI21_X1 i_0_1_1106 (.ZN (n_0_703), .A (n_0_1_590), .B1 (n_0_1_600), .B2 (slo__n1812));
AOI222_X1 i_0_1_1103 (.ZN (n_0_1_588), .A1 (\A_imm_2s_complement[21] ), .A2 (slo__n4931)
    , .B1 (opt_ipo_n5312), .B2 (opt_ipo_n5196), .C1 (opt_ipo_n5785), .C2 (n_0_1_599));
OAI21_X1 i_0_1_1102 (.ZN (n_0_701), .A (n_0_1_588), .B1 (n_0_1_600), .B2 (opt_ipo_n5145));
AOI222_X1 i_0_1_1101 (.ZN (n_0_1_587), .A1 (opt_ipo_n5339), .A2 (slo__n4931), .B1 (opt_ipo_n5311)
    , .B2 (opt_ipo_n5303), .C1 (spw__n7776), .C2 (opt_ipo_n5373));
OAI21_X1 i_0_1_1100 (.ZN (n_0_700), .A (n_0_1_587), .B1 (n_0_1_600), .B2 (opt_ipo_n5195));
AOI222_X2 i_0_1_1099 (.ZN (n_0_1_586), .A1 (opt_ipo_n5373), .A2 (slo__n4931), .B1 (opt_ipo_n5312)
    , .B2 (slo__n2915), .C1 (spw__n7776), .C2 (\A_imm_2s_complement[18] ));
OAI21_X1 i_0_1_1098 (.ZN (n_0_699), .A (n_0_1_586), .B1 (n_0_1_600), .B2 (opt_ipo_n5307));
AOI222_X2 i_0_1_1097 (.ZN (n_0_1_585), .A1 (\A_imm_2s_complement[18] ), .A2 (slo__n4931)
    , .B1 (opt_ipo_n5312), .B2 (slo__n3402), .C1 (CLOCK_opt_ipo_n5880), .C2 (n_0_1_599));
OAI21_X1 i_0_1_1096 (.ZN (n_0_698), .A (n_0_1_585), .B1 (n_0_1_600), .B2 (slo__xsl_n1425));
AOI222_X2 i_0_1_1095 (.ZN (n_0_1_584), .A1 (opt_ipo_n5411), .A2 (slo__n4931), .B1 (opt_ipo_n5311)
    , .B2 (slo__n3547), .C1 (n_0_1_599), .C2 (\A_imm_2s_complement[16] ));
OAI21_X1 i_0_1_1094 (.ZN (n_0_697), .A (n_0_1_584), .B1 (n_0_1_600), .B2 (slo__xsl_n1366));
AOI222_X1 i_0_1_1093 (.ZN (n_0_1_583), .A1 (opt_ipo_n5162), .A2 (opt_ipo_n5151), .B1 (opt_ipo_n5312)
    , .B2 (opt_ipo_n5415), .C1 (n_0_1_599), .C2 (\A_imm_2s_complement[15] ));
OAI21_X1 i_0_1_1092 (.ZN (n_0_696), .A (n_0_1_583), .B1 (n_0_1_600), .B2 (slo__n1493));
AOI222_X1 i_0_1_1091 (.ZN (n_0_1_582), .A1 (sgo__n895), .A2 (opt_ipo_n5151), .B1 (opt_ipo_n5311)
    , .B2 (\A_imm[14] ), .C1 (n_0_1_599), .C2 (opt_ipo_n5672));
OAI21_X1 i_0_1_1090 (.ZN (n_0_695), .A (n_0_1_582), .B1 (n_0_1_600), .B2 (slo__n1828));
AOI222_X1 i_0_1_1089 (.ZN (n_0_1_581), .A1 (\A_imm_2s_complement[14] ), .A2 (opt_ipo_n5151)
    , .B1 (opt_ipo_n5312), .B2 (\A_imm[13] ), .C1 (\A_imm_2s_complement[13] ), .C2 (slo__n3030));
OAI21_X1 i_0_1_1088 (.ZN (n_0_694), .A (n_0_1_581), .B1 (n_0_1_600), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_1087 (.ZN (n_0_1_580), .A1 (opt_ipo_n5710), .A2 (opt_ipo_n5151), .B1 (opt_ipo_n5311)
    , .B2 (slo__n3230), .C1 (n_0_1_599), .C2 (\A_imm_2s_complement[12] ));
OAI21_X1 i_0_1_1086 (.ZN (n_0_693), .A (n_0_1_580), .B1 (n_0_1_600), .B2 (slo__n1559));
AOI222_X1 i_0_1_1085 (.ZN (n_0_1_579), .A1 (\A_imm_2s_complement[12] ), .A2 (n_0_1_920)
    , .B1 (opt_ipo_n5312), .B2 (opt_ipo_n5297), .C1 (\A_imm_2s_complement[11] ), .C2 (n_0_1_599));
OAI21_X1 i_0_1_1084 (.ZN (n_0_692), .A (n_0_1_579), .B1 (n_0_1_600), .B2 (slo__n1402));
AOI222_X1 i_0_1_1083 (.ZN (n_0_1_578), .A1 (slo__n3026), .A2 (opt_ipo_n5151), .B1 (opt_ipo_n5311)
    , .B2 (opt_ipo_n5164), .C1 (n_0_1_599), .C2 (opt_ipo_n5466));
OAI21_X1 i_0_1_1082 (.ZN (n_0_691), .A (n_0_1_578), .B1 (n_0_1_600), .B2 (slo___n3458));
AOI222_X1 i_0_1_1081 (.ZN (n_0_1_577), .A1 (opt_ipo_n5466), .A2 (opt_ipo_n5151), .B1 (opt_ipo_n5312)
    , .B2 (\A_imm[9] ), .C1 (slo__n3030), .C2 (opt_ipo_n5198));
BUF_X4 slo__c1796 (.Z (slo__n1615), .A (n_0_1_167));
AOI222_X1 i_0_1_1079 (.ZN (n_0_1_576), .A1 (opt_ipo_n5197), .A2 (opt_ipo_n5151), .B1 (opt_ipo_n5312)
    , .B2 (slo__n3281), .C1 (n_0_1_599), .C2 (\A_imm_2s_complement[8] ));
OAI21_X1 i_0_1_1078 (.ZN (n_0_689), .A (n_0_1_576), .B1 (n_0_1_600), .B2 (n_0_1_792));
AOI222_X1 i_0_1_1077 (.ZN (n_0_1_575), .A1 (\A_imm_2s_complement[8] ), .A2 (opt_ipo_n5151)
    , .B1 (opt_ipo_n5312), .B2 (slo__n1788), .C1 (slo__n3614), .C2 (\A_imm_2s_complement[7] ));
OAI21_X1 i_0_1_1076 (.ZN (n_0_688), .A (n_0_1_575), .B1 (n_0_1_600), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_1075 (.ZN (n_0_1_574), .A1 (CLOCK_spw__n7291), .A2 (opt_ipo_n5151)
    , .B1 (opt_ipo_n5311), .B2 (\A_imm[6] ), .C1 (slo__n3614), .C2 (opt_ipo_n5205));
OAI21_X1 i_0_1_1074 (.ZN (n_0_687), .A (n_0_1_574), .B1 (n_0_1_600), .B2 (sgo__n874));
AOI222_X1 i_0_1_1073 (.ZN (n_0_1_573), .A1 (opt_ipo_n5205), .A2 (n_0_1_920), .B1 (opt_ipo_n5312)
    , .B2 (slo__n3378), .C1 (n_0_1_599), .C2 (\A_imm_2s_complement[5] ));
OAI21_X1 i_0_1_1072 (.ZN (n_0_686), .A (n_0_1_573), .B1 (n_0_1_600), .B2 (slo__xsl_n1694));
NAND2_X1 slo__sro_c3687 (.ZN (slo__sro_n3370), .A1 (n_0_1_969), .A2 (n_0_1_842));
OAI21_X1 i_0_1_1070 (.ZN (n_0_685), .A (slo__sro_n3317), .B1 (n_0_1_600), .B2 (n_0_1_784));
AOI222_X2 i_0_1_1069 (.ZN (n_0_1_571), .A1 (n_0_1_920), .A2 (slo__n2805), .B1 (opt_ipo_n5312)
    , .B2 (slo__n1801), .C1 (slo__n3030), .C2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_1068 (.ZN (n_0_684), .A (n_0_1_571), .B1 (n_0_1_600), .B2 (sgo__n959));
AOI222_X1 i_0_1_1067 (.ZN (n_0_1_570), .A1 (\A_imm_2s_complement[3] ), .A2 (n_0_1_920)
    , .B1 (opt_ipo_n5312), .B2 (sgo__n1053), .C1 (n_0_1_599), .C2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_1066 (.ZN (n_0_683), .A (n_0_1_570), .B1 (n_0_1_600), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_1065 (.ZN (n_0_1_569), .A1 (\A_imm_2s_complement[2] ), .A2 (opt_ipo_n5151)
    , .B1 (opt_ipo_n5312), .B2 (opt_ipo_n5459), .C1 (n_0_1_599), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_1064 (.ZN (n_0_682), .A (n_0_1_569), .B1 (n_0_1_600), .B2 (sgo__n1043));
NAND2_X1 i_0_1_1063 (.ZN (n_0_1_568), .A1 (\A_imm_2s_complement[1] ), .A2 (opt_ipo_n5151));
OAI21_X1 i_0_1_1062 (.ZN (n_0_1_567), .A (sgo__n759), .B1 (opt_ipo_n5311), .B2 (n_0_1_599));
OAI211_X1 i_0_1_1061 (.ZN (n_0_681), .A (n_0_1_568), .B (n_0_1_567), .C1 (n_0_1_776), .C2 (n_0_1_600));
AND2_X1 i_0_1_1060 (.ZN (n_0_680), .A1 (n_0_1_603), .A2 (sgo__n759));
MUX2_X2 i_0_1_1059 (.Z (n_0_1_566), .A (n_0_175), .B (n_0_41), .S (drc_ipo_n58));
INV_X2 i_0_1_1058 (.ZN (n_0_1_565), .A (n_0_1_566));
CLKBUF_X1 slo___L1_c3387 (.Z (slo___n3078), .A (n_0_1_259));
OAI21_X1 i_0_1_1056 (.ZN (n_0_1_563), .A (\A_imm[31] ), .B1 (opt_ipo_n5314), .B2 (slo__sro_n2959));
NAND2_X1 i_0_1_1055 (.ZN (n_0_1_562), .A1 (n_0_1_607), .A2 (slo__sro_n2959));
NAND3_X1 i_0_1_1054 (.ZN (n_0_1_561), .A1 (n_0_1_562), .A2 (\A_imm_2s_complement[31] ), .A3 (n_0_1_566));
OAI21_X2 i_0_1_1053 (.ZN (n_0_679), .A (n_0_1_561), .B1 (n_0_1_563), .B2 (slo___n3489));
XNOR2_X1 i_0_1_1052 (.ZN (n_0_1_560), .A (opt_ipo_n5315), .B (slo__sro_n2959));
AOI222_X1 i_0_1_1043 (.ZN (n_0_1_553), .A1 (sgo__n1241), .A2 (slo___n2464), .B1 (opt_ipo_n5774)
    , .B2 (\A_imm[28] ), .C1 (opt_ipo_n5258), .C2 (sgo__n678));
OAI21_X1 i_0_1_1042 (.ZN (n_0_676), .A (n_0_1_553), .B1 (n_0_1_557), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_1041 (.ZN (n_0_1_552), .A1 (sgo__n678), .A2 (slo___n2464), .B1 (opt_ipo_n5774)
    , .B2 (\A_imm[27] ), .C1 (\A_imm_2s_complement[27] ), .C2 (opt_ipo_n5258));
OAI21_X1 i_0_1_1040 (.ZN (n_0_675), .A (n_0_1_552), .B1 (n_0_1_557), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_1039 (.ZN (n_0_1_551), .A1 (sgo__n877), .A2 (slo___n2464), .B1 (opt_ipo_n5774)
    , .B2 (slo__n1897), .C1 (opt_ipo_n5258), .C2 (\A_imm_2s_complement[26] ));
OAI21_X1 i_0_1_1038 (.ZN (n_0_674), .A (n_0_1_551), .B1 (n_0_1_557), .B2 (slo__n2762));
BUF_X4 slo__c3332 (.Z (slo__n3026), .A (\A_imm_2s_complement[11] ));
OAI21_X1 i_0_1_1036 (.ZN (n_0_673), .A (slo__sro_n2992), .B1 (n_0_1_557), .B2 (slo__xsl_n1889));
AOI222_X2 i_0_1_1035 (.ZN (n_0_1_549), .A1 (sgo__n1339), .A2 (slo___n2464), .B1 (opt_ipo_n5774)
    , .B2 (slo__n2216), .C1 (opt_ipo_n5258), .C2 (\A_imm_2s_complement[24] ));
OAI21_X1 i_0_1_1034 (.ZN (n_0_672), .A (n_0_1_549), .B1 (n_0_1_557), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_1033 (.ZN (n_0_1_548), .A1 (slo__n1550), .A2 (slo___n2464), .B1 (opt_ipo_n5774)
    , .B2 (slo__n3760), .C1 (opt_ipo_n5258), .C2 (sgo__n839));
OAI21_X1 i_0_1_1032 (.ZN (n_0_671), .A (n_0_1_548), .B1 (n_0_1_557), .B2 (sgo__n1238));
AOI222_X1 i_0_1_1031 (.ZN (n_0_1_547), .A1 (sgo__n839), .A2 (slo___n2464), .B1 (opt_ipo_n5774)
    , .B2 (slo__n1649), .C1 (opt_ipo_n5258), .C2 (sgo__n836));
OAI21_X1 i_0_1_1030 (.ZN (n_0_670), .A (n_0_1_547), .B1 (n_0_1_557), .B2 (slo__n1812));
AOI222_X1 i_0_1_1029 (.ZN (n_0_1_546), .A1 (\A_imm_2s_complement[22] ), .A2 (slo___n2464)
    , .B1 (opt_ipo_n5423), .B2 (opt_ipo_n5135), .C1 (\A_imm_2s_complement[21] ), .C2 (opt_ipo_n5258));
OAI21_X1 i_0_1_1028 (.ZN (n_0_669), .A (n_0_1_546), .B1 (n_0_1_557), .B2 (slo__xsl_n1641));
AOI222_X2 i_0_1_1027 (.ZN (n_0_1_545), .A1 (sgo__n1009), .A2 (slo___n2464), .B1 (opt_ipo_n5774)
    , .B2 (opt_ipo_n5196), .C1 (opt_ipo_n5258), .C2 (opt_ipo_n5339));
OAI21_X1 i_0_1_1026 (.ZN (n_0_668), .A (n_0_1_545), .B1 (n_0_1_557), .B2 (opt_ipo_n5145));
INV_X1 opt_ipo_c6237 (.ZN (opt_ipo_n5682), .A (opt_ipo_n5683));
OAI21_X2 i_0_1_1024 (.ZN (n_0_667), .A (n_0_1_544), .B1 (n_0_1_557), .B2 (opt_ipo_n5195));
AOI222_X2 i_0_1_1023 (.ZN (n_0_1_543), .A1 (\A_imm_2s_complement[19] ), .A2 (slo___n2464)
    , .B1 (opt_ipo_n5774), .B2 (slo__n2915), .C1 (\A_imm_2s_complement[18] ), .C2 (opt_ipo_n5258));
OAI21_X1 i_0_1_1022 (.ZN (n_0_666), .A (n_0_1_543), .B1 (n_0_1_557), .B2 (opt_ipo_n5307));
AOI222_X1 i_0_1_1021 (.ZN (n_0_1_542), .A1 (\A_imm_2s_complement[18] ), .A2 (slo___n2464)
    , .B1 (opt_ipo_n5774), .B2 (slo__n3402), .C1 (opt_ipo_n5258), .C2 (opt_ipo_n5411));
OAI21_X1 i_0_1_1020 (.ZN (n_0_665), .A (n_0_1_542), .B1 (n_0_1_557), .B2 (slo__xsl_n1425));
AOI222_X1 i_0_1_1019 (.ZN (n_0_1_541), .A1 (opt_ipo_n5411), .A2 (slo__n3696), .B1 (opt_ipo_n5423)
    , .B2 (slo__n3547), .C1 (\A_imm_2s_complement[16] ), .C2 (opt_ipo_n5258));
OAI21_X1 i_0_1_1018 (.ZN (n_0_664), .A (n_0_1_541), .B1 (n_0_1_557), .B2 (slo__xsl_n1366));
AOI222_X1 i_0_1_1017 (.ZN (n_0_1_540), .A1 (\A_imm_2s_complement[16] ), .A2 (slo__n3696)
    , .B1 (opt_ipo_n5423), .B2 (opt_ipo_n5415), .C1 (opt_ipo_n5258), .C2 (\A_imm_2s_complement[15] ));
OAI21_X1 i_0_1_1016 (.ZN (n_0_663), .A (n_0_1_540), .B1 (n_0_1_557), .B2 (slo__n1493));
AOI222_X1 i_0_1_1015 (.ZN (n_0_1_539), .A1 (sgo__n895), .A2 (slo___n2464), .B1 (opt_ipo_n5774)
    , .B2 (\A_imm[14] ), .C1 (opt_ipo_n5258), .C2 (\A_imm_2s_complement[14] ));
OAI21_X1 i_0_1_1014 (.ZN (n_0_662), .A (n_0_1_539), .B1 (n_0_1_557), .B2 (slo__n1828));
AOI222_X1 i_0_1_1013 (.ZN (n_0_1_538), .A1 (opt_ipo_n5672), .A2 (opt_ipo_n5438), .B1 (opt_ipo_n5774)
    , .B2 (\A_imm[13] ), .C1 (opt_ipo_n5258), .C2 (\A_imm_2s_complement[13] ));
OAI21_X1 i_0_1_1012 (.ZN (n_0_661), .A (n_0_1_538), .B1 (n_0_1_557), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_1011 (.ZN (n_0_1_537), .A1 (opt_ipo_n5710), .A2 (opt_ipo_n5438), .B1 (opt_ipo_n5774)
    , .B2 (slo__n3230), .C1 (opt_ipo_n5258), .C2 (\A_imm_2s_complement[12] ));
OAI21_X1 i_0_1_1010 (.ZN (n_0_660), .A (n_0_1_537), .B1 (n_0_1_557), .B2 (slo__n1559));
AOI222_X1 i_0_1_1009 (.ZN (n_0_1_536), .A1 (\A_imm_2s_complement[12] ), .A2 (opt_ipo_n5438)
    , .B1 (opt_ipo_n5423), .B2 (opt_ipo_n5297), .C1 (opt_ipo_n5258), .C2 (\A_imm_2s_complement[11] ));
OAI21_X1 i_0_1_1008 (.ZN (n_0_659), .A (n_0_1_536), .B1 (n_0_1_557), .B2 (slo__n1402));
AOI222_X1 i_0_1_1007 (.ZN (n_0_1_535), .A1 (slo__n3026), .A2 (opt_ipo_n5438), .B1 (opt_ipo_n5774)
    , .B2 (opt_ipo_n5164), .C1 (opt_ipo_n5258), .C2 (opt_ipo_n5466));
OAI21_X1 i_0_1_1006 (.ZN (n_0_658), .A (n_0_1_535), .B1 (n_0_1_557), .B2 (slo___n3458));
AOI222_X1 i_0_1_1005 (.ZN (n_0_1_534), .A1 (opt_ipo_n5466), .A2 (opt_ipo_n5438), .B1 (opt_ipo_n5423)
    , .B2 (\A_imm[9] ), .C1 (slo__n4197), .C2 (opt_ipo_n5198));
OAI21_X1 i_0_1_1004 (.ZN (n_0_657), .A (n_0_1_534), .B1 (n_0_1_557), .B2 (opt_ipo_n5165));
AOI222_X1 i_0_1_1003 (.ZN (n_0_1_533), .A1 (opt_ipo_n5197), .A2 (opt_ipo_n5438), .B1 (opt_ipo_n5774)
    , .B2 (slo__n3281), .C1 (opt_ipo_n5258), .C2 (\A_imm_2s_complement[8] ));
OAI21_X1 i_0_1_1002 (.ZN (n_0_656), .A (n_0_1_533), .B1 (n_0_1_557), .B2 (n_0_1_792));
INV_X2 opt_ipo_c6258 (.ZN (opt_ipo_n5703), .A (n_0_149));
OAI21_X1 i_0_1_1000 (.ZN (n_0_655), .A (slo__sro_n2477), .B1 (n_0_1_557), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_999 (.ZN (n_0_1_531), .A1 (\A_imm_2s_complement[7] ), .A2 (opt_ipo_n5438)
    , .B1 (opt_ipo_n5423), .B2 (\A_imm[6] ), .C1 (opt_ipo_n5258), .C2 (opt_ipo_n5205));
OAI21_X1 i_0_1_998 (.ZN (n_0_654), .A (n_0_1_531), .B1 (n_0_1_557), .B2 (sgo__n874));
AOI222_X2 i_0_1_997 (.ZN (n_0_1_530), .A1 (opt_ipo_n5205), .A2 (opt_ipo_n5438), .B1 (opt_ipo_n5774)
    , .B2 (slo__n3378), .C1 (opt_ipo_n5258), .C2 (\A_imm_2s_complement[5] ));
OAI21_X1 i_0_1_996 (.ZN (n_0_653), .A (n_0_1_530), .B1 (n_0_1_557), .B2 (slo__xsl_n1694));
AOI222_X1 i_0_1_995 (.ZN (n_0_1_529), .A1 (slo__n3910), .A2 (opt_ipo_n5438), .B1 (opt_ipo_n5774)
    , .B2 (sgo__n962), .C1 (opt_ipo_n5258), .C2 (slo__n2805));
OAI21_X1 i_0_1_994 (.ZN (n_0_652), .A (n_0_1_529), .B1 (n_0_1_557), .B2 (n_0_1_784));
AOI222_X1 i_0_1_993 (.ZN (n_0_1_528), .A1 (slo__n2805), .A2 (n_0_1_559), .B1 (n_0_1_558)
    , .B2 (slo__n1801), .C1 (slo__n4197), .C2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_992 (.ZN (n_0_651), .A (n_0_1_528), .B1 (n_0_1_557), .B2 (sgo__n959));
AOI222_X1 i_0_1_991 (.ZN (n_0_1_527), .A1 (\A_imm_2s_complement[3] ), .A2 (n_0_1_559)
    , .B1 (n_0_1_558), .B2 (sgo__n1053), .C1 (slo__n4197), .C2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_990 (.ZN (n_0_650), .A (n_0_1_527), .B1 (n_0_1_557), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_989 (.ZN (n_0_1_526), .A1 (\A_imm_2s_complement[2] ), .A2 (n_0_1_559)
    , .B1 (n_0_1_558), .B2 (opt_ipo_n5459), .C1 (slo__n4197), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_988 (.ZN (n_0_649), .A (n_0_1_526), .B1 (n_0_1_557), .B2 (sgo__n1043));
NAND2_X1 i_0_1_987 (.ZN (n_0_1_525), .A1 (\A_imm_2s_complement[1] ), .A2 (opt_ipo_n5438));
OAI21_X1 i_0_1_986 (.ZN (n_0_1_524), .A (sgo__n759), .B1 (opt_ipo_n5423), .B2 (opt_ipo_n5258));
OAI211_X1 i_0_1_985 (.ZN (n_0_648), .A (n_0_1_525), .B (n_0_1_524), .C1 (n_0_1_776), .C2 (n_0_1_557));
AND2_X1 i_0_1_984 (.ZN (n_0_647), .A1 (n_0_1_560), .A2 (sgo__n759));
MUX2_X2 i_0_1_983 (.Z (n_0_1_523), .A (n_0_173), .B (n_0_43), .S (drc_ipo_n58));
INV_X4 i_0_1_982 (.ZN (n_0_1_522), .A (n_0_1_523));
MUX2_X1 i_0_1_981 (.Z (n_0_1_521), .A (n_0_174), .B (n_0_42), .S (drc_ipo_n58));
OAI21_X1 i_0_1_980 (.ZN (n_0_1_520), .A (\A_imm[31] ), .B1 (slo___n3489), .B2 (n_0_1_521));
NAND2_X1 i_0_1_979 (.ZN (n_0_1_519), .A1 (slo___n3489), .A2 (n_0_1_521));
NAND3_X1 i_0_1_978 (.ZN (n_0_1_518), .A1 (n_0_1_519), .A2 (\A_imm_2s_complement[31] ), .A3 (n_0_1_523));
OAI21_X1 i_0_1_977 (.ZN (n_0_646), .A (n_0_1_518), .B1 (n_0_1_520), .B2 (n_0_1_523));
XNOR2_X1 i_0_1_976 (.ZN (n_0_1_517), .A (n_0_1_565), .B (n_0_1_521));
AND2_X4 i_0_1_975 (.ZN (n_0_1_516), .A1 (slo__n3522), .A2 (n_0_1_523));
BUF_X2 slo___L1_c2747 (.Z (slo___n2464), .A (slo__n3696));
NAND2_X4 i_0_1_973 (.ZN (n_0_1_514), .A1 (n_0_1_517), .A2 (n_0_1_522));
NOR3_X1 i_0_1_972 (.ZN (n_0_1_513), .A1 (slo___n3489), .A2 (n_0_1_521), .A3 (n_0_1_522));
AOI222_X1 i_0_1_971 (.ZN (n_0_1_512), .A1 (sgo__n731), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (\A_imm[30] ), .C1 (CLOCK_spw__n7329), .C2 (sgo__n844));
OAI21_X1 i_0_1_970 (.ZN (n_0_645), .A (n_0_1_512), .B1 (n_0_1_514), .B2 (n_0_1_836));
AOI222_X1 i_0_1_969 (.ZN (n_0_1_511), .A1 (\A_imm_2s_complement[30] ), .A2 (n_0_1_516)
    , .B1 (slo__mro_n1860), .B2 (\A_imm[29] ), .C1 (CLOCK_spw__n7329), .C2 (\A_imm_2s_complement[29] ));
OAI21_X1 i_0_1_968 (.ZN (n_0_644), .A (n_0_1_511), .B1 (n_0_1_514), .B2 (sgo__n734));
AOI222_X1 i_0_1_967 (.ZN (n_0_1_510), .A1 (\A_imm_2s_complement[29] ), .A2 (n_0_1_516)
    , .B1 (slo__mro_n1860), .B2 (\A_imm[28] ), .C1 (\A_imm_2s_complement[28] ), .C2 (CLOCK_spw__n7329));
OAI21_X1 i_0_1_966 (.ZN (n_0_643), .A (n_0_1_510), .B1 (n_0_1_514), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_965 (.ZN (n_0_1_509), .A1 (sgo__n678), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (\A_imm[27] ), .C1 (CLOCK_spw__n7329), .C2 (\A_imm_2s_complement[27] ));
OAI21_X1 i_0_1_964 (.ZN (n_0_642), .A (n_0_1_509), .B1 (n_0_1_514), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_963 (.ZN (n_0_1_508), .A1 (sgo__n877), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (slo__n1897), .C1 (CLOCK_spw__n7329), .C2 (sgo__n943));
OAI21_X1 i_0_1_962 (.ZN (n_0_641), .A (n_0_1_508), .B1 (n_0_1_514), .B2 (slo__n2762));
AOI222_X1 i_0_1_961 (.ZN (n_0_1_507), .A1 (sgo__n943), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (opt_ipo_n5362), .C1 (CLOCK_spw__n7329), .C2 (\A_imm_2s_complement[25] ));
OAI21_X1 i_0_1_960 (.ZN (n_0_640), .A (n_0_1_507), .B1 (n_0_1_514), .B2 (slo__xsl_n1889));
AOI222_X1 i_0_1_959 (.ZN (n_0_1_506), .A1 (sgo__n1339), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (slo__n2216), .C1 (drc_ipo_n52), .C2 (slo__n1550));
OAI21_X1 i_0_1_958 (.ZN (n_0_639), .A (n_0_1_506), .B1 (n_0_1_514), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_957 (.ZN (n_0_1_505), .A1 (\A_imm_2s_complement[24] ), .A2 (n_0_1_516)
    , .B1 (slo__mro_n1860), .B2 (slo__n3760), .C1 (CLOCK_spw__n7329), .C2 (\A_imm_2s_complement[23] ));
OAI21_X1 i_0_1_956 (.ZN (n_0_638), .A (n_0_1_505), .B1 (n_0_1_514), .B2 (sgo__n1238));
AOI222_X1 i_0_1_955 (.ZN (n_0_1_504), .A1 (sgo__n839), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (slo__n1649), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[22] ));
OAI21_X1 i_0_1_954 (.ZN (n_0_637), .A (n_0_1_504), .B1 (n_0_1_514), .B2 (slo__n1812));
AOI222_X1 i_0_1_953 (.ZN (n_0_1_503), .A1 (sgo__n836), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (opt_ipo_n5135), .C1 (CLOCK_spw__n7329), .C2 (sgo__n1009));
OAI21_X1 i_0_1_952 (.ZN (n_0_636), .A (n_0_1_503), .B1 (n_0_1_514), .B2 (slo__xsl_n1641));
AOI222_X1 i_0_1_951 (.ZN (n_0_1_502), .A1 (\A_imm_2s_complement[21] ), .A2 (n_0_1_516)
    , .B1 (slo__mro_n1860), .B2 (opt_ipo_n5196), .C1 (opt_ipo_n5785), .C2 (drc_ipo_n52));
OAI21_X1 i_0_1_950 (.ZN (n_0_635), .A (n_0_1_502), .B1 (n_0_1_514), .B2 (opt_ipo_n5145));
AOI222_X1 i_0_1_949 (.ZN (n_0_1_501), .A1 (opt_ipo_n5339), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (opt_ipo_n5303), .C1 (\A_imm_2s_complement[19] ), .C2 (drc_ipo_n52));
OAI21_X1 i_0_1_948 (.ZN (n_0_634), .A (n_0_1_501), .B1 (n_0_1_514), .B2 (opt_ipo_n5195));
AOI222_X1 i_0_1_947 (.ZN (n_0_1_500), .A1 (opt_ipo_n5373), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (slo__n2915), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[18] ));
OAI21_X1 i_0_1_946 (.ZN (n_0_633), .A (n_0_1_500), .B1 (n_0_1_514), .B2 (opt_ipo_n5307));
AOI222_X2 i_0_1_945 (.ZN (n_0_1_499), .A1 (\A_imm_2s_complement[18] ), .A2 (n_0_1_516)
    , .B1 (slo__mro_n1860), .B2 (slo__n3402), .C1 (CLOCK_opt_ipo_n5880), .C2 (drc_ipo_n52));
OAI21_X1 i_0_1_944 (.ZN (n_0_632), .A (n_0_1_499), .B1 (n_0_1_514), .B2 (slo__xsl_n1425));
AOI222_X1 i_0_1_943 (.ZN (n_0_1_498), .A1 (opt_ipo_n5411), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (slo__n3547), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[16] ));
OAI21_X1 i_0_1_942 (.ZN (n_0_631), .A (n_0_1_498), .B1 (n_0_1_514), .B2 (slo__xsl_n1366));
AOI222_X1 i_0_1_941 (.ZN (n_0_1_497), .A1 (sgo__n1056), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (opt_ipo_n5415), .C1 (drc_ipo_n52), .C2 (sgo__n895));
OAI21_X1 i_0_1_940 (.ZN (n_0_630), .A (n_0_1_497), .B1 (n_0_1_514), .B2 (slo__n1493));
AOI222_X1 i_0_1_939 (.ZN (n_0_1_496), .A1 (sgo__n895), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (\A_imm[14] ), .C1 (\A_imm_2s_complement[14] ), .C2 (drc_ipo_n52));
OAI21_X1 i_0_1_938 (.ZN (n_0_629), .A (n_0_1_496), .B1 (n_0_1_514), .B2 (slo__n1828));
AOI222_X2 i_0_1_937 (.ZN (n_0_1_495), .A1 (\A_imm_2s_complement[14] ), .A2 (n_0_1_516)
    , .B1 (slo__mro_n1860), .B2 (\A_imm[13] ), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[13] ));
OAI21_X1 i_0_1_936 (.ZN (n_0_628), .A (n_0_1_495), .B1 (n_0_1_514), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_935 (.ZN (n_0_1_494), .A1 (opt_ipo_n5710), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (slo__n3230), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[12] ));
OAI21_X1 i_0_1_934 (.ZN (n_0_627), .A (n_0_1_494), .B1 (n_0_1_514), .B2 (slo__n1559));
AOI222_X1 i_0_1_933 (.ZN (n_0_1_493), .A1 (slo__n1702), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (opt_ipo_n5297), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[11] ));
OAI21_X1 i_0_1_932 (.ZN (n_0_626), .A (n_0_1_493), .B1 (n_0_1_514), .B2 (slo__n1402));
AOI222_X1 i_0_1_931 (.ZN (n_0_1_492), .A1 (slo__n3026), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (opt_ipo_n5164), .C1 (drc_ipo_n52), .C2 (opt_ipo_n5466));
OAI21_X1 i_0_1_930 (.ZN (n_0_625), .A (n_0_1_492), .B1 (n_0_1_514), .B2 (slo___n3458));
AOI222_X1 i_0_1_929 (.ZN (n_0_1_491), .A1 (opt_ipo_n5466), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (\A_imm[9] ), .C1 (drc_ipo_n52), .C2 (opt_ipo_n5198));
OAI21_X1 i_0_1_928 (.ZN (n_0_624), .A (n_0_1_491), .B1 (n_0_1_514), .B2 (opt_ipo_n5165));
AOI222_X1 i_0_1_927 (.ZN (n_0_1_490), .A1 (opt_ipo_n5197), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (slo__n3281), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[8] ));
OAI21_X1 i_0_1_926 (.ZN (n_0_623), .A (n_0_1_490), .B1 (n_0_1_514), .B2 (n_0_1_792));
AOI222_X1 i_0_1_925 (.ZN (n_0_1_489), .A1 (\A_imm_2s_complement[8] ), .A2 (n_0_1_516)
    , .B1 (slo__mro_n1860), .B2 (slo__n1788), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[7] ));
OAI21_X1 i_0_1_924 (.ZN (n_0_622), .A (n_0_1_489), .B1 (n_0_1_514), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_923 (.ZN (n_0_1_488), .A1 (CLOCK_spw__n7291), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (\A_imm[6] ), .C1 (drc_ipo_n52), .C2 (opt_ipo_n5204));
OAI21_X1 i_0_1_922 (.ZN (n_0_621), .A (n_0_1_488), .B1 (n_0_1_514), .B2 (sgo__n874));
AOI222_X1 i_0_1_921 (.ZN (n_0_1_487), .A1 (n_0_1_516), .A2 (opt_ipo_n5205), .B1 (slo__mro_n1860)
    , .B2 (slo__n3378), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[5] ));
OAI21_X1 i_0_1_920 (.ZN (n_0_620), .A (n_0_1_487), .B1 (n_0_1_514), .B2 (slo__xsl_n1694));
AOI222_X1 i_0_1_919 (.ZN (n_0_1_486), .A1 (\A_imm_2s_complement[5] ), .A2 (n_0_1_516)
    , .B1 (slo__mro_n1860), .B2 (sgo__n962), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[4] ));
OAI21_X1 i_0_1_918 (.ZN (n_0_619), .A (n_0_1_486), .B1 (n_0_1_514), .B2 (n_0_1_784));
AOI222_X1 i_0_1_917 (.ZN (n_0_1_485), .A1 (slo__n2805), .A2 (n_0_1_516), .B1 (slo__mro_n1860)
    , .B2 (slo__n1801), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_916 (.ZN (n_0_618), .A (n_0_1_485), .B1 (n_0_1_514), .B2 (sgo__n959));
AOI222_X1 i_0_1_915 (.ZN (n_0_1_484), .A1 (\A_imm_2s_complement[3] ), .A2 (n_0_1_516)
    , .B1 (slo__mro_n1860), .B2 (sgo__n1053), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_914 (.ZN (n_0_617), .A (n_0_1_484), .B1 (n_0_1_514), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_913 (.ZN (n_0_1_483), .A1 (n_0_1_516), .A2 (\A_imm_2s_complement[2] )
    , .B1 (slo__mro_n1860), .B2 (opt_ipo_n5459), .C1 (drc_ipo_n52), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_912 (.ZN (n_0_616), .A (n_0_1_483), .B1 (n_0_1_514), .B2 (sgo__n1043));
NAND2_X1 i_0_1_911 (.ZN (n_0_1_482), .A1 (\A_imm_2s_complement[1] ), .A2 (n_0_1_516));
OAI21_X1 i_0_1_910 (.ZN (n_0_1_481), .A (sgo__n759), .B1 (slo__mro_n1860), .B2 (drc_ipo_n52));
OAI211_X1 i_0_1_909 (.ZN (n_0_615), .A (n_0_1_482), .B (n_0_1_481), .C1 (n_0_1_776), .C2 (n_0_1_514));
AND2_X1 i_0_1_908 (.ZN (n_0_614), .A1 (n_0_1_517), .A2 (sgo__n759));
MUX2_X2 i_0_1_907 (.Z (n_0_1_480), .A (n_0_172), .B (n_0_44), .S (drc_ipo_n58));
NAND2_X2 i_0_1_906 (.ZN (n_0_1_479), .A1 (slo__n3640), .A2 (n_0_1_480));
MUX2_X2 i_0_1_905 (.Z (n_0_1_478), .A (n_0_171), .B (opt_ipo_n5223), .S (drc_ipo_n58));
INV_X2 i_0_1_904 (.ZN (n_0_1_477), .A (n_0_1_478));
NAND3_X1 i_0_1_903 (.ZN (n_0_1_476), .A1 (n_0_1_479), .A2 (slo__xsl_n1963), .A3 (\A_imm_2s_complement[31] ));
OAI21_X1 i_0_1_902 (.ZN (n_0_1_475), .A (\A_imm[31] ), .B1 (slo__n3640), .B2 (n_0_1_480));
OAI21_X2 i_0_1_901 (.ZN (n_0_613), .A (n_0_1_476), .B1 (n_0_1_475), .B2 (slo__xsl_n1963));
XNOR2_X1 i_0_1_900 (.ZN (n_0_1_474), .A (n_0_1_522), .B (n_0_1_480));
CLKBUF_X1 CLOCK_slh__c7905 (.Z (CLOCK_slh__n7195), .A (CLOCK_slh__n7194));
NOR2_X2 i_0_1_898 (.ZN (n_0_1_472), .A1 (n_0_1_479), .A2 (slo__xsl_n1963));
NAND2_X4 i_0_1_897 (.ZN (n_0_1_471), .A1 (n_0_1_474), .A2 (n_0_1_477));
NOR3_X4 i_0_1_896 (.ZN (n_0_1_470), .A1 (slo__n2885), .A2 (n_0_1_477), .A3 (n_0_1_480));
AOI222_X1 i_0_1_895 (.ZN (n_0_1_469), .A1 (sgo__n731), .A2 (spw__n7730), .B1 (slo___n2245)
    , .B2 (\A_imm[30] ), .C1 (drc_ipo_n53), .C2 (sgo__n844));
OAI21_X1 i_0_1_894 (.ZN (n_0_612), .A (n_0_1_469), .B1 (n_0_1_471), .B2 (n_0_1_836));
AOI222_X1 i_0_1_893 (.ZN (n_0_1_468), .A1 (sgo__n844), .A2 (spw__n7730), .B1 (slo___n2245)
    , .B2 (\A_imm[29] ), .C1 (drc_ipo_n53), .C2 (sgo__n1241));
OAI21_X1 i_0_1_892 (.ZN (n_0_611), .A (n_0_1_468), .B1 (n_0_1_471), .B2 (sgo__n734));
AOI222_X1 i_0_1_891 (.ZN (n_0_1_467), .A1 (sgo__n1241), .A2 (spw__n7730), .B1 (slo___n2245)
    , .B2 (\A_imm[28] ), .C1 (drc_ipo_n53), .C2 (sgo__n678));
OAI21_X1 i_0_1_890 (.ZN (n_0_610), .A (n_0_1_467), .B1 (n_0_1_471), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_889 (.ZN (n_0_1_466), .A1 (\A_imm_2s_complement[28] ), .A2 (spw__n7730)
    , .B1 (slo___n2245), .B2 (\A_imm[27] ), .C1 (drc_ipo_n53), .C2 (\A_imm_2s_complement[27] ));
OAI21_X1 i_0_1_888 (.ZN (n_0_609), .A (n_0_1_466), .B1 (n_0_1_471), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_887 (.ZN (n_0_1_465), .A1 (\A_imm_2s_complement[27] ), .A2 (spw__n7729)
    , .B1 (slo___n2245), .B2 (slo__n1897), .C1 (\A_imm_2s_complement[26] ), .C2 (drc_ipo_n53));
OAI21_X1 i_0_1_886 (.ZN (n_0_608), .A (n_0_1_465), .B1 (n_0_1_471), .B2 (slo__n2762));
AOI222_X1 i_0_1_885 (.ZN (n_0_1_464), .A1 (sgo__n943), .A2 (spw__n7729), .B1 (slo___n2245)
    , .B2 (opt_ipo_n5362), .C1 (drc_ipo_n53), .C2 (\A_imm_2s_complement[25] ));
OAI21_X1 i_0_1_884 (.ZN (n_0_607), .A (n_0_1_464), .B1 (n_0_1_471), .B2 (slo__xsl_n1889));
AOI222_X1 i_0_1_883 (.ZN (n_0_1_463), .A1 (sgo__n1339), .A2 (spw__n7729), .B1 (slo___n2245)
    , .B2 (slo__n2216), .C1 (drc_ipo_n53), .C2 (slo__n1550));
OAI21_X1 i_0_1_882 (.ZN (n_0_606), .A (n_0_1_463), .B1 (n_0_1_471), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_881 (.ZN (n_0_1_462), .A1 (slo__n1550), .A2 (spw__n7730), .B1 (slo___n2245)
    , .B2 (slo__n3760), .C1 (drc_ipo_n53), .C2 (sgo__n839));
OAI21_X1 i_0_1_880 (.ZN (n_0_605), .A (n_0_1_462), .B1 (n_0_1_471), .B2 (sgo__n1238));
AOI222_X1 i_0_1_879 (.ZN (n_0_1_461), .A1 (sgo__n839), .A2 (spw__n7729), .B1 (slo___n2245)
    , .B2 (slo__n1649), .C1 (drc_ipo_n53), .C2 (sgo__n836));
OAI21_X1 i_0_1_878 (.ZN (n_0_604), .A (n_0_1_461), .B1 (n_0_1_471), .B2 (slo__n1812));
AOI222_X1 i_0_1_877 (.ZN (n_0_1_460), .A1 (sgo__n836), .A2 (spw__n7729), .B1 (slo___n2245)
    , .B2 (opt_ipo_n5135), .C1 (drc_ipo_n53), .C2 (\A_imm_2s_complement[21] ));
OAI21_X1 i_0_1_876 (.ZN (n_0_603), .A (n_0_1_460), .B1 (n_0_1_471), .B2 (slo__xsl_n1641));
AOI222_X1 i_0_1_875 (.ZN (n_0_1_459), .A1 (sgo__n1009), .A2 (opt_ipo_n5285), .B1 (slo___n2245)
    , .B2 (opt_ipo_n5196), .C1 (drc_ipo_n53), .C2 (opt_ipo_n5785));
OAI21_X1 i_0_1_874 (.ZN (n_0_602), .A (n_0_1_459), .B1 (n_0_1_471), .B2 (opt_ipo_n5145));
AOI222_X1 i_0_1_873 (.ZN (n_0_1_458), .A1 (opt_ipo_n5339), .A2 (spw__n7729), .B1 (slo___n2245)
    , .B2 (opt_ipo_n5303), .C1 (drc_ipo_n53), .C2 (opt_ipo_n5373));
OAI21_X1 i_0_1_872 (.ZN (n_0_601), .A (n_0_1_458), .B1 (n_0_1_471), .B2 (opt_ipo_n5195));
AOI222_X2 i_0_1_871 (.ZN (n_0_1_457), .A1 (opt_ipo_n5373), .A2 (opt_ipo_n5285), .B1 (slo___n2245)
    , .B2 (slo__n2915), .C1 (drc_ipo_n53), .C2 (\A_imm_2s_complement[18] ));
OAI21_X1 i_0_1_870 (.ZN (n_0_600), .A (n_0_1_457), .B1 (n_0_1_471), .B2 (opt_ipo_n5307));
AOI222_X1 i_0_1_869 (.ZN (n_0_1_456), .A1 (\A_imm_2s_complement[18] ), .A2 (opt_ipo_n5285)
    , .B1 (slo___n2244), .B2 (slo__n3402), .C1 (CLOCK_opt_ipo_n5880), .C2 (drc_ipo_n53));
OAI21_X1 i_0_1_868 (.ZN (n_0_599), .A (n_0_1_456), .B1 (n_0_1_471), .B2 (slo__xsl_n1425));
AOI222_X1 i_0_1_867 (.ZN (n_0_1_455), .A1 (opt_ipo_n5411), .A2 (opt_ipo_n5285), .B1 (slo___n2244)
    , .B2 (slo__n3547), .C1 (drc_ipo_n53), .C2 (\A_imm_2s_complement[16] ));
OAI21_X1 i_0_1_866 (.ZN (n_0_598), .A (n_0_1_455), .B1 (n_0_1_471), .B2 (slo__xsl_n1366));
AOI222_X1 i_0_1_865 (.ZN (n_0_1_454), .A1 (\A_imm_2s_complement[16] ), .A2 (n_0_1_473)
    , .B1 (slo___n2244), .B2 (opt_ipo_n5415), .C1 (\A_imm_2s_complement[15] ), .C2 (drc_ipo_n53));
OAI21_X1 i_0_1_864 (.ZN (n_0_597), .A (n_0_1_454), .B1 (n_0_1_471), .B2 (slo__n1493));
AOI222_X1 i_0_1_863 (.ZN (n_0_1_453), .A1 (sgo__n895), .A2 (opt_ipo_n5285), .B1 (slo___n2244)
    , .B2 (\A_imm[14] ), .C1 (drc_ipo_n53), .C2 (\A_imm_2s_complement[14] ));
OAI21_X1 i_0_1_862 (.ZN (n_0_596), .A (n_0_1_453), .B1 (n_0_1_471), .B2 (slo__n1828));
AOI222_X1 i_0_1_861 (.ZN (n_0_1_452), .A1 (slo__n2107), .A2 (opt_ipo_n5285), .B1 (slo___n2244)
    , .B2 (\A_imm[13] ), .C1 (drc_ipo_n53), .C2 (\A_imm_2s_complement[13] ));
OAI21_X1 i_0_1_860 (.ZN (n_0_595), .A (n_0_1_452), .B1 (n_0_1_471), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_859 (.ZN (n_0_1_451), .A1 (opt_ipo_n5710), .A2 (n_0_1_473), .B1 (slo___n2244)
    , .B2 (slo__n3230), .C1 (\A_imm_2s_complement[12] ), .C2 (drc_ipo_n53));
OAI21_X1 i_0_1_858 (.ZN (n_0_594), .A (n_0_1_451), .B1 (n_0_1_471), .B2 (slo__n1559));
AOI222_X2 i_0_1_857 (.ZN (n_0_1_450), .A1 (\A_imm_2s_complement[12] ), .A2 (opt_ipo_n5285)
    , .B1 (slo___n2244), .B2 (opt_ipo_n5297), .C1 (drc_ipo_n53), .C2 (\A_imm_2s_complement[11] ));
OAI21_X1 i_0_1_856 (.ZN (n_0_593), .A (n_0_1_450), .B1 (n_0_1_471), .B2 (slo__n1402));
AOI222_X1 i_0_1_855 (.ZN (n_0_1_449), .A1 (slo__n3026), .A2 (opt_ipo_n5285), .B1 (slo___n2244)
    , .B2 (opt_ipo_n5164), .C1 (drc_ipo_n53), .C2 (opt_ipo_n5466));
OAI21_X1 i_0_1_854 (.ZN (n_0_592), .A (n_0_1_449), .B1 (n_0_1_471), .B2 (slo___n3458));
AOI222_X1 i_0_1_853 (.ZN (n_0_1_448), .A1 (opt_ipo_n5466), .A2 (opt_ipo_n5285), .B1 (n_0_1_472)
    , .B2 (\A_imm[9] ), .C1 (drc_ipo_n53), .C2 (opt_ipo_n5198));
OAI21_X1 i_0_1_852 (.ZN (n_0_591), .A (n_0_1_448), .B1 (n_0_1_471), .B2 (opt_ipo_n5165));
AOI222_X1 i_0_1_851 (.ZN (n_0_1_447), .A1 (opt_ipo_n5197), .A2 (n_0_1_473), .B1 (slo___n2248)
    , .B2 (slo__n3281), .C1 (\A_imm_2s_complement[8] ), .C2 (drc_ipo_n53));
OAI21_X1 i_0_1_850 (.ZN (n_0_590), .A (n_0_1_447), .B1 (n_0_1_471), .B2 (n_0_1_792));
AOI222_X1 i_0_1_849 (.ZN (n_0_1_446), .A1 (\A_imm_2s_complement[8] ), .A2 (n_0_1_473)
    , .B1 (slo___n2248), .B2 (slo__n1788), .C1 (\A_imm_2s_complement[7] ), .C2 (drc_ipo_n53));
OAI21_X1 i_0_1_848 (.ZN (n_0_589), .A (n_0_1_446), .B1 (n_0_1_471), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_847 (.ZN (n_0_1_445), .A1 (CLOCK_spw__n7291), .A2 (opt_ipo_n5285)
    , .B1 (slo___n2247), .B2 (\A_imm[6] ), .C1 (drc_ipo_n53), .C2 (opt_ipo_n5205));
OAI21_X1 i_0_1_846 (.ZN (n_0_588), .A (n_0_1_445), .B1 (n_0_1_471), .B2 (sgo__n874));
AOI222_X1 i_0_1_845 (.ZN (n_0_1_444), .A1 (opt_ipo_n5205), .A2 (n_0_1_473), .B1 (slo___n2248)
    , .B2 (slo__n3378), .C1 (drc_ipo_n53), .C2 (\A_imm_2s_complement[5] ));
OAI21_X1 i_0_1_844 (.ZN (n_0_587), .A (n_0_1_444), .B1 (n_0_1_471), .B2 (slo__xsl_n1694));
AOI222_X2 i_0_1_843 (.ZN (n_0_1_443), .A1 (n_0_1_473), .A2 (\A_imm_2s_complement[5] )
    , .B1 (n_0_1_472), .B2 (sgo__n962), .C1 (n_0_1_470), .C2 (\A_imm_2s_complement[4] ));
OAI21_X1 i_0_1_842 (.ZN (n_0_586), .A (n_0_1_443), .B1 (n_0_1_471), .B2 (n_0_1_784));
AOI222_X1 i_0_1_841 (.ZN (n_0_1_442), .A1 (\A_imm_2s_complement[4] ), .A2 (n_0_1_473)
    , .B1 (slo___n2247), .B2 (slo__n1801), .C1 (drc_ipo_n53), .C2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_840 (.ZN (n_0_585), .A (n_0_1_442), .B1 (n_0_1_471), .B2 (sgo__n959));
AOI222_X1 i_0_1_839 (.ZN (n_0_1_441), .A1 (\A_imm_2s_complement[3] ), .A2 (n_0_1_473)
    , .B1 (slo___n2247), .B2 (sgo__n1053), .C1 (drc_ipo_n53), .C2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_838 (.ZN (n_0_584), .A (n_0_1_441), .B1 (n_0_1_471), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_837 (.ZN (n_0_1_440), .A1 (\A_imm_2s_complement[2] ), .A2 (opt_ipo_n5285)
    , .B1 (slo___n2247), .B2 (opt_ipo_n5459), .C1 (drc_ipo_n53), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_836 (.ZN (n_0_583), .A (n_0_1_440), .B1 (n_0_1_471), .B2 (sgo__n1043));
NAND2_X1 i_0_1_835 (.ZN (n_0_1_439), .A1 (\A_imm_2s_complement[1] ), .A2 (opt_ipo_n5285));
OAI21_X1 i_0_1_834 (.ZN (n_0_1_438), .A (sgo__n759), .B1 (slo___n2247), .B2 (drc_ipo_n53));
OAI211_X1 i_0_1_833 (.ZN (n_0_582), .A (n_0_1_439), .B (n_0_1_438), .C1 (n_0_1_776), .C2 (n_0_1_471));
AND2_X1 i_0_1_832 (.ZN (n_0_581), .A1 (n_0_1_474), .A2 (sgo__n759));
MUX2_X2 i_0_1_831 (.Z (n_0_1_437), .A (n_0_170), .B (n_0_46), .S (drc_ipo_n58));
NAND2_X2 i_0_1_830 (.ZN (n_0_1_436), .A1 (slo__xsl_n1963), .A2 (n_0_1_437));
MUX2_X2 i_0_1_829 (.Z (n_0_1_435), .A (n_0_169), .B (n_0_47), .S (drc_ipo_n58));
INV_X4 i_0_1_828 (.ZN (n_0_1_434), .A (slo__n3134));
NAND3_X1 i_0_1_827 (.ZN (n_0_1_433), .A1 (n_0_1_436), .A2 (n_0_1_435), .A3 (sgo__n731));
OAI21_X1 i_0_1_826 (.ZN (n_0_1_432), .A (\A_imm[31] ), .B1 (slo__xsl_n1963), .B2 (n_0_1_437));
OAI21_X1 i_0_1_825 (.ZN (n_0_580), .A (n_0_1_433), .B1 (n_0_1_432), .B2 (n_0_1_435));
XNOR2_X2 i_0_1_824 (.ZN (n_0_1_431), .A (n_0_1_477), .B (n_0_1_437));
AND2_X2 i_0_1_823 (.ZN (n_0_1_430), .A1 (n_0_1_435), .A2 (n_0_1_431));
MUX2_X2 slo__c3023 (.Z (slo__n2712), .A (n_0_161), .B (n_0_55), .S (drc_ipo_n58));
NAND2_X4 i_0_1_821 (.ZN (n_0_1_428), .A1 (n_0_1_431), .A2 (n_0_1_434));
NOR3_X2 i_0_1_820 (.ZN (n_0_1_427), .A1 (n_0_1_434), .A2 (n_0_1_437), .A3 (slo__xsl_n1963));
AOI222_X1 i_0_1_819 (.ZN (n_0_1_426), .A1 (sgo__n731), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (\A_imm[30] ), .C1 (opt_ipo_n5419), .C2 (opt_ipo_n5358));
OAI21_X1 i_0_1_818 (.ZN (n_0_579), .A (n_0_1_426), .B1 (n_0_1_428), .B2 (n_0_1_836));
AOI222_X1 i_0_1_817 (.ZN (n_0_1_425), .A1 (\A_imm_2s_complement[30] ), .A2 (sgo__n779)
    , .B1 (opt_ipo_n5686), .B2 (\A_imm[29] ), .C1 (opt_ipo_n5419), .C2 (\A_imm_2s_complement[29] ));
OAI21_X1 i_0_1_816 (.ZN (n_0_578), .A (n_0_1_425), .B1 (n_0_1_428), .B2 (sgo__n734));
AOI222_X1 i_0_1_815 (.ZN (n_0_1_424), .A1 (sgo__n1241), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (\A_imm[28] ), .C1 (opt_ipo_n5419), .C2 (sgo__n678));
OAI21_X1 i_0_1_814 (.ZN (n_0_577), .A (n_0_1_424), .B1 (n_0_1_428), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_813 (.ZN (n_0_1_423), .A1 (sgo__n678), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (\A_imm[27] ), .C1 (opt_ipo_n5419), .C2 (sgo__n877));
OAI21_X1 i_0_1_812 (.ZN (n_0_576), .A (n_0_1_423), .B1 (n_0_1_428), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_811 (.ZN (n_0_1_422), .A1 (\A_imm_2s_complement[27] ), .A2 (sgo__n779)
    , .B1 (opt_ipo_n5686), .B2 (slo__n1897), .C1 (opt_ipo_n5419), .C2 (\A_imm_2s_complement[26] ));
OAI21_X1 i_0_1_810 (.ZN (n_0_575), .A (n_0_1_422), .B1 (n_0_1_428), .B2 (slo__n2762));
AOI222_X1 i_0_1_809 (.ZN (n_0_1_421), .A1 (sgo__n943), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (opt_ipo_n5362), .C1 (opt_ipo_n5419), .C2 (\A_imm_2s_complement[25] ));
OAI21_X1 i_0_1_808 (.ZN (n_0_574), .A (n_0_1_421), .B1 (n_0_1_428), .B2 (slo__xsl_n1889));
AOI222_X1 i_0_1_807 (.ZN (n_0_1_420), .A1 (\A_imm_2s_complement[25] ), .A2 (sgo__n779)
    , .B1 (opt_ipo_n5686), .B2 (slo__n2216), .C1 (\A_imm_2s_complement[24] ), .C2 (opt_ipo_n5419));
OAI21_X1 i_0_1_806 (.ZN (n_0_573), .A (n_0_1_420), .B1 (n_0_1_428), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_805 (.ZN (n_0_1_419), .A1 (slo__n1550), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (slo__n3760), .C1 (opt_ipo_n5419), .C2 (sgo__n839));
OAI21_X1 i_0_1_804 (.ZN (n_0_572), .A (n_0_1_419), .B1 (n_0_1_428), .B2 (sgo__n1238));
AOI222_X1 i_0_1_803 (.ZN (n_0_1_418), .A1 (sgo__n839), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (slo__n1649), .C1 (opt_ipo_n5419), .C2 (sgo__n836));
OAI21_X1 i_0_1_802 (.ZN (n_0_571), .A (n_0_1_418), .B1 (n_0_1_428), .B2 (slo__n1812));
AOI222_X1 i_0_1_801 (.ZN (n_0_1_417), .A1 (sgo__n836), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (opt_ipo_n5135), .C1 (opt_ipo_n5419), .C2 (sgo__n1009));
OAI21_X1 i_0_1_800 (.ZN (n_0_570), .A (n_0_1_417), .B1 (n_0_1_428), .B2 (slo__xsl_n1641));
AOI222_X1 i_0_1_799 (.ZN (n_0_1_416), .A1 (\A_imm_2s_complement[21] ), .A2 (sgo__n779)
    , .B1 (opt_ipo_n5686), .B2 (opt_ipo_n5196), .C1 (opt_ipo_n5419), .C2 (opt_ipo_n5785));
OAI21_X1 i_0_1_798 (.ZN (n_0_569), .A (n_0_1_416), .B1 (n_0_1_428), .B2 (opt_ipo_n5145));
AOI222_X1 i_0_1_797 (.ZN (n_0_1_415), .A1 (opt_ipo_n5339), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (opt_ipo_n5303), .C1 (opt_ipo_n5419), .C2 (opt_ipo_n5373));
OAI21_X1 i_0_1_796 (.ZN (n_0_568), .A (n_0_1_415), .B1 (n_0_1_428), .B2 (opt_ipo_n5195));
AOI222_X1 i_0_1_795 (.ZN (n_0_1_414), .A1 (opt_ipo_n5373), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (slo__n2915), .C1 (\A_imm_2s_complement[18] ), .C2 (opt_ipo_n5419));
OAI21_X1 i_0_1_794 (.ZN (n_0_567), .A (n_0_1_414), .B1 (n_0_1_428), .B2 (opt_ipo_n5307));
AOI222_X1 i_0_1_793 (.ZN (n_0_1_413), .A1 (\A_imm_2s_complement[18] ), .A2 (sgo__n779)
    , .B1 (opt_ipo_n5686), .B2 (slo__n3402), .C1 (opt_ipo_n5419), .C2 (opt_ipo_n5411));
OAI21_X1 i_0_1_792 (.ZN (n_0_566), .A (n_0_1_413), .B1 (n_0_1_428), .B2 (slo__xsl_n1425));
AOI222_X1 i_0_1_791 (.ZN (n_0_1_412), .A1 (opt_ipo_n5411), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (slo__n3547), .C1 (opt_ipo_n5419), .C2 (\A_imm_2s_complement[16] ));
OAI21_X1 i_0_1_790 (.ZN (n_0_565), .A (n_0_1_412), .B1 (n_0_1_428), .B2 (slo__xsl_n1366));
AOI222_X1 i_0_1_789 (.ZN (n_0_1_411), .A1 (opt_ipo_n5162), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (opt_ipo_n5415), .C1 (opt_ipo_n5419), .C2 (opt_ipo_n5653));
OAI21_X1 i_0_1_788 (.ZN (n_0_564), .A (n_0_1_411), .B1 (n_0_1_428), .B2 (slo__n1493));
AOI222_X1 i_0_1_787 (.ZN (n_0_1_410), .A1 (sgo__n895), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (\A_imm[14] ), .C1 (opt_ipo_n5419), .C2 (opt_ipo_n5672));
OAI21_X1 i_0_1_786 (.ZN (n_0_563), .A (n_0_1_410), .B1 (n_0_1_428), .B2 (slo__n1828));
AOI222_X2 i_0_1_785 (.ZN (n_0_1_409), .A1 (\A_imm_2s_complement[14] ), .A2 (n_0_1_430)
    , .B1 (opt_ipo_n5686), .B2 (\A_imm[13] ), .C1 (\A_imm_2s_complement[13] ), .C2 (drc_ipo_n54));
OAI21_X1 i_0_1_784 (.ZN (n_0_562), .A (n_0_1_409), .B1 (n_0_1_428), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_783 (.ZN (n_0_1_408), .A1 (opt_ipo_n5710), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (slo__n3230), .C1 (opt_ipo_n5419), .C2 (\A_imm_2s_complement[12] ));
OAI21_X1 i_0_1_782 (.ZN (n_0_561), .A (n_0_1_408), .B1 (n_0_1_428), .B2 (slo__n1559));
AOI222_X2 i_0_1_781 (.ZN (n_0_1_407), .A1 (slo__n1702), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (opt_ipo_n5297), .C1 (opt_ipo_n5419), .C2 (slo__n3026));
OAI21_X1 i_0_1_780 (.ZN (n_0_560), .A (n_0_1_407), .B1 (n_0_1_428), .B2 (slo__n1402));
AOI222_X2 i_0_1_779 (.ZN (n_0_1_406), .A1 (\A_imm_2s_complement[11] ), .A2 (n_0_1_430)
    , .B1 (opt_ipo_n5686), .B2 (opt_ipo_n5164), .C1 (opt_ipo_n5466), .C2 (opt_ipo_n5419));
OAI21_X1 i_0_1_778 (.ZN (n_0_559), .A (n_0_1_406), .B1 (n_0_1_428), .B2 (slo___n3458));
AOI222_X1 i_0_1_777 (.ZN (n_0_1_405), .A1 (opt_ipo_n5466), .A2 (n_0_1_430), .B1 (opt_ipo_n5686)
    , .B2 (\A_imm[9] ), .C1 (opt_ipo_n5419), .C2 (opt_ipo_n5198));
OAI21_X1 i_0_1_776 (.ZN (n_0_558), .A (n_0_1_405), .B1 (n_0_1_428), .B2 (opt_ipo_n5165));
AOI222_X1 i_0_1_775 (.ZN (n_0_1_404), .A1 (opt_ipo_n5197), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (slo__n3281), .C1 (opt_ipo_n5419), .C2 (\A_imm_2s_complement[8] ));
OAI21_X1 i_0_1_774 (.ZN (n_0_557), .A (n_0_1_404), .B1 (n_0_1_428), .B2 (n_0_1_792));
AOI222_X1 i_0_1_773 (.ZN (n_0_1_403), .A1 (slo__n2969), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (slo__n1788), .C1 (opt_ipo_n5419), .C2 (\A_imm_2s_complement[7] ));
OAI21_X1 i_0_1_772 (.ZN (n_0_556), .A (n_0_1_403), .B1 (n_0_1_428), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_771 (.ZN (n_0_1_402), .A1 (\A_imm_2s_complement[7] ), .A2 (n_0_1_430)
    , .B1 (opt_ipo_n5686), .B2 (spw__n7740), .C1 (opt_ipo_n5419), .C2 (opt_ipo_n5205));
OAI21_X1 i_0_1_770 (.ZN (n_0_555), .A (n_0_1_402), .B1 (n_0_1_428), .B2 (sgo__n874));
BUF_X1 spw__L1_c8575 (.Z (spw__n7776), .A (n_0_1_599));
OAI21_X1 i_0_1_768 (.ZN (n_0_554), .A (n_0_1_401), .B1 (n_0_1_428), .B2 (slo__xsl_n1694));
AOI222_X1 i_0_1_767 (.ZN (n_0_1_400), .A1 (slo__n3910), .A2 (sgo__n779), .B1 (opt_ipo_n5686)
    , .B2 (sgo__n962), .C1 (opt_ipo_n5419), .C2 (slo__n2805));
OAI21_X1 i_0_1_766 (.ZN (n_0_553), .A (n_0_1_400), .B1 (n_0_1_428), .B2 (n_0_1_784));
AOI222_X1 i_0_1_765 (.ZN (n_0_1_399), .A1 (slo__n2805), .A2 (n_0_1_430), .B1 (n_0_1_429)
    , .B2 (slo__n1801), .C1 (drc_ipo_n54), .C2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_764 (.ZN (n_0_552), .A (n_0_1_399), .B1 (n_0_1_428), .B2 (sgo__n959));
BUF_X4 sgo__c822 (.Z (sgo__n844), .A (\A_imm_2s_complement[30] ));
OAI21_X1 i_0_1_762 (.ZN (n_0_551), .A (sgo__sro_n769), .B1 (n_0_1_428), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_761 (.ZN (n_0_1_397), .A1 (\A_imm_2s_complement[2] ), .A2 (n_0_1_430)
    , .B1 (opt_ipo_n5686), .B2 (opt_ipo_n5459), .C1 (opt_ipo_n5419), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_760 (.ZN (n_0_550), .A (n_0_1_397), .B1 (n_0_1_428), .B2 (sgo__n1043));
NAND2_X1 i_0_1_759 (.ZN (n_0_1_396), .A1 (\A_imm_2s_complement[1] ), .A2 (n_0_1_430));
OAI21_X1 i_0_1_758 (.ZN (n_0_1_395), .A (sgo__n759), .B1 (opt_ipo_n5686), .B2 (opt_ipo_n5419));
OAI211_X1 i_0_1_757 (.ZN (n_0_549), .A (n_0_1_396), .B (n_0_1_395), .C1 (n_0_1_776), .C2 (n_0_1_428));
AND2_X1 i_0_1_756 (.ZN (n_0_548), .A1 (n_0_1_431), .A2 (sgo__n759));
INV_X1 CLOCK_slo__sro_c7468 (.ZN (CLOCK_slo__sro_n6743), .A (n_0_1_686));
INV_X2 i_0_1_754 (.ZN (n_0_1_393), .A (n_0_1_394));
MUX2_X2 i_0_1_753 (.Z (n_0_1_392), .A (n_0_168), .B (n_0_48), .S (drc_ipo_n58));
OAI21_X1 i_0_1_752 (.ZN (n_0_1_391), .A (\A_imm[31] ), .B1 (n_0_1_435), .B2 (opt_ipo_n5720));
NAND2_X1 i_0_1_751 (.ZN (n_0_1_390), .A1 (slo__n3134), .A2 (n_0_1_392));
NAND3_X1 i_0_1_750 (.ZN (n_0_1_389), .A1 (n_0_1_390), .A2 (sgo__n731), .A3 (n_0_1_394));
OAI21_X2 i_0_1_749 (.ZN (n_0_547), .A (n_0_1_389), .B1 (n_0_1_391), .B2 (n_0_1_394));
XNOR2_X2 i_0_1_748 (.ZN (n_0_1_388), .A (n_0_1_434), .B (n_0_1_392));
AND2_X4 i_0_1_747 (.ZN (n_0_1_387), .A1 (n_0_1_394), .A2 (n_0_1_388));
NOR2_X1 i_0_1_746 (.ZN (n_0_1_386), .A1 (n_0_1_394), .A2 (n_0_1_390));
NAND2_X1 i_0_1_745 (.ZN (n_0_1_385), .A1 (n_0_1_388), .A2 (n_0_1_393));
NOR3_X4 i_0_1_744 (.ZN (n_0_1_384), .A1 (n_0_1_393), .A2 (opt_ipo_n5720), .A3 (n_0_1_435));
AOI222_X1 i_0_1_743 (.ZN (n_0_1_383), .A1 (sgo__n731), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (\A_imm[30] ), .C1 (opt_ipo_n5719), .C2 (opt_ipo_n5358));
OAI21_X1 i_0_1_742 (.ZN (n_0_546), .A (n_0_1_383), .B1 (CLOCK_spw__n7321), .B2 (n_0_1_836));
AOI222_X1 i_0_1_741 (.ZN (n_0_1_382), .A1 (opt_ipo_n5358), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (\A_imm[29] ), .C1 (opt_ipo_n5719), .C2 (sgo__n1241));
OAI21_X1 i_0_1_740 (.ZN (n_0_545), .A (n_0_1_382), .B1 (CLOCK_spw__n7321), .B2 (sgo__n734));
AOI222_X1 i_0_1_739 (.ZN (n_0_1_381), .A1 (sgo__n1241), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (\A_imm[28] ), .C1 (opt_ipo_n5719), .C2 (sgo__n678));
OAI21_X1 i_0_1_738 (.ZN (n_0_544), .A (n_0_1_381), .B1 (CLOCK_spw__n7321), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_737 (.ZN (n_0_1_380), .A1 (sgo__n678), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (\A_imm[27] ), .C1 (opt_ipo_n5719), .C2 (\A_imm_2s_complement[27] ));
OAI21_X1 i_0_1_736 (.ZN (n_0_543), .A (n_0_1_380), .B1 (CLOCK_spw__n7321), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_735 (.ZN (n_0_1_379), .A1 (sgo__n877), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (slo__n1897), .C1 (opt_ipo_n5719), .C2 (sgo__n943));
OAI21_X1 i_0_1_734 (.ZN (n_0_542), .A (n_0_1_379), .B1 (CLOCK_spw__n7321), .B2 (slo__n2762));
AOI222_X1 i_0_1_733 (.ZN (n_0_1_378), .A1 (sgo__n943), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (opt_ipo_n5362), .C1 (sgo__n1339), .C2 (opt_ipo_n5719));
OAI21_X1 i_0_1_732 (.ZN (n_0_541), .A (n_0_1_378), .B1 (CLOCK_spw__n7321), .B2 (slo__xsl_n1889));
AOI222_X1 i_0_1_731 (.ZN (n_0_1_377), .A1 (sgo__n1339), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (slo__n2216), .C1 (slo__n1550), .C2 (opt_ipo_n5719));
OAI21_X1 i_0_1_730 (.ZN (n_0_540), .A (n_0_1_377), .B1 (CLOCK_spw__n7321), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_729 (.ZN (n_0_1_376), .A1 (slo__n1550), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (slo__n3760), .C1 (opt_ipo_n5719), .C2 (sgo__n839));
OAI21_X1 i_0_1_728 (.ZN (n_0_539), .A (n_0_1_376), .B1 (CLOCK_spw__n7321), .B2 (sgo__n1238));
AOI222_X1 i_0_1_727 (.ZN (n_0_1_375), .A1 (sgo__n839), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (slo__n1649), .C1 (opt_ipo_n5719), .C2 (\A_imm_2s_complement[22] ));
OAI21_X1 i_0_1_726 (.ZN (n_0_538), .A (n_0_1_375), .B1 (CLOCK_spw__n7321), .B2 (slo__n1812));
AOI222_X1 i_0_1_725 (.ZN (n_0_1_374), .A1 (sgo__n836), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (opt_ipo_n5135), .C1 (opt_ipo_n5719), .C2 (sgo__n1009));
OAI21_X1 i_0_1_724 (.ZN (n_0_537), .A (n_0_1_374), .B1 (CLOCK_spw__n7321), .B2 (slo__xsl_n1641));
AOI222_X1 i_0_1_723 (.ZN (n_0_1_373), .A1 (sgo__n1009), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (opt_ipo_n5196), .C1 (opt_ipo_n5719), .C2 (opt_ipo_n5339));
OAI21_X1 i_0_1_722 (.ZN (n_0_536), .A (n_0_1_373), .B1 (CLOCK_spw__n7321), .B2 (opt_ipo_n5145));
AOI222_X1 i_0_1_721 (.ZN (n_0_1_372), .A1 (opt_ipo_n5339), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (opt_ipo_n5303), .C1 (opt_ipo_n5373), .C2 (opt_ipo_n5719));
OAI21_X1 i_0_1_720 (.ZN (n_0_535), .A (n_0_1_372), .B1 (CLOCK_spw__n7321), .B2 (opt_ipo_n5195));
AOI222_X1 i_0_1_719 (.ZN (n_0_1_371), .A1 (opt_ipo_n5373), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (slo__n2915), .C1 (opt_ipo_n5719), .C2 (\A_imm_2s_complement[18] ));
OAI21_X1 i_0_1_718 (.ZN (n_0_534), .A (n_0_1_371), .B1 (CLOCK_spw__n7321), .B2 (opt_ipo_n5307));
AOI222_X1 i_0_1_717 (.ZN (n_0_1_370), .A1 (\A_imm_2s_complement[18] ), .A2 (slo___n3116)
    , .B1 (slo___n3416), .B2 (slo__n3402), .C1 (opt_ipo_n5719), .C2 (opt_ipo_n5411));
OAI21_X1 i_0_1_716 (.ZN (n_0_533), .A (n_0_1_370), .B1 (CLOCK_spw__n7321), .B2 (slo__xsl_n1425));
AOI222_X1 i_0_1_715 (.ZN (n_0_1_369), .A1 (opt_ipo_n5411), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (slo__n3547), .C1 (opt_ipo_n5719), .C2 (\A_imm_2s_complement[16] ));
OAI21_X1 i_0_1_714 (.ZN (n_0_532), .A (n_0_1_369), .B1 (CLOCK_spw__n7321), .B2 (slo__xsl_n1366));
AOI222_X1 i_0_1_713 (.ZN (n_0_1_368), .A1 (sgo__n1056), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (opt_ipo_n5415), .C1 (opt_ipo_n5719), .C2 (sgo__n895));
OAI21_X1 i_0_1_712 (.ZN (n_0_531), .A (n_0_1_368), .B1 (CLOCK_spw__n7321), .B2 (slo__n1493));
AOI222_X1 i_0_1_711 (.ZN (n_0_1_367), .A1 (sgo__n895), .A2 (slo___n3116), .B1 (slo___n3416)
    , .B2 (\A_imm[14] ), .C1 (n_0_1_384), .C2 (\A_imm_2s_complement[14] ));
OAI21_X1 i_0_1_710 (.ZN (n_0_530), .A (n_0_1_367), .B1 (CLOCK_spw__n7320), .B2 (slo__n1828));
AOI222_X1 i_0_1_709 (.ZN (n_0_1_366), .A1 (slo__n2107), .A2 (slo___n3116), .B1 (opt_ipo_n5159)
    , .B2 (\A_imm[13] ), .C1 (opt_ipo_n5719), .C2 (opt_ipo_n5710));
OAI21_X1 i_0_1_708 (.ZN (n_0_529), .A (n_0_1_366), .B1 (CLOCK_spw__n7320), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_707 (.ZN (n_0_1_365), .A1 (opt_ipo_n5710), .A2 (slo___n3116), .B1 (opt_ipo_n5159)
    , .B2 (slo__n3230), .C1 (opt_ipo_n5719), .C2 (\A_imm_2s_complement[12] ));
OAI21_X1 i_0_1_706 (.ZN (n_0_528), .A (n_0_1_365), .B1 (CLOCK_spw__n7320), .B2 (slo__n1559));
AOI222_X1 i_0_1_705 (.ZN (n_0_1_364), .A1 (\A_imm_2s_complement[12] ), .A2 (slo___n3116)
    , .B1 (opt_ipo_n5159), .B2 (opt_ipo_n5297), .C1 (n_0_1_384), .C2 (\A_imm_2s_complement[11] ));
OAI21_X1 i_0_1_704 (.ZN (n_0_527), .A (n_0_1_364), .B1 (CLOCK_spw__n7320), .B2 (slo__n1402));
AOI222_X1 i_0_1_703 (.ZN (n_0_1_363), .A1 (slo__n3026), .A2 (slo___n3116), .B1 (opt_ipo_n5159)
    , .B2 (opt_ipo_n5164), .C1 (n_0_1_384), .C2 (opt_ipo_n5466));
OAI21_X1 i_0_1_702 (.ZN (n_0_526), .A (n_0_1_363), .B1 (CLOCK_spw__n7320), .B2 (slo___n3458));
AOI222_X1 i_0_1_701 (.ZN (n_0_1_362), .A1 (opt_ipo_n5465), .A2 (n_0_1_387), .B1 (opt_ipo_n5159)
    , .B2 (\A_imm[9] ), .C1 (opt_ipo_n5719), .C2 (opt_ipo_n5197));
OAI21_X1 i_0_1_700 (.ZN (n_0_525), .A (n_0_1_362), .B1 (CLOCK_spw__n7322), .B2 (opt_ipo_n5165));
AOI222_X1 i_0_1_699 (.ZN (n_0_1_361), .A1 (opt_ipo_n5197), .A2 (n_0_1_387), .B1 (opt_ipo_n5159)
    , .B2 (slo__n3281), .C1 (n_0_1_384), .C2 (\A_imm_2s_complement[8] ));
OAI21_X1 i_0_1_698 (.ZN (n_0_524), .A (n_0_1_361), .B1 (CLOCK_spw__n7320), .B2 (n_0_1_792));
AOI222_X1 i_0_1_697 (.ZN (n_0_1_360), .A1 (slo__n2969), .A2 (n_0_1_387), .B1 (opt_ipo_n5159)
    , .B2 (slo__n1788), .C1 (n_0_1_384), .C2 (\A_imm_2s_complement[7] ));
OAI21_X1 i_0_1_696 (.ZN (n_0_523), .A (n_0_1_360), .B1 (CLOCK_spw__n7320), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_695 (.ZN (n_0_1_359), .A1 (CLOCK_spw__n7292), .A2 (n_0_1_387), .B1 (opt_ipo_n5159)
    , .B2 (spw__n7740), .C1 (opt_ipo_n5719), .C2 (opt_ipo_n5205));
OAI21_X1 i_0_1_694 (.ZN (n_0_522), .A (n_0_1_359), .B1 (CLOCK_spw__n7322), .B2 (sgo__n874));
AOI222_X1 i_0_1_693 (.ZN (n_0_1_358), .A1 (opt_ipo_n5204), .A2 (n_0_1_387), .B1 (opt_ipo_n5159)
    , .B2 (slo__n3378), .C1 (opt_ipo_n5719), .C2 (slo__n3910));
OAI21_X1 i_0_1_692 (.ZN (n_0_521), .A (n_0_1_358), .B1 (n_0_1_385), .B2 (slo__xsl_n1694));
AOI222_X1 i_0_1_691 (.ZN (n_0_1_357), .A1 (\A_imm_2s_complement[5] ), .A2 (n_0_1_387)
    , .B1 (opt_ipo_n5159), .B2 (sgo__n962), .C1 (opt_ipo_n5719), .C2 (\A_imm_2s_complement[4] ));
OAI21_X1 i_0_1_690 (.ZN (n_0_520), .A (n_0_1_357), .B1 (n_0_1_385), .B2 (n_0_1_784));
AOI222_X1 i_0_1_689 (.ZN (n_0_1_356), .A1 (slo__n2805), .A2 (n_0_1_387), .B1 (opt_ipo_n5159)
    , .B2 (slo__n1801), .C1 (n_0_1_384), .C2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_688 (.ZN (n_0_519), .A (n_0_1_356), .B1 (n_0_1_385), .B2 (sgo__n959));
AOI222_X1 i_0_1_687 (.ZN (n_0_1_355), .A1 (\A_imm_2s_complement[3] ), .A2 (n_0_1_387)
    , .B1 (opt_ipo_n5159), .B2 (sgo__n1053), .C1 (opt_ipo_n5719), .C2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_686 (.ZN (n_0_518), .A (n_0_1_355), .B1 (n_0_1_385), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_685 (.ZN (n_0_1_354), .A1 (\A_imm_2s_complement[2] ), .A2 (n_0_1_387)
    , .B1 (opt_ipo_n5159), .B2 (opt_ipo_n5459), .C1 (n_0_1_384), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_684 (.ZN (n_0_517), .A (n_0_1_354), .B1 (n_0_1_385), .B2 (sgo__n1043));
NAND2_X1 i_0_1_683 (.ZN (n_0_1_353), .A1 (n_0_1_387), .A2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_682 (.ZN (n_0_1_352), .A (sgo__n759), .B1 (opt_ipo_n5159), .B2 (n_0_1_384));
OAI211_X2 i_0_1_681 (.ZN (n_0_516), .A (n_0_1_353), .B (n_0_1_352), .C1 (n_0_1_776), .C2 (n_0_1_385));
AND2_X1 i_0_1_680 (.ZN (n_0_515), .A1 (n_0_1_388), .A2 (sgo__n759));
MUX2_X1 i_0_1_679 (.Z (n_0_1_351), .A (n_0_166), .B (n_0_50), .S (drc_ipo_n58));
OAI21_X1 i_0_1_678 (.ZN (n_0_1_350), .A (\A_imm[31] ), .B1 (n_0_1_394), .B2 (n_0_1_351));
MUX2_X2 i_0_1_677 (.Z (n_0_1_349), .A (n_0_165), .B (n_0_51), .S (drc_ipo_n58));
INV_X2 i_0_1_676 (.ZN (n_0_1_348), .A (slo__n3204));
NAND2_X1 i_0_1_675 (.ZN (n_0_1_347), .A1 (n_0_1_394), .A2 (n_0_1_351));
NAND3_X1 i_0_1_674 (.ZN (n_0_1_346), .A1 (n_0_1_347), .A2 (sgo__n731), .A3 (n_0_1_349));
OAI21_X1 i_0_1_673 (.ZN (n_0_514), .A (n_0_1_346), .B1 (n_0_1_349), .B2 (n_0_1_350));
XNOR2_X2 i_0_1_672 (.ZN (n_0_1_345), .A (n_0_1_351), .B (n_0_1_393));
NAND3_X1 CLOCK_slo__mro_c7544 (.ZN (CLOCK_slo__mro_n6798), .A1 (CLOCK_slo__mro_n6799)
    , .A2 (sgo__sro_n697), .A3 (sgo__sro_n722));
NOR2_X4 i_0_1_670 (.ZN (n_0_1_343), .A1 (n_0_1_349), .A2 (n_0_1_347));
NAND2_X4 i_0_1_669 (.ZN (n_0_1_342), .A1 (n_0_1_345), .A2 (n_0_1_348));
NAND2_X4 CLOCK_slo__mro_c7450 (.ZN (CLOCK_slo__mro_n6730), .A1 (n_0_1_345), .A2 (n_0_1_349));
AOI222_X1 i_0_1_667 (.ZN (n_0_1_340), .A1 (sgo__n731), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (\A_imm[30] ), .C1 (opt_ipo_n5332), .C2 (opt_ipo_n5358));
OAI21_X1 i_0_1_666 (.ZN (n_0_513), .A (n_0_1_340), .B1 (n_0_1_342), .B2 (n_0_1_836));
AOI222_X1 i_0_1_665 (.ZN (n_0_1_339), .A1 (opt_ipo_n5358), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (\A_imm[29] ), .C1 (opt_ipo_n5332), .C2 (sgo__n1241));
OAI21_X1 i_0_1_664 (.ZN (n_0_512), .A (n_0_1_339), .B1 (n_0_1_342), .B2 (sgo__n734));
AOI222_X1 i_0_1_663 (.ZN (n_0_1_338), .A1 (sgo__n1241), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (\A_imm[28] ), .C1 (opt_ipo_n5332), .C2 (sgo__n678));
OAI21_X1 i_0_1_662 (.ZN (n_0_511), .A (n_0_1_338), .B1 (n_0_1_342), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_661 (.ZN (n_0_1_337), .A1 (sgo__n678), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (\A_imm[27] ), .C1 (opt_ipo_n5332), .C2 (sgo__n877));
OAI21_X1 i_0_1_660 (.ZN (n_0_510), .A (n_0_1_337), .B1 (n_0_1_342), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_659 (.ZN (n_0_1_336), .A1 (sgo__n877), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (slo__n1897), .C1 (opt_ipo_n5332), .C2 (sgo__n943));
OAI21_X1 i_0_1_658 (.ZN (n_0_509), .A (n_0_1_336), .B1 (n_0_1_342), .B2 (slo__n2762));
AOI222_X2 i_0_1_657 (.ZN (n_0_1_335), .A1 (sgo__n943), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (opt_ipo_n5362), .C1 (sgo__n1339), .C2 (opt_ipo_n5332));
OAI21_X1 i_0_1_656 (.ZN (n_0_508), .A (n_0_1_335), .B1 (n_0_1_342), .B2 (slo__xsl_n1889));
AOI222_X1 i_0_1_655 (.ZN (n_0_1_334), .A1 (sgo__n1339), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (slo__n2216), .C1 (opt_ipo_n5332), .C2 (slo__n1550));
OAI21_X1 i_0_1_654 (.ZN (n_0_507), .A (n_0_1_334), .B1 (n_0_1_342), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_653 (.ZN (n_0_1_333), .A1 (slo__n1550), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (slo__n3760), .C1 (opt_ipo_n5332), .C2 (sgo__n839));
OAI21_X1 i_0_1_652 (.ZN (n_0_506), .A (n_0_1_333), .B1 (n_0_1_342), .B2 (sgo__n1238));
AOI222_X1 i_0_1_651 (.ZN (n_0_1_332), .A1 (sgo__n839), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (slo__n1649), .C1 (opt_ipo_n5332), .C2 (sgo__n836));
OAI21_X1 i_0_1_650 (.ZN (n_0_505), .A (n_0_1_332), .B1 (n_0_1_342), .B2 (slo__n1812));
AOI222_X1 i_0_1_649 (.ZN (n_0_1_331), .A1 (sgo__n836), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (opt_ipo_n5135), .C1 (opt_ipo_n5332), .C2 (sgo__n1009));
OAI21_X1 i_0_1_648 (.ZN (n_0_504), .A (n_0_1_331), .B1 (n_0_1_342), .B2 (slo__xsl_n1641));
AOI222_X1 i_0_1_647 (.ZN (n_0_1_330), .A1 (\A_imm_2s_complement[21] ), .A2 (n_0_1_344)
    , .B1 (n_0_1_343), .B2 (opt_ipo_n5196), .C1 (opt_ipo_n5339), .C2 (opt_ipo_n5332));
OAI21_X1 i_0_1_646 (.ZN (n_0_503), .A (n_0_1_330), .B1 (n_0_1_342), .B2 (opt_ipo_n5145));
AOI222_X1 i_0_1_645 (.ZN (n_0_1_329), .A1 (opt_ipo_n5339), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (opt_ipo_n5303), .C1 (opt_ipo_n5332), .C2 (opt_ipo_n5373));
OAI21_X1 i_0_1_644 (.ZN (n_0_502), .A (n_0_1_329), .B1 (n_0_1_342), .B2 (opt_ipo_n5195));
AOI222_X1 i_0_1_643 (.ZN (n_0_1_328), .A1 (opt_ipo_n5373), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (slo__n2915), .C1 (opt_ipo_n5332), .C2 (\A_imm_2s_complement[18] ));
OAI21_X1 i_0_1_642 (.ZN (n_0_501), .A (n_0_1_328), .B1 (n_0_1_342), .B2 (opt_ipo_n5307));
AOI222_X1 i_0_1_641 (.ZN (n_0_1_327), .A1 (\A_imm_2s_complement[18] ), .A2 (n_0_1_344)
    , .B1 (n_0_1_343), .B2 (slo__n3402), .C1 (opt_ipo_n5332), .C2 (opt_ipo_n5411));
OAI21_X1 i_0_1_640 (.ZN (n_0_500), .A (n_0_1_327), .B1 (n_0_1_342), .B2 (slo__xsl_n1425));
AOI222_X1 i_0_1_639 (.ZN (n_0_1_326), .A1 (opt_ipo_n5411), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (slo__n3547), .C1 (opt_ipo_n5332), .C2 (\A_imm_2s_complement[16] ));
OAI21_X1 i_0_1_638 (.ZN (n_0_499), .A (n_0_1_326), .B1 (n_0_1_342), .B2 (slo__xsl_n1366));
AOI222_X1 i_0_1_637 (.ZN (n_0_1_325), .A1 (opt_ipo_n5162), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (opt_ipo_n5415), .C1 (sgo__n895), .C2 (opt_ipo_n5332));
OAI21_X1 i_0_1_636 (.ZN (n_0_498), .A (n_0_1_325), .B1 (n_0_1_342), .B2 (slo__n1493));
AOI222_X1 i_0_1_635 (.ZN (n_0_1_324), .A1 (sgo__n895), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (\A_imm[14] ), .C1 (opt_ipo_n5332), .C2 (\A_imm_2s_complement[14] ));
OAI21_X1 i_0_1_634 (.ZN (n_0_497), .A (n_0_1_324), .B1 (n_0_1_342), .B2 (slo__n1828));
AOI222_X1 i_0_1_633 (.ZN (n_0_1_323), .A1 (slo__n2107), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (\A_imm[13] ), .C1 (opt_ipo_n5332), .C2 (opt_ipo_n5710));
OAI21_X1 i_0_1_632 (.ZN (n_0_496), .A (n_0_1_323), .B1 (n_0_1_342), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_631 (.ZN (n_0_1_322), .A1 (opt_ipo_n5710), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (slo__n3230), .C1 (slo__sro_n2149), .C2 (\A_imm_2s_complement[12] ));
OAI21_X1 i_0_1_630 (.ZN (n_0_495), .A (n_0_1_322), .B1 (n_0_1_342), .B2 (slo__n1559));
AOI222_X1 i_0_1_629 (.ZN (n_0_1_321), .A1 (slo__n1702), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (opt_ipo_n5297), .C1 (slo__sro_n2149), .C2 (slo__n3026));
OAI21_X1 i_0_1_628 (.ZN (n_0_494), .A (n_0_1_321), .B1 (n_0_1_342), .B2 (slo__n1402));
AOI222_X1 i_0_1_627 (.ZN (n_0_1_320), .A1 (slo__n3026), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (opt_ipo_n5164), .C1 (opt_ipo_n5332), .C2 (opt_ipo_n5466));
OAI21_X1 i_0_1_626 (.ZN (n_0_493), .A (n_0_1_320), .B1 (n_0_1_342), .B2 (slo___n3458));
AOI222_X1 i_0_1_625 (.ZN (n_0_1_319), .A1 (opt_ipo_n5466), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (\A_imm[9] ), .C1 (slo__sro_n2149), .C2 (opt_ipo_n5198));
OAI21_X1 i_0_1_624 (.ZN (n_0_492), .A (n_0_1_319), .B1 (n_0_1_342), .B2 (opt_ipo_n5165));
AOI222_X1 i_0_1_623 (.ZN (n_0_1_318), .A1 (opt_ipo_n5197), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (slo__n3281), .C1 (slo__sro_n2149), .C2 (\A_imm_2s_complement[8] ));
OAI21_X1 i_0_1_622 (.ZN (n_0_491), .A (n_0_1_318), .B1 (n_0_1_342), .B2 (n_0_1_792));
AOI222_X1 i_0_1_621 (.ZN (n_0_1_317), .A1 (slo__n2969), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (slo__n1788), .C1 (slo__sro_n2149), .C2 (CLOCK_spw__n7292));
OAI21_X1 i_0_1_620 (.ZN (n_0_490), .A (n_0_1_317), .B1 (n_0_1_342), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_619 (.ZN (n_0_1_316), .A1 (\A_imm_2s_complement[7] ), .A2 (n_0_1_344)
    , .B1 (n_0_1_343), .B2 (spw__n7740), .C1 (slo__sro_n2149), .C2 (opt_ipo_n5205));
OAI21_X1 i_0_1_618 (.ZN (n_0_489), .A (n_0_1_316), .B1 (n_0_1_342), .B2 (sgo__n874));
AOI222_X1 i_0_1_617 (.ZN (n_0_1_315), .A1 (opt_ipo_n5204), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (slo__n3378), .C1 (slo__sro_n2149), .C2 (slo__n3910));
OAI21_X1 i_0_1_616 (.ZN (n_0_488), .A (n_0_1_315), .B1 (n_0_1_342), .B2 (slo__xsl_n1694));
AOI222_X1 i_0_1_615 (.ZN (n_0_1_314), .A1 (slo__n3910), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (sgo__n962), .C1 (slo__sro_n2149), .C2 (slo__n2805));
OAI21_X1 i_0_1_614 (.ZN (n_0_487), .A (n_0_1_314), .B1 (n_0_1_342), .B2 (n_0_1_784));
AOI222_X1 i_0_1_613 (.ZN (n_0_1_313), .A1 (slo__n2805), .A2 (n_0_1_344), .B1 (n_0_1_343)
    , .B2 (slo__n1801), .C1 (slo__sro_n2149), .C2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_612 (.ZN (n_0_486), .A (n_0_1_313), .B1 (n_0_1_342), .B2 (sgo__n959));
AOI222_X1 i_0_1_611 (.ZN (n_0_1_312), .A1 (n_0_1_344), .A2 (\A_imm_2s_complement[3] )
    , .B1 (n_0_1_343), .B2 (sgo__n1053), .C1 (slo__sro_n2149), .C2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_610 (.ZN (n_0_485), .A (n_0_1_312), .B1 (n_0_1_342), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_609 (.ZN (n_0_1_311), .A1 (\A_imm_2s_complement[2] ), .A2 (n_0_1_344)
    , .B1 (n_0_1_343), .B2 (opt_ipo_n5459), .C1 (slo__sro_n2149), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_608 (.ZN (n_0_484), .A (n_0_1_311), .B1 (n_0_1_342), .B2 (sgo__n1043));
NAND2_X1 i_0_1_607 (.ZN (n_0_1_310), .A1 (\A_imm_2s_complement[1] ), .A2 (n_0_1_344));
OAI21_X1 i_0_1_606 (.ZN (n_0_1_309), .A (sgo__n759), .B1 (n_0_1_343), .B2 (opt_ipo_n5332));
OAI211_X1 i_0_1_605 (.ZN (n_0_483), .A (n_0_1_310), .B (n_0_1_309), .C1 (n_0_1_776), .C2 (n_0_1_342));
AND2_X1 i_0_1_604 (.ZN (n_0_482), .A1 (n_0_1_345), .A2 (sgo__n759));
MUX2_X2 i_0_1_603 (.Z (n_0_1_308), .A (n_0_164), .B (n_0_52), .S (drc_ipo_n58));
NOR2_X2 slo__sro_c4063 (.ZN (n_0_1_170), .A1 (n_0_1_174), .A2 (n_0_1_178));
MUX2_X1 i_0_1_601 (.Z (n_0_1_306), .A (n_0_163), .B (n_0_53), .S (drc_ipo_n58));
INV_X1 i_0_1_600 (.ZN (n_0_1_305), .A (n_0_1_306));
NAND3_X1 i_0_1_599 (.ZN (n_0_1_304), .A1 (slo__sro_n3685), .A2 (slo__xsl_n4223), .A3 (sgo__n731));
OAI21_X1 i_0_1_598 (.ZN (n_0_1_303), .A (\A_imm[31] ), .B1 (n_0_1_349), .B2 (n_0_1_308));
OAI21_X1 i_0_1_597 (.ZN (n_0_481), .A (n_0_1_304), .B1 (n_0_1_303), .B2 (slo__xsl_n4223));
XNOR2_X2 i_0_1_596 (.ZN (n_0_1_302), .A (n_0_1_348), .B (n_0_1_308));
AND2_X4 i_0_1_595 (.ZN (n_0_1_301), .A1 (slo__xsl_n4223), .A2 (n_0_1_302));
NOR2_X2 i_0_1_594 (.ZN (n_0_1_300), .A1 (slo__sro_n3685), .A2 (slo__xsl_n4223));
NAND2_X4 i_0_1_593 (.ZN (n_0_1_299), .A1 (n_0_1_302), .A2 (n_0_1_305));
NOR3_X2 i_0_1_592 (.ZN (n_0_1_298), .A1 (n_0_1_305), .A2 (n_0_1_308), .A3 (n_0_1_349));
AOI222_X1 i_0_1_591 (.ZN (n_0_1_297), .A1 (sgo__n731), .A2 (slo__n1475), .B1 (opt_ipo_n5224)
    , .B2 (\A_imm[30] ), .C1 (drc_ipo_n48), .C2 (opt_ipo_n5358));
OAI21_X1 i_0_1_590 (.ZN (n_0_480), .A (n_0_1_297), .B1 (n_0_1_299), .B2 (n_0_1_836));
AOI222_X1 i_0_1_589 (.ZN (n_0_1_296), .A1 (opt_ipo_n5358), .A2 (slo__n1475), .B1 (opt_ipo_n5224)
    , .B2 (\A_imm[29] ), .C1 (drc_ipo_n48), .C2 (sgo__n1241));
OAI21_X1 i_0_1_588 (.ZN (n_0_479), .A (n_0_1_296), .B1 (n_0_1_299), .B2 (sgo__n734));
AOI222_X1 i_0_1_587 (.ZN (n_0_1_295), .A1 (sgo__n1241), .A2 (slo__n1475), .B1 (opt_ipo_n5224)
    , .B2 (\A_imm[28] ), .C1 (drc_ipo_n48), .C2 (sgo__n678));
OAI21_X1 i_0_1_586 (.ZN (n_0_478), .A (n_0_1_295), .B1 (n_0_1_299), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_585 (.ZN (n_0_1_294), .A1 (sgo__n678), .A2 (slo__n1475), .B1 (opt_ipo_n5224)
    , .B2 (\A_imm[27] ), .C1 (drc_ipo_n48), .C2 (sgo__n877));
OAI21_X1 i_0_1_584 (.ZN (n_0_477), .A (n_0_1_294), .B1 (n_0_1_299), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_583 (.ZN (n_0_1_293), .A1 (sgo__n877), .A2 (slo__n1475), .B1 (opt_ipo_n5224)
    , .B2 (slo__n1897), .C1 (drc_ipo_n48), .C2 (sgo__n943));
OAI21_X1 i_0_1_582 (.ZN (n_0_476), .A (n_0_1_293), .B1 (n_0_1_299), .B2 (slo__n2762));
AOI222_X1 i_0_1_581 (.ZN (n_0_1_292), .A1 (sgo__n943), .A2 (slo__n1475), .B1 (opt_ipo_n5224)
    , .B2 (opt_ipo_n5362), .C1 (drc_ipo_n48), .C2 (sgo__n1339));
OAI21_X1 i_0_1_580 (.ZN (n_0_475), .A (n_0_1_292), .B1 (n_0_1_299), .B2 (slo__xsl_n1889));
AOI222_X1 i_0_1_579 (.ZN (n_0_1_291), .A1 (sgo__n1339), .A2 (slo__n1475), .B1 (opt_ipo_n5224)
    , .B2 (slo__n2216), .C1 (drc_ipo_n48), .C2 (slo__n1550));
OAI21_X1 i_0_1_578 (.ZN (n_0_474), .A (n_0_1_291), .B1 (n_0_1_299), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_577 (.ZN (n_0_1_290), .A1 (slo__n1550), .A2 (slo__n1475), .B1 (opt_ipo_n5224)
    , .B2 (slo__n3760), .C1 (drc_ipo_n48), .C2 (sgo__n839));
OAI21_X1 i_0_1_576 (.ZN (n_0_473), .A (n_0_1_290), .B1 (n_0_1_299), .B2 (sgo__n1238));
AOI222_X1 i_0_1_575 (.ZN (n_0_1_289), .A1 (sgo__n839), .A2 (slo__n1475), .B1 (opt_ipo_n5224)
    , .B2 (slo__n1649), .C1 (drc_ipo_n48), .C2 (sgo__n836));
OAI21_X1 i_0_1_574 (.ZN (n_0_472), .A (n_0_1_289), .B1 (n_0_1_299), .B2 (slo__n1812));
AOI222_X1 i_0_1_573 (.ZN (n_0_1_288), .A1 (sgo__n836), .A2 (slo__n1475), .B1 (opt_ipo_n5224)
    , .B2 (opt_ipo_n5135), .C1 (drc_ipo_n48), .C2 (sgo__n1009));
OAI21_X1 i_0_1_572 (.ZN (n_0_471), .A (n_0_1_288), .B1 (n_0_1_299), .B2 (slo__xsl_n1641));
AOI222_X2 i_0_1_571 (.ZN (n_0_1_287), .A1 (sgo__n1009), .A2 (slo__n1475), .B1 (opt_ipo_n5224)
    , .B2 (opt_ipo_n5196), .C1 (drc_ipo_n48), .C2 (opt_ipo_n5339));
OAI21_X1 i_0_1_570 (.ZN (n_0_470), .A (n_0_1_287), .B1 (n_0_1_299), .B2 (opt_ipo_n5145));
AOI222_X1 i_0_1_569 (.ZN (n_0_1_286), .A1 (opt_ipo_n5339), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (opt_ipo_n5303), .C1 (\A_imm_2s_complement[19] ), .C2 (drc_ipo_n48));
OAI21_X1 i_0_1_568 (.ZN (n_0_469), .A (n_0_1_286), .B1 (n_0_1_299), .B2 (opt_ipo_n5195));
AOI222_X1 i_0_1_567 (.ZN (n_0_1_285), .A1 (opt_ipo_n5373), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (slo__n2915), .C1 (drc_ipo_n48), .C2 (\A_imm_2s_complement[18] ));
OAI21_X1 i_0_1_566 (.ZN (n_0_468), .A (n_0_1_285), .B1 (n_0_1_299), .B2 (opt_ipo_n5307));
AOI222_X1 i_0_1_565 (.ZN (n_0_1_284), .A1 (\A_imm_2s_complement[18] ), .A2 (slo__n1475)
    , .B1 (opt_ipo_n5224), .B2 (slo__n3402), .C1 (drc_ipo_n48), .C2 (opt_ipo_n5411));
OAI21_X1 i_0_1_564 (.ZN (n_0_467), .A (n_0_1_284), .B1 (n_0_1_299), .B2 (slo__xsl_n1425));
AOI222_X1 i_0_1_563 (.ZN (n_0_1_283), .A1 (opt_ipo_n5411), .A2 (slo__n1475), .B1 (opt_ipo_n5224)
    , .B2 (slo__n3547), .C1 (drc_ipo_n48), .C2 (sgo__n1056));
OAI21_X1 i_0_1_562 (.ZN (n_0_466), .A (n_0_1_283), .B1 (n_0_1_299), .B2 (slo__xsl_n1366));
AOI222_X1 i_0_1_561 (.ZN (n_0_1_282), .A1 (sgo__n1056), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (opt_ipo_n5415), .C1 (drc_ipo_n48), .C2 (sgo__n895));
OAI21_X1 i_0_1_560 (.ZN (n_0_465), .A (n_0_1_282), .B1 (n_0_1_299), .B2 (slo__n1493));
AOI222_X1 i_0_1_559 (.ZN (n_0_1_281), .A1 (sgo__n895), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (\A_imm[14] ), .C1 (drc_ipo_n48), .C2 (\A_imm_2s_complement[14] ));
OAI21_X1 i_0_1_558 (.ZN (n_0_464), .A (n_0_1_281), .B1 (n_0_1_299), .B2 (slo__n1828));
AOI222_X1 i_0_1_557 (.ZN (n_0_1_280), .A1 (slo__n2107), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (\A_imm[13] ), .C1 (opt_ipo_n5710), .C2 (drc_ipo_n48));
OAI21_X1 i_0_1_556 (.ZN (n_0_463), .A (n_0_1_280), .B1 (n_0_1_299), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_555 (.ZN (n_0_1_279), .A1 (opt_ipo_n5710), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (slo__n3230), .C1 (drc_ipo_n48), .C2 (\A_imm_2s_complement[12] ));
OAI21_X1 i_0_1_554 (.ZN (n_0_462), .A (n_0_1_279), .B1 (n_0_1_299), .B2 (slo__n1559));
AOI222_X1 i_0_1_553 (.ZN (n_0_1_278), .A1 (slo__n1702), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (opt_ipo_n5297), .C1 (drc_ipo_n48), .C2 (slo__n3026));
OAI21_X1 i_0_1_552 (.ZN (n_0_461), .A (n_0_1_278), .B1 (n_0_1_299), .B2 (slo__n1402));
AOI222_X1 i_0_1_551 (.ZN (n_0_1_277), .A1 (slo__n3026), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (opt_ipo_n5164), .C1 (drc_ipo_n48), .C2 (opt_ipo_n5466));
OAI21_X1 i_0_1_550 (.ZN (n_0_460), .A (n_0_1_277), .B1 (n_0_1_299), .B2 (slo___n3458));
AOI222_X1 i_0_1_549 (.ZN (n_0_1_276), .A1 (opt_ipo_n5465), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (\A_imm[9] ), .C1 (drc_ipo_n48), .C2 (opt_ipo_n5197));
OAI21_X1 i_0_1_548 (.ZN (n_0_459), .A (n_0_1_276), .B1 (n_0_1_299), .B2 (opt_ipo_n5165));
AOI222_X1 i_0_1_547 (.ZN (n_0_1_275), .A1 (opt_ipo_n5197), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (slo__n3281), .C1 (drc_ipo_n48), .C2 (slo__n2969));
OAI21_X1 i_0_1_546 (.ZN (n_0_458), .A (n_0_1_275), .B1 (n_0_1_299), .B2 (n_0_1_792));
AOI222_X1 i_0_1_545 (.ZN (n_0_1_274), .A1 (slo__n2969), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (slo__n1788), .C1 (drc_ipo_n48), .C2 (\A_imm_2s_complement[7] ));
OAI21_X1 i_0_1_544 (.ZN (n_0_457), .A (n_0_1_274), .B1 (n_0_1_299), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_543 (.ZN (n_0_1_273), .A1 (CLOCK_spw__n7292), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (spw__n7739), .C1 (drc_ipo_n48), .C2 (opt_ipo_n5205));
OAI21_X1 i_0_1_542 (.ZN (n_0_456), .A (n_0_1_273), .B1 (n_0_1_299), .B2 (sgo__n874));
AOI222_X1 i_0_1_541 (.ZN (n_0_1_272), .A1 (opt_ipo_n5204), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (slo__n3378), .C1 (drc_ipo_n48), .C2 (slo__n3910));
OAI21_X1 i_0_1_540 (.ZN (n_0_455), .A (n_0_1_272), .B1 (n_0_1_299), .B2 (slo__xsl_n1694));
AOI222_X2 i_0_1_539 (.ZN (n_0_1_271), .A1 (n_0_1_301), .A2 (\A_imm_2s_complement[5] )
    , .B1 (opt_ipo_n5224), .B2 (sgo__n962), .C1 (drc_ipo_n48), .C2 (\A_imm_2s_complement[4] ));
OAI21_X1 i_0_1_538 (.ZN (n_0_454), .A (n_0_1_271), .B1 (n_0_1_299), .B2 (n_0_1_784));
AOI222_X1 i_0_1_537 (.ZN (n_0_1_270), .A1 (slo__n2805), .A2 (n_0_1_301), .B1 (opt_ipo_n5224)
    , .B2 (slo__n1801), .C1 (drc_ipo_n48), .C2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_536 (.ZN (n_0_453), .A (n_0_1_270), .B1 (n_0_1_299), .B2 (sgo__n959));
AOI222_X1 i_0_1_535 (.ZN (n_0_1_269), .A1 (\A_imm_2s_complement[3] ), .A2 (n_0_1_301)
    , .B1 (opt_ipo_n5224), .B2 (sgo__n1053), .C1 (drc_ipo_n48), .C2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_534 (.ZN (n_0_452), .A (n_0_1_269), .B1 (n_0_1_299), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_533 (.ZN (n_0_1_268), .A1 (\A_imm_2s_complement[2] ), .A2 (n_0_1_301)
    , .B1 (opt_ipo_n5224), .B2 (opt_ipo_n5459), .C1 (drc_ipo_n48), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_532 (.ZN (n_0_451), .A (n_0_1_268), .B1 (n_0_1_299), .B2 (sgo__n1043));
NAND2_X1 i_0_1_531 (.ZN (n_0_1_267), .A1 (\A_imm_2s_complement[1] ), .A2 (n_0_1_301));
INV_X1 slo__c4036 (.ZN (slo__n3696), .A (n_0_1_914));
OAI211_X1 i_0_1_529 (.ZN (n_0_450), .A (n_0_1_267), .B (slo__sro_n3675), .C1 (n_0_1_299), .C2 (n_0_1_776));
AND2_X1 i_0_1_528 (.ZN (n_0_449), .A1 (n_0_1_302), .A2 (sgo__n759));
MUX2_X1 i_0_1_527 (.Z (n_0_1_265), .A (n_0_162), .B (n_0_54), .S (drc_ipo_n58));
NAND2_X2 i_0_1_526 (.ZN (n_0_1_264), .A1 (slo__xsl_n4223), .A2 (n_0_1_265));
MUX2_X2 i_0_1_525 (.Z (n_0_1_263), .A (n_0_161), .B (n_0_55), .S (drc_ipo_n58));
INV_X4 i_0_1_524 (.ZN (n_0_1_262), .A (slo__n2712));
NAND3_X1 i_0_1_523 (.ZN (n_0_1_261), .A1 (n_0_1_264), .A2 (n_0_1_263), .A3 (sgo__n731));
OAI21_X1 i_0_1_522 (.ZN (n_0_1_260), .A (\A_imm[31] ), .B1 (slo__xsl_n4223), .B2 (n_0_1_265));
OAI21_X1 i_0_1_521 (.ZN (n_0_448), .A (n_0_1_261), .B1 (n_0_1_260), .B2 (n_0_1_263));
XNOR2_X1 i_0_1_520 (.ZN (n_0_1_259), .A (n_0_1_305), .B (n_0_1_265));
AND2_X4 i_0_1_519 (.ZN (n_0_1_258), .A1 (n_0_1_263), .A2 (n_0_1_259));
NOR2_X4 i_0_1_518 (.ZN (n_0_1_257), .A1 (n_0_1_264), .A2 (n_0_1_263));
NAND2_X4 i_0_1_517 (.ZN (n_0_1_256), .A1 (slo___n3078), .A2 (n_0_1_262));
NOR3_X1 i_0_1_516 (.ZN (n_0_1_255), .A1 (n_0_1_262), .A2 (n_0_1_265), .A3 (slo__xsl_n4223));
AOI222_X1 i_0_1_515 (.ZN (n_0_1_254), .A1 (sgo__n731), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (\A_imm[30] ), .C1 (opt_ipo_n5125), .C2 (opt_ipo_n5358));
OAI21_X1 i_0_1_514 (.ZN (n_0_447), .A (n_0_1_254), .B1 (n_0_1_256), .B2 (n_0_1_836));
AOI222_X1 i_0_1_513 (.ZN (n_0_1_253), .A1 (opt_ipo_n5358), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (\A_imm[29] ), .C1 (opt_ipo_n5125), .C2 (sgo__n1241));
OAI21_X1 i_0_1_512 (.ZN (n_0_446), .A (n_0_1_253), .B1 (n_0_1_256), .B2 (sgo__n734));
AOI222_X1 i_0_1_511 (.ZN (n_0_1_252), .A1 (sgo__n1241), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (\A_imm[28] ), .C1 (opt_ipo_n5125), .C2 (sgo__n678));
OAI21_X1 i_0_1_510 (.ZN (n_0_445), .A (n_0_1_252), .B1 (n_0_1_256), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_509 (.ZN (n_0_1_251), .A1 (sgo__n678), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (\A_imm[27] ), .C1 (opt_ipo_n5125), .C2 (sgo__n877));
OAI21_X1 i_0_1_508 (.ZN (n_0_444), .A (n_0_1_251), .B1 (n_0_1_256), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_507 (.ZN (n_0_1_250), .A1 (sgo__n877), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (slo__n1897), .C1 (opt_ipo_n5125), .C2 (sgo__n943));
OAI21_X1 i_0_1_506 (.ZN (n_0_443), .A (n_0_1_250), .B1 (n_0_1_256), .B2 (slo__n2762));
AOI222_X1 i_0_1_505 (.ZN (n_0_1_249), .A1 (sgo__n943), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (opt_ipo_n5362), .C1 (opt_ipo_n5125), .C2 (sgo__n1339));
OAI21_X1 i_0_1_504 (.ZN (n_0_442), .A (n_0_1_249), .B1 (n_0_1_256), .B2 (slo__xsl_n1889));
AOI222_X1 i_0_1_503 (.ZN (n_0_1_248), .A1 (sgo__n1339), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (slo__n2216), .C1 (opt_ipo_n5125), .C2 (slo__n1550));
OAI21_X1 i_0_1_502 (.ZN (n_0_441), .A (n_0_1_248), .B1 (n_0_1_256), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_501 (.ZN (n_0_1_247), .A1 (slo__n1550), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (slo__n3760), .C1 (opt_ipo_n5125), .C2 (sgo__n839));
OAI21_X1 i_0_1_500 (.ZN (n_0_440), .A (n_0_1_247), .B1 (n_0_1_256), .B2 (sgo__n1238));
AOI222_X1 i_0_1_499 (.ZN (n_0_1_246), .A1 (sgo__n839), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (slo__n1649), .C1 (opt_ipo_n5125), .C2 (sgo__n836));
OAI21_X1 i_0_1_498 (.ZN (n_0_439), .A (n_0_1_246), .B1 (n_0_1_256), .B2 (slo__n1812));
AOI222_X1 i_0_1_497 (.ZN (n_0_1_245), .A1 (sgo__n836), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (opt_ipo_n5135), .C1 (opt_ipo_n5125), .C2 (sgo__n1009));
OAI21_X1 i_0_1_496 (.ZN (n_0_438), .A (n_0_1_245), .B1 (n_0_1_256), .B2 (slo__xsl_n1641));
AOI222_X1 i_0_1_495 (.ZN (n_0_1_244), .A1 (sgo__n1009), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (opt_ipo_n5196), .C1 (opt_ipo_n5125), .C2 (opt_ipo_n5339));
OAI21_X1 i_0_1_494 (.ZN (n_0_437), .A (n_0_1_244), .B1 (n_0_1_256), .B2 (opt_ipo_n5145));
AOI222_X1 i_0_1_493 (.ZN (n_0_1_243), .A1 (opt_ipo_n5339), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (opt_ipo_n5303), .C1 (opt_ipo_n5125), .C2 (opt_ipo_n5373));
OAI21_X1 i_0_1_492 (.ZN (n_0_436), .A (n_0_1_243), .B1 (n_0_1_256), .B2 (opt_ipo_n5195));
AOI222_X1 i_0_1_491 (.ZN (n_0_1_242), .A1 (opt_ipo_n5373), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (slo__n2915), .C1 (opt_ipo_n5125), .C2 (\A_imm_2s_complement[18] ));
OAI21_X1 i_0_1_490 (.ZN (n_0_435), .A (n_0_1_242), .B1 (n_0_1_256), .B2 (opt_ipo_n5307));
AOI222_X2 i_0_1_489 (.ZN (n_0_1_241), .A1 (\A_imm_2s_complement[18] ), .A2 (n_0_1_258)
    , .B1 (n_0_1_257), .B2 (slo__n3402), .C1 (opt_ipo_n5411), .C2 (opt_ipo_n5125));
OAI21_X1 i_0_1_488 (.ZN (n_0_434), .A (n_0_1_241), .B1 (n_0_1_256), .B2 (slo__xsl_n1425));
AOI222_X1 i_0_1_487 (.ZN (n_0_1_240), .A1 (opt_ipo_n5411), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (slo__n3547), .C1 (opt_ipo_n5125), .C2 (opt_ipo_n5162));
OAI21_X1 i_0_1_486 (.ZN (n_0_433), .A (n_0_1_240), .B1 (n_0_1_256), .B2 (slo__xsl_n1366));
AOI222_X1 i_0_1_485 (.ZN (n_0_1_239), .A1 (sgo__n1056), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (opt_ipo_n5415), .C1 (opt_ipo_n5125), .C2 (sgo__n895));
OAI21_X1 i_0_1_484 (.ZN (n_0_432), .A (n_0_1_239), .B1 (n_0_1_256), .B2 (slo__n1493));
AOI222_X1 i_0_1_483 (.ZN (n_0_1_238), .A1 (sgo__n895), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (\A_imm[14] ), .C1 (opt_ipo_n5125), .C2 (slo__n2107));
OAI21_X1 i_0_1_482 (.ZN (n_0_431), .A (n_0_1_238), .B1 (n_0_1_256), .B2 (slo__n1828));
AOI222_X1 i_0_1_481 (.ZN (n_0_1_237), .A1 (slo__n2107), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (\A_imm[13] ), .C1 (opt_ipo_n5125), .C2 (opt_ipo_n5710));
OAI21_X1 i_0_1_480 (.ZN (n_0_430), .A (n_0_1_237), .B1 (n_0_1_256), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_479 (.ZN (n_0_1_236), .A1 (n_0_1_258), .A2 (opt_ipo_n5710), .B1 (n_0_1_257)
    , .B2 (slo__n3230), .C1 (opt_ipo_n5125), .C2 (\A_imm_2s_complement[12] ));
OAI21_X1 i_0_1_478 (.ZN (n_0_429), .A (n_0_1_236), .B1 (n_0_1_256), .B2 (slo__n1559));
AOI222_X1 i_0_1_477 (.ZN (n_0_1_235), .A1 (slo__n1702), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (opt_ipo_n5297), .C1 (slo__n3026), .C2 (opt_ipo_n5125));
OAI21_X1 i_0_1_476 (.ZN (n_0_428), .A (n_0_1_235), .B1 (n_0_1_256), .B2 (slo__n1402));
AOI222_X1 i_0_1_475 (.ZN (n_0_1_234), .A1 (slo__n3026), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (opt_ipo_n5164), .C1 (opt_ipo_n5125), .C2 (opt_ipo_n5466));
OAI21_X1 i_0_1_474 (.ZN (n_0_427), .A (n_0_1_234), .B1 (n_0_1_256), .B2 (slo___n3458));
AOI222_X1 i_0_1_473 (.ZN (n_0_1_233), .A1 (opt_ipo_n5465), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (\A_imm[9] ), .C1 (opt_ipo_n5125), .C2 (opt_ipo_n5197));
OAI21_X1 i_0_1_472 (.ZN (n_0_426), .A (n_0_1_233), .B1 (n_0_1_256), .B2 (opt_ipo_n5165));
AOI222_X1 i_0_1_471 (.ZN (n_0_1_232), .A1 (opt_ipo_n5197), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (slo__n3281), .C1 (opt_ipo_n5125), .C2 (\A_imm_2s_complement[8] ));
OAI21_X1 i_0_1_470 (.ZN (n_0_425), .A (n_0_1_232), .B1 (n_0_1_256), .B2 (n_0_1_792));
AOI222_X1 i_0_1_469 (.ZN (n_0_1_231), .A1 (slo__n2969), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (slo__n1788), .C1 (opt_ipo_n5125), .C2 (\A_imm_2s_complement[7] ));
OAI21_X1 i_0_1_468 (.ZN (n_0_424), .A (n_0_1_231), .B1 (n_0_1_256), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_467 (.ZN (n_0_1_230), .A1 (CLOCK_spw__n7292), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (spw__n7740), .C1 (opt_ipo_n5125), .C2 (opt_ipo_n5204));
OAI21_X1 i_0_1_466 (.ZN (n_0_423), .A (n_0_1_230), .B1 (n_0_1_256), .B2 (sgo__n874));
AOI222_X1 i_0_1_465 (.ZN (n_0_1_229), .A1 (opt_ipo_n5204), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (slo__n3378), .C1 (opt_ipo_n5125), .C2 (\A_imm_2s_complement[5] ));
OAI21_X1 i_0_1_464 (.ZN (n_0_422), .A (n_0_1_229), .B1 (n_0_1_256), .B2 (slo__xsl_n1694));
AOI222_X1 i_0_1_463 (.ZN (n_0_1_228), .A1 (slo__n3910), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (sgo__n962), .C1 (opt_ipo_n5125), .C2 (slo__n2805));
OAI21_X1 i_0_1_462 (.ZN (n_0_421), .A (n_0_1_228), .B1 (n_0_1_256), .B2 (n_0_1_784));
AOI222_X1 i_0_1_461 (.ZN (n_0_1_227), .A1 (slo__n2805), .A2 (n_0_1_258), .B1 (n_0_1_257)
    , .B2 (slo__n1801), .C1 (opt_ipo_n5125), .C2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_460 (.ZN (n_0_420), .A (n_0_1_227), .B1 (n_0_1_256), .B2 (sgo__n959));
AOI222_X1 i_0_1_459 (.ZN (n_0_1_226), .A1 (\A_imm_2s_complement[3] ), .A2 (n_0_1_258)
    , .B1 (n_0_1_257), .B2 (sgo__n1053), .C1 (opt_ipo_n5125), .C2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_458 (.ZN (n_0_419), .A (n_0_1_226), .B1 (n_0_1_256), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_457 (.ZN (n_0_1_225), .A1 (\A_imm_2s_complement[2] ), .A2 (n_0_1_258)
    , .B1 (n_0_1_257), .B2 (opt_ipo_n5459), .C1 (opt_ipo_n5125), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_456 (.ZN (n_0_418), .A (n_0_1_225), .B1 (n_0_1_256), .B2 (sgo__n1043));
NAND2_X1 i_0_1_455 (.ZN (n_0_1_224), .A1 (\A_imm_2s_complement[1] ), .A2 (n_0_1_258));
OAI21_X1 i_0_1_454 (.ZN (n_0_1_223), .A (sgo__n759), .B1 (n_0_1_257), .B2 (opt_ipo_n5125));
OAI211_X1 i_0_1_453 (.ZN (n_0_417), .A (n_0_1_224), .B (n_0_1_223), .C1 (n_0_1_776), .C2 (n_0_1_256));
AND2_X1 i_0_1_452 (.ZN (n_0_416), .A1 (n_0_1_259), .A2 (sgo__n759));
MUX2_X1 i_0_1_451 (.Z (n_0_1_222), .A (n_0_160), .B (n_0_56), .S (drc_ipo_n58));
NAND2_X1 i_0_1_450 (.ZN (n_0_1_221), .A1 (slo__n2712), .A2 (n_0_1_222));
NOR2_X1 slo__c1812 (.ZN (slo__n1627), .A1 (n_0_1_179), .A2 (n_0_1_220));
BUF_X1 opt_ipo_c6208 (.Z (opt_ipo_n5653), .A (\A_imm_2s_complement[15] ));
NAND3_X1 i_0_1_447 (.ZN (n_0_1_218), .A1 (n_0_1_221), .A2 (opt_ipo_n5107), .A3 (sgo__n731));
OAI21_X1 i_0_1_446 (.ZN (n_0_1_217), .A (\A_imm[31] ), .B1 (n_0_1_263), .B2 (n_0_1_222));
OAI21_X1 i_0_1_445 (.ZN (n_0_415), .A (n_0_1_218), .B1 (n_0_1_217), .B2 (opt_ipo_n5107));
XNOR2_X2 i_0_1_444 (.ZN (n_0_1_216), .A (n_0_1_262), .B (n_0_1_222));
AND2_X4 i_0_1_443 (.ZN (n_0_1_215), .A1 (n_0_1_216), .A2 (opt_ipo_n5107));
NOR2_X4 i_0_1_442 (.ZN (n_0_1_214), .A1 (n_0_1_221), .A2 (opt_ipo_n5107));
NAND2_X1 i_0_1_441 (.ZN (n_0_1_213), .A1 (n_0_1_216), .A2 (opt_ipo_n5108));
NOR3_X1 i_0_1_440 (.ZN (n_0_1_212), .A1 (opt_ipo_n5108), .A2 (n_0_1_222), .A3 (n_0_1_263));
AOI222_X1 i_0_1_439 (.ZN (n_0_1_211), .A1 (sgo__n731), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (\A_imm[30] ), .C1 (opt_ipo_n5433), .C2 (opt_ipo_n5358));
OAI21_X1 i_0_1_438 (.ZN (n_0_414), .A (n_0_1_211), .B1 (opt_ipo_n5230), .B2 (n_0_1_836));
AOI222_X1 i_0_1_437 (.ZN (n_0_1_210), .A1 (opt_ipo_n5358), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (\A_imm[29] ), .C1 (opt_ipo_n5433), .C2 (sgo__n1241));
OAI21_X1 i_0_1_436 (.ZN (n_0_413), .A (n_0_1_210), .B1 (opt_ipo_n5230), .B2 (sgo__n734));
AOI222_X1 i_0_1_435 (.ZN (n_0_1_209), .A1 (sgo__n1241), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (\A_imm[28] ), .C1 (opt_ipo_n5433), .C2 (sgo__n678));
OAI21_X1 i_0_1_434 (.ZN (n_0_412), .A (n_0_1_209), .B1 (opt_ipo_n5230), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_433 (.ZN (n_0_1_208), .A1 (sgo__n678), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (\A_imm[27] ), .C1 (opt_ipo_n5433), .C2 (sgo__n877));
OAI21_X1 i_0_1_432 (.ZN (n_0_411), .A (n_0_1_208), .B1 (opt_ipo_n5230), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_431 (.ZN (n_0_1_207), .A1 (sgo__n877), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (slo__n1897), .C1 (opt_ipo_n5433), .C2 (sgo__n943));
OAI21_X1 i_0_1_430 (.ZN (n_0_410), .A (n_0_1_207), .B1 (opt_ipo_n5230), .B2 (slo__n2762));
AOI222_X1 i_0_1_429 (.ZN (n_0_1_206), .A1 (sgo__n943), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (opt_ipo_n5362), .C1 (opt_ipo_n5433), .C2 (sgo__n1339));
OAI21_X1 i_0_1_428 (.ZN (n_0_409), .A (n_0_1_206), .B1 (opt_ipo_n5230), .B2 (slo__xsl_n1889));
AOI222_X1 i_0_1_427 (.ZN (n_0_1_205), .A1 (sgo__n1339), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (slo__n2216), .C1 (opt_ipo_n5433), .C2 (slo__n1550));
OAI21_X1 i_0_1_426 (.ZN (n_0_408), .A (n_0_1_205), .B1 (opt_ipo_n5230), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_425 (.ZN (n_0_1_204), .A1 (slo__n1550), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (slo__n3760), .C1 (opt_ipo_n5433), .C2 (sgo__n839));
OAI21_X1 i_0_1_424 (.ZN (n_0_407), .A (n_0_1_204), .B1 (opt_ipo_n5230), .B2 (sgo__n1238));
AOI222_X1 i_0_1_423 (.ZN (n_0_1_203), .A1 (sgo__n839), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (slo__n1649), .C1 (opt_ipo_n5433), .C2 (sgo__n836));
OAI21_X1 i_0_1_422 (.ZN (n_0_406), .A (n_0_1_203), .B1 (opt_ipo_n5230), .B2 (slo__n1812));
AOI222_X1 i_0_1_421 (.ZN (n_0_1_202), .A1 (sgo__n836), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (opt_ipo_n5135), .C1 (opt_ipo_n5433), .C2 (sgo__n1009));
OAI21_X1 i_0_1_420 (.ZN (n_0_405), .A (n_0_1_202), .B1 (opt_ipo_n5230), .B2 (slo__xsl_n1641));
AOI222_X1 i_0_1_419 (.ZN (n_0_1_201), .A1 (sgo__n1009), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (opt_ipo_n5196), .C1 (opt_ipo_n5433), .C2 (opt_ipo_n5339));
OAI21_X1 i_0_1_418 (.ZN (n_0_404), .A (n_0_1_201), .B1 (opt_ipo_n5230), .B2 (opt_ipo_n5145));
AOI222_X1 i_0_1_417 (.ZN (n_0_1_200), .A1 (opt_ipo_n5339), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (opt_ipo_n5303), .C1 (opt_ipo_n5433), .C2 (opt_ipo_n5373));
OAI21_X1 i_0_1_416 (.ZN (n_0_403), .A (n_0_1_200), .B1 (opt_ipo_n5230), .B2 (opt_ipo_n5195));
AOI222_X1 i_0_1_415 (.ZN (n_0_1_199), .A1 (opt_ipo_n5373), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (slo__n2915), .C1 (opt_ipo_n5433), .C2 (\A_imm_2s_complement[18] ));
OAI21_X1 i_0_1_414 (.ZN (n_0_402), .A (n_0_1_199), .B1 (opt_ipo_n5230), .B2 (opt_ipo_n5307));
AOI222_X1 i_0_1_413 (.ZN (n_0_1_198), .A1 (\A_imm_2s_complement[18] ), .A2 (slo__n1936)
    , .B1 (CLOCK_sgo__n6468), .B2 (slo__n3402), .C1 (opt_ipo_n5433), .C2 (opt_ipo_n5411));
OAI21_X1 i_0_1_412 (.ZN (n_0_401), .A (n_0_1_198), .B1 (opt_ipo_n5230), .B2 (slo__xsl_n1425));
AOI222_X1 i_0_1_411 (.ZN (n_0_1_197), .A1 (opt_ipo_n5411), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (slo__n3547), .C1 (opt_ipo_n5433), .C2 (sgo__n1056));
OAI21_X1 i_0_1_410 (.ZN (n_0_400), .A (n_0_1_197), .B1 (opt_ipo_n5230), .B2 (slo__xsl_n1366));
AOI222_X1 i_0_1_409 (.ZN (n_0_1_196), .A1 (sgo__n1056), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (opt_ipo_n5415), .C1 (opt_ipo_n5433), .C2 (sgo__n895));
OAI21_X1 i_0_1_408 (.ZN (n_0_399), .A (n_0_1_196), .B1 (opt_ipo_n5230), .B2 (slo__n1493));
AOI222_X1 i_0_1_407 (.ZN (n_0_1_195), .A1 (sgo__n895), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (\A_imm[14] ), .C1 (opt_ipo_n5433), .C2 (slo__n2107));
OAI21_X1 i_0_1_406 (.ZN (n_0_398), .A (n_0_1_195), .B1 (opt_ipo_n5230), .B2 (slo__n1828));
AOI222_X1 i_0_1_405 (.ZN (n_0_1_194), .A1 (slo__n2107), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (\A_imm[13] ), .C1 (opt_ipo_n5433), .C2 (opt_ipo_n5710));
OAI21_X1 i_0_1_404 (.ZN (n_0_397), .A (n_0_1_194), .B1 (opt_ipo_n5230), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_403 (.ZN (n_0_1_193), .A1 (opt_ipo_n5710), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (slo__n3230), .C1 (opt_ipo_n5433), .C2 (slo__n1702));
OAI21_X1 i_0_1_402 (.ZN (n_0_396), .A (n_0_1_193), .B1 (opt_ipo_n5230), .B2 (slo__n1559));
AOI222_X1 i_0_1_401 (.ZN (n_0_1_192), .A1 (slo__n1702), .A2 (n_0_1_215), .B1 (CLOCK_sgo__n6468)
    , .B2 (opt_ipo_n5297), .C1 (opt_ipo_n5433), .C2 (\A_imm_2s_complement[11] ));
OAI21_X1 i_0_1_400 (.ZN (n_0_395), .A (n_0_1_192), .B1 (opt_ipo_n5230), .B2 (slo__n1402));
AOI222_X1 i_0_1_399 (.ZN (n_0_1_191), .A1 (slo__n3026), .A2 (n_0_1_215), .B1 (CLOCK_sgo__n6468)
    , .B2 (opt_ipo_n5164), .C1 (drc_ipo_n50), .C2 (opt_ipo_n5466));
OAI21_X1 i_0_1_398 (.ZN (n_0_394), .A (n_0_1_191), .B1 (opt_ipo_n5230), .B2 (slo___n3458));
AOI222_X2 i_0_1_397 (.ZN (n_0_1_190), .A1 (opt_ipo_n5465), .A2 (slo__n1936), .B1 (CLOCK_sgo__n6468)
    , .B2 (\A_imm[9] ), .C1 (opt_ipo_n5433), .C2 (opt_ipo_n5197));
OAI21_X1 i_0_1_396 (.ZN (n_0_393), .A (n_0_1_190), .B1 (opt_ipo_n5230), .B2 (opt_ipo_n5165));
AOI222_X1 i_0_1_395 (.ZN (n_0_1_189), .A1 (opt_ipo_n5197), .A2 (n_0_1_215), .B1 (n_0_1_214)
    , .B2 (slo__n3281), .C1 (drc_ipo_n50), .C2 (\A_imm_2s_complement[8] ));
OAI21_X1 i_0_1_394 (.ZN (n_0_392), .A (n_0_1_189), .B1 (opt_ipo_n5230), .B2 (n_0_1_792));
AOI222_X1 i_0_1_393 (.ZN (n_0_1_188), .A1 (slo__n2969), .A2 (slo__n1936), .B1 (n_0_1_214)
    , .B2 (slo__n1788), .C1 (opt_ipo_n5433), .C2 (CLOCK_spw__n7292));
OAI21_X1 i_0_1_392 (.ZN (n_0_391), .A (n_0_1_188), .B1 (opt_ipo_n5230), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_391 (.ZN (n_0_1_187), .A1 (CLOCK_spw__n7292), .A2 (n_0_1_215), .B1 (n_0_1_214)
    , .B2 (spw__n7739), .C1 (drc_ipo_n50), .C2 (opt_ipo_n5205));
OAI21_X1 i_0_1_390 (.ZN (n_0_390), .A (n_0_1_187), .B1 (opt_ipo_n5230), .B2 (sgo__n874));
AOI222_X1 i_0_1_389 (.ZN (n_0_1_186), .A1 (opt_ipo_n5204), .A2 (n_0_1_215), .B1 (n_0_1_214)
    , .B2 (slo__n3378), .C1 (drc_ipo_n50), .C2 (slo__n3910));
OAI21_X1 i_0_1_388 (.ZN (n_0_389), .A (n_0_1_186), .B1 (opt_ipo_n5230), .B2 (slo__xsl_n1694));
AOI222_X1 i_0_1_387 (.ZN (n_0_1_185), .A1 (\A_imm_2s_complement[5] ), .A2 (n_0_1_215)
    , .B1 (n_0_1_214), .B2 (sgo__n962), .C1 (drc_ipo_n50), .C2 (\A_imm_2s_complement[4] ));
OAI21_X1 i_0_1_386 (.ZN (n_0_388), .A (n_0_1_185), .B1 (opt_ipo_n5230), .B2 (n_0_1_784));
AOI222_X1 i_0_1_385 (.ZN (n_0_1_184), .A1 (slo__n2805), .A2 (n_0_1_215), .B1 (n_0_1_214)
    , .B2 (slo__n1801), .C1 (drc_ipo_n50), .C2 (\A_imm_2s_complement[3] ));
OAI21_X1 i_0_1_384 (.ZN (n_0_387), .A (n_0_1_184), .B1 (opt_ipo_n5230), .B2 (sgo__n959));
AOI222_X1 i_0_1_383 (.ZN (n_0_1_183), .A1 (\A_imm_2s_complement[3] ), .A2 (n_0_1_215)
    , .B1 (n_0_1_214), .B2 (sgo__n1053), .C1 (drc_ipo_n50), .C2 (\A_imm_2s_complement[2] ));
OAI21_X1 i_0_1_382 (.ZN (n_0_386), .A (n_0_1_183), .B1 (opt_ipo_n5230), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_381 (.ZN (n_0_1_182), .A1 (\A_imm_2s_complement[2] ), .A2 (slo__n1936)
    , .B1 (n_0_1_214), .B2 (opt_ipo_n5459), .C1 (drc_ipo_n50), .C2 (\A_imm_2s_complement[1] ));
OAI21_X1 i_0_1_380 (.ZN (n_0_385), .A (n_0_1_182), .B1 (opt_ipo_n5230), .B2 (sgo__n1043));
NAND2_X1 i_0_1_379 (.ZN (n_0_1_181), .A1 (\A_imm_2s_complement[1] ), .A2 (slo__n1936));
OAI21_X1 i_0_1_378 (.ZN (n_0_1_180), .A (sgo__n759), .B1 (n_0_1_214), .B2 (opt_ipo_n5433));
OAI211_X1 i_0_1_377 (.ZN (n_0_384), .A (n_0_1_181), .B (n_0_1_180), .C1 (n_0_1_776), .C2 (opt_ipo_n5230));
AND2_X1 i_0_1_376 (.ZN (n_0_383), .A1 (n_0_1_216), .A2 (sgo__n759));
MUX2_X2 i_0_1_375 (.Z (n_0_1_179), .A (n_0_158), .B (n_0_58), .S (drc_ipo_n58));
NAND2_X1 i_0_1_374 (.ZN (n_0_1_178), .A1 (n_0_1_179), .A2 (n_0_1_220));
NAND2_X1 i_0_1_373 (.ZN (n_0_1_177), .A1 (drc_ipo_n58), .A2 (n_0_59));
NOR2_X1 i_0_1_372 (.ZN (n_0_1_176), .A1 (n_0_1_868), .A2 (drc_ipo_n58));
AOI21_X2 i_0_1_371 (.ZN (n_0_1_175), .A (n_0_1_176), .B1 (n_0_59), .B2 (drc_ipo_n58));
NAND3_X1 i_0_1_369 (.ZN (n_0_1_173), .A1 (n_0_1_178), .A2 (n_0_1_174), .A3 (sgo__n731));
BUF_X1 slo__c1840 (.Z (slo__n1649), .A (\A_imm[22] ));
NAND3_X1 i_0_1_367 (.ZN (n_0_1_171), .A1 (n_0_1_172), .A2 (n_0_1_175), .A3 (\A_imm[31] ));
NAND2_X1 i_0_1_366 (.ZN (n_0_382), .A1 (n_0_1_173), .A2 (n_0_1_171));
CLKBUF_X2 slo__c4106 (.Z (slo__n3760), .A (\A_imm[23] ));
XNOR2_X2 i_0_1_364 (.ZN (n_0_1_169), .A (opt_ipo_n5108), .B (n_0_1_179));
AND2_X4 i_0_1_363 (.ZN (n_0_1_168), .A1 (n_0_1_174), .A2 (n_0_1_169));
NOR2_X2 i_0_1_362 (.ZN (n_0_1_167), .A1 (n_0_1_172), .A2 (n_0_1_175));
AOI222_X1 i_0_1_361 (.ZN (n_0_1_166), .A1 (sgo__n731), .A2 (n_0_1_168), .B1 (slo__n1615)
    , .B2 (opt_ipo_n5358), .C1 (\A_imm[30] ), .C2 (opt_ipo_n5385));
NAND2_X1 i_0_1_360 (.ZN (n_0_1_165), .A1 (n_0_1_169), .A2 (n_0_1_175));
OAI21_X1 i_0_1_359 (.ZN (n_0_381), .A (n_0_1_166), .B1 (opt_ipo_n5103), .B2 (n_0_1_836));
AOI222_X1 i_0_1_358 (.ZN (n_0_1_164), .A1 (opt_ipo_n5358), .A2 (n_0_1_168), .B1 (slo__n1615)
    , .B2 (sgo__n1241), .C1 (\A_imm[29] ), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_357 (.ZN (n_0_380), .A (n_0_1_164), .B1 (opt_ipo_n5103), .B2 (sgo__n734));
AOI222_X1 i_0_1_356 (.ZN (n_0_1_163), .A1 (sgo__n1241), .A2 (n_0_1_168), .B1 (slo__n1615)
    , .B2 (sgo__n678), .C1 (\A_imm[28] ), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_355 (.ZN (n_0_379), .A (n_0_1_163), .B1 (opt_ipo_n5103), .B2 (slo__xsl_n1736));
AOI222_X1 i_0_1_354 (.ZN (n_0_1_162), .A1 (sgo__n678), .A2 (n_0_1_168), .B1 (slo__n1615)
    , .B2 (sgo__n877), .C1 (\A_imm[27] ), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_353 (.ZN (n_0_378), .A (n_0_1_162), .B1 (opt_ipo_n5103), .B2 (slo__xsl_n1669));
AOI222_X1 i_0_1_352 (.ZN (n_0_1_161), .A1 (sgo__n877), .A2 (n_0_1_168), .B1 (slo__n1615)
    , .B2 (sgo__n943), .C1 (slo__n1897), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_351 (.ZN (n_0_377), .A (n_0_1_161), .B1 (opt_ipo_n5103), .B2 (slo__n2762));
AOI222_X1 i_0_1_350 (.ZN (n_0_1_160), .A1 (sgo__n943), .A2 (n_0_1_168), .B1 (slo__n1615)
    , .B2 (sgo__n1339), .C1 (opt_ipo_n5362), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_349 (.ZN (n_0_376), .A (n_0_1_160), .B1 (opt_ipo_n5103), .B2 (slo__xsl_n1889));
AOI222_X1 i_0_1_348 (.ZN (n_0_1_159), .A1 (sgo__n1339), .A2 (n_0_1_168), .B1 (slo__n1615)
    , .B2 (slo__n1550), .C1 (slo__n2216), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_347 (.ZN (n_0_375), .A (n_0_1_159), .B1 (opt_ipo_n5103), .B2 (slo__xsl_n2010));
AOI222_X1 i_0_1_346 (.ZN (n_0_1_158), .A1 (slo__n1550), .A2 (n_0_1_168), .B1 (slo__n1615)
    , .B2 (sgo__n839), .C1 (slo__n3760), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_345 (.ZN (n_0_374), .A (n_0_1_158), .B1 (opt_ipo_n5103), .B2 (sgo__n1238));
AOI222_X1 i_0_1_344 (.ZN (n_0_1_157), .A1 (sgo__n839), .A2 (CLOCK_sgo__n6410), .B1 (slo__n1615)
    , .B2 (sgo__n836), .C1 (slo__n1649), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_343 (.ZN (n_0_373), .A (n_0_1_157), .B1 (opt_ipo_n5103), .B2 (slo__n1812));
AOI222_X1 i_0_1_342 (.ZN (n_0_1_156), .A1 (sgo__n836), .A2 (CLOCK_sgo__n6410), .B1 (slo__n1615)
    , .B2 (sgo__n1009), .C1 (opt_ipo_n5135), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_341 (.ZN (n_0_372), .A (n_0_1_156), .B1 (opt_ipo_n5103), .B2 (slo__xsl_n1641));
AOI222_X1 i_0_1_340 (.ZN (n_0_1_155), .A1 (sgo__n1009), .A2 (CLOCK_sgo__n6410), .B1 (slo__n1615)
    , .B2 (opt_ipo_n5339), .C1 (opt_ipo_n5196), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_339 (.ZN (n_0_371), .A (n_0_1_155), .B1 (opt_ipo_n5103), .B2 (opt_ipo_n5145));
AOI222_X1 i_0_1_338 (.ZN (n_0_1_154), .A1 (opt_ipo_n5339), .A2 (CLOCK_sgo__n6410)
    , .B1 (slo__n1615), .B2 (opt_ipo_n5373), .C1 (opt_ipo_n5303), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_337 (.ZN (n_0_370), .A (n_0_1_154), .B1 (opt_ipo_n5103), .B2 (opt_ipo_n5195));
AOI222_X1 i_0_1_336 (.ZN (n_0_1_153), .A1 (opt_ipo_n5373), .A2 (CLOCK_sgo__n6410)
    , .B1 (slo__n1615), .B2 (\A_imm_2s_complement[18] ), .C1 (slo__n2915), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_335 (.ZN (n_0_369), .A (n_0_1_153), .B1 (opt_ipo_n5103), .B2 (opt_ipo_n5307));
AOI222_X1 i_0_1_334 (.ZN (n_0_1_152), .A1 (\A_imm_2s_complement[18] ), .A2 (CLOCK_sgo__n6410)
    , .B1 (slo__n1615), .B2 (opt_ipo_n5411), .C1 (slo__n3402), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_333 (.ZN (n_0_368), .A (n_0_1_152), .B1 (opt_ipo_n5103), .B2 (slo__xsl_n1425));
AOI222_X1 i_0_1_332 (.ZN (n_0_1_151), .A1 (opt_ipo_n5411), .A2 (CLOCK_sgo__n6410)
    , .B1 (slo__n1615), .B2 (sgo__n1056), .C1 (slo__n3547), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_331 (.ZN (n_0_367), .A (n_0_1_151), .B1 (opt_ipo_n5103), .B2 (slo__xsl_n1366));
AOI222_X1 i_0_1_330 (.ZN (n_0_1_150), .A1 (sgo__n1056), .A2 (CLOCK_sgo__n6410), .B1 (slo__n1615)
    , .B2 (sgo__n895), .C1 (opt_ipo_n5415), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_329 (.ZN (n_0_366), .A (n_0_1_150), .B1 (opt_ipo_n5103), .B2 (slo__n1493));
AOI222_X1 i_0_1_328 (.ZN (n_0_1_149), .A1 (sgo__n895), .A2 (CLOCK_sgo__n6410), .B1 (slo__n1615)
    , .B2 (slo__n2107), .C1 (\A_imm[14] ), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_327 (.ZN (n_0_365), .A (n_0_1_149), .B1 (opt_ipo_n5103), .B2 (slo__n1828));
AOI222_X1 i_0_1_326 (.ZN (n_0_1_148), .A1 (slo__n2107), .A2 (CLOCK_sgo__n6410), .B1 (slo__n1615)
    , .B2 (opt_ipo_n5710), .C1 (\A_imm[13] ), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_325 (.ZN (n_0_364), .A (n_0_1_148), .B1 (opt_ipo_n5103), .B2 (slo__xsl_n4487));
AOI222_X1 i_0_1_324 (.ZN (n_0_1_147), .A1 (opt_ipo_n5710), .A2 (CLOCK_sgo__n6410)
    , .B1 (slo__n1615), .B2 (slo__n1702), .C1 (slo__n3230), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_323 (.ZN (n_0_363), .A (n_0_1_147), .B1 (opt_ipo_n5103), .B2 (slo__n1559));
AOI222_X1 i_0_1_322 (.ZN (n_0_1_146), .A1 (slo__n1702), .A2 (CLOCK_sgo__n6410), .B1 (slo__n1615)
    , .B2 (slo__n3026), .C1 (opt_ipo_n5297), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_321 (.ZN (n_0_362), .A (n_0_1_146), .B1 (opt_ipo_n5103), .B2 (slo__n1402));
AOI222_X1 i_0_1_320 (.ZN (n_0_1_145), .A1 (slo__n3026), .A2 (CLOCK_sgo__n6410), .B1 (slo__n1615)
    , .B2 (opt_ipo_n5465), .C1 (opt_ipo_n5164), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_319 (.ZN (n_0_361), .A (n_0_1_145), .B1 (opt_ipo_n5103), .B2 (slo___n3458));
AOI222_X1 i_0_1_318 (.ZN (n_0_1_144), .A1 (opt_ipo_n5465), .A2 (CLOCK_sgo__n6410)
    , .B1 (slo__n1615), .B2 (opt_ipo_n5197), .C1 (opt_ipo_n5385), .C2 (\A_imm[9] ));
OAI21_X1 i_0_1_317 (.ZN (n_0_360), .A (n_0_1_144), .B1 (opt_ipo_n5103), .B2 (opt_ipo_n5165));
AOI222_X1 i_0_1_316 (.ZN (n_0_1_143), .A1 (opt_ipo_n5197), .A2 (n_0_1_168), .B1 (slo__n1615)
    , .B2 (slo__n2969), .C1 (slo__n3281), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_315 (.ZN (n_0_359), .A (n_0_1_143), .B1 (opt_ipo_n5103), .B2 (n_0_1_792));
AOI222_X1 i_0_1_314 (.ZN (n_0_1_142), .A1 (slo__n2969), .A2 (n_0_1_168), .B1 (slo__n1615)
    , .B2 (CLOCK_spw__n7292), .C1 (slo__n1788), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_313 (.ZN (n_0_358), .A (n_0_1_142), .B1 (opt_ipo_n5103), .B2 (opt_ipo_n5794));
AOI222_X1 i_0_1_312 (.ZN (n_0_1_141), .A1 (CLOCK_spw__n7292), .A2 (n_0_1_168), .B1 (n_0_1_167)
    , .B2 (opt_ipo_n5205), .C1 (spw__n7740), .C2 (n_0_1_170));
OAI21_X1 i_0_1_311 (.ZN (n_0_357), .A (n_0_1_141), .B1 (opt_ipo_n5103), .B2 (sgo__n874));
AOI222_X1 i_0_1_310 (.ZN (n_0_1_140), .A1 (opt_ipo_n5204), .A2 (n_0_1_168), .B1 (slo__n1615)
    , .B2 (slo__n3910), .C1 (slo__n3378), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_309 (.ZN (n_0_356), .A (n_0_1_140), .B1 (opt_ipo_n5103), .B2 (slo__xsl_n1694));
AOI222_X1 i_0_1_308 (.ZN (n_0_1_139), .A1 (slo__n3910), .A2 (n_0_1_168), .B1 (n_0_1_167)
    , .B2 (slo__n2805), .C1 (sgo__n962), .C2 (n_0_1_170));
OAI21_X1 i_0_1_307 (.ZN (n_0_355), .A (n_0_1_139), .B1 (opt_ipo_n5103), .B2 (n_0_1_784));
AOI222_X1 i_0_1_306 (.ZN (n_0_1_138), .A1 (slo__n2805), .A2 (n_0_1_168), .B1 (n_0_1_167)
    , .B2 (\A_imm_2s_complement[3] ), .C1 (slo__n1801), .C2 (opt_ipo_n5385));
OAI21_X1 i_0_1_305 (.ZN (n_0_354), .A (n_0_1_138), .B1 (opt_ipo_n5103), .B2 (sgo__n959));
BUF_X2 opt_ipo_c6227 (.Z (opt_ipo_n5672), .A (\A_imm_2s_complement[14] ));
OAI21_X1 i_0_1_303 (.ZN (n_0_353), .A (n_0_1_137), .B1 (opt_ipo_n5103), .B2 (slo__xsl_n3900));
AOI222_X1 i_0_1_302 (.ZN (n_0_1_136), .A1 (\A_imm_2s_complement[2] ), .A2 (n_0_1_168)
    , .B1 (n_0_1_167), .B2 (\A_imm_2s_complement[1] ), .C1 (opt_ipo_n5459), .C2 (n_0_1_170));
OAI21_X1 i_0_1_301 (.ZN (n_0_352), .A (n_0_1_136), .B1 (opt_ipo_n5103), .B2 (sgo__n1043));
NAND2_X1 i_0_1_300 (.ZN (n_0_1_135), .A1 (\A_imm_2s_complement[1] ), .A2 (n_0_1_168));
OAI21_X1 i_0_1_299 (.ZN (n_0_1_134), .A (sgo__n759), .B1 (opt_ipo_n5385), .B2 (slo__n1615));
OAI211_X1 i_0_1_298 (.ZN (n_0_351), .A (n_0_1_135), .B (n_0_1_134), .C1 (n_0_1_776), .C2 (opt_ipo_n5103));
AND2_X1 i_0_1_297 (.ZN (n_0_350), .A1 (n_0_1_169), .A2 (sgo__n759));
NAND2_X1 i_0_1_296 (.ZN (n_0_1_133), .A1 (drc_ipo_n58), .A2 (n_0_61));
MUX2_X1 i_0_1_295 (.Z (n_0_1_132), .A (n_0_156), .B (n_0_60), .S (drc_ipo_n58));
XNOR2_X2 i_0_1_294 (.ZN (n_0_1_131), .A (n_0_1_132), .B (n_0_1_175));
INV_X1 i_0_1_293 (.ZN (n_0_1_130), .A (n_0_1_131));
NAND2_X4 i_0_1_292 (.ZN (n_0_1_129), .A1 (n_0_1_133), .A2 (n_0_1_131));
NOR2_X1 i_0_1_291 (.ZN (n_0_1_128), .A1 (n_0_1_129), .A2 (n_0_1_836));
NOR2_X2 i_0_1_290 (.ZN (n_0_1_127), .A1 (n_0_1_130), .A2 (n_0_1_133));
AOI21_X1 i_0_1_289 (.ZN (n_0_1_126), .A (n_0_1_128), .B1 (slo__n2069), .B2 (sgo__n731));
NAND3_X4 i_0_1_288 (.ZN (n_0_1_125), .A1 (n_0_1_174), .A2 (n_0_1_133), .A3 (n_0_1_132));
INV_X1 i_0_1_287 (.ZN (n_0_1_124), .A (n_0_1_125));
NOR3_X1 i_0_1_286 (.ZN (n_0_1_123), .A1 (n_0_1_133), .A2 (n_0_59), .A3 (n_0_60));
NAND2_X1 i_0_1_285 (.ZN (n_0_1_122), .A1 (sgo__n731), .A2 (drc_ipo_n56));
OAI211_X1 i_0_1_284 (.ZN (n_0_349), .A (n_0_1_126), .B (n_0_1_122), .C1 (n_0_1_125), .C2 (n_0_1_836));
AOI22_X1 i_0_1_283 (.ZN (n_0_1_121), .A1 (n_0_1_124), .A2 (\A_imm[30] ), .B1 (opt_ipo_n5358), .B2 (drc_ipo_n56));
NAND2_X1 i_0_1_282 (.ZN (n_0_348), .A1 (n_0_1_126), .A2 (n_0_1_121));
AOI22_X1 i_0_1_281 (.ZN (n_0_1_120), .A1 (opt_ipo_n5358), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (sgo__n1241));
OAI221_X1 i_0_1_280 (.ZN (n_0_347), .A (n_0_1_120), .B1 (n_0_1_125), .B2 (slo__xsl_n1736)
    , .C1 (sgo__n734), .C2 (n_0_1_129));
AOI22_X1 i_0_1_279 (.ZN (n_0_1_119), .A1 (sgo__n1241), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (sgo__n678));
OAI221_X1 i_0_1_278 (.ZN (n_0_346), .A (n_0_1_119), .B1 (n_0_1_125), .B2 (slo__xsl_n1669)
    , .C1 (slo__xsl_n1736), .C2 (n_0_1_129));
AOI22_X1 i_0_1_277 (.ZN (n_0_1_118), .A1 (sgo__n678), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (sgo__n877));
OAI221_X1 i_0_1_276 (.ZN (n_0_345), .A (n_0_1_118), .B1 (n_0_1_125), .B2 (slo__n2762)
    , .C1 (slo__xsl_n1669), .C2 (n_0_1_129));
AOI22_X1 i_0_1_275 (.ZN (n_0_1_117), .A1 (sgo__n877), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (sgo__n943));
OAI221_X1 i_0_1_274 (.ZN (n_0_344), .A (n_0_1_117), .B1 (n_0_1_125), .B2 (slo__xsl_n1889)
    , .C1 (slo__n2762), .C2 (n_0_1_129));
AOI22_X1 i_0_1_273 (.ZN (n_0_1_116), .A1 (sgo__n943), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (sgo__n1339));
OAI221_X1 i_0_1_272 (.ZN (n_0_343), .A (n_0_1_116), .B1 (n_0_1_125), .B2 (slo__xsl_n2010)
    , .C1 (slo__xsl_n1889), .C2 (n_0_1_129));
AOI22_X1 i_0_1_271 (.ZN (n_0_1_115), .A1 (sgo__n1339), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (slo__n1550));
OAI221_X1 i_0_1_270 (.ZN (n_0_342), .A (n_0_1_115), .B1 (n_0_1_125), .B2 (sgo__n1238)
    , .C1 (slo__xsl_n2010), .C2 (n_0_1_129));
AOI22_X1 i_0_1_269 (.ZN (n_0_1_114), .A1 (slo__n1550), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (sgo__n839));
OAI221_X1 i_0_1_268 (.ZN (n_0_341), .A (n_0_1_114), .B1 (n_0_1_125), .B2 (slo__n1812)
    , .C1 (sgo__n1238), .C2 (n_0_1_129));
AOI22_X1 i_0_1_267 (.ZN (n_0_1_113), .A1 (sgo__n839), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (sgo__n836));
OAI221_X1 i_0_1_266 (.ZN (n_0_340), .A (n_0_1_113), .B1 (n_0_1_125), .B2 (slo__xsl_n1641)
    , .C1 (slo__n1812), .C2 (n_0_1_129));
AOI22_X1 i_0_1_265 (.ZN (n_0_1_112), .A1 (sgo__n836), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (sgo__n1009));
OAI221_X1 i_0_1_264 (.ZN (n_0_339), .A (n_0_1_112), .B1 (n_0_1_125), .B2 (opt_ipo_n5145)
    , .C1 (slo__xsl_n1641), .C2 (n_0_1_129));
AOI22_X1 i_0_1_263 (.ZN (n_0_1_111), .A1 (sgo__n1009), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (opt_ipo_n5339));
OAI221_X1 i_0_1_262 (.ZN (n_0_338), .A (n_0_1_111), .B1 (n_0_1_125), .B2 (opt_ipo_n5195)
    , .C1 (opt_ipo_n5145), .C2 (n_0_1_129));
AOI22_X1 i_0_1_261 (.ZN (n_0_1_110), .A1 (opt_ipo_n5339), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (opt_ipo_n5373));
OAI221_X1 i_0_1_260 (.ZN (n_0_337), .A (n_0_1_110), .B1 (n_0_1_125), .B2 (opt_ipo_n5307)
    , .C1 (opt_ipo_n5195), .C2 (n_0_1_129));
AOI22_X1 i_0_1_259 (.ZN (n_0_1_109), .A1 (opt_ipo_n5373), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (\A_imm_2s_complement[18] ));
OAI221_X1 i_0_1_258 (.ZN (n_0_336), .A (n_0_1_109), .B1 (n_0_1_125), .B2 (slo__xsl_n1425)
    , .C1 (opt_ipo_n5307), .C2 (n_0_1_129));
AOI22_X1 i_0_1_257 (.ZN (n_0_1_108), .A1 (\A_imm_2s_complement[18] ), .A2 (slo__n2069)
    , .B1 (drc_ipo_n56), .B2 (opt_ipo_n5411));
OAI221_X1 i_0_1_256 (.ZN (n_0_335), .A (n_0_1_108), .B1 (n_0_1_125), .B2 (slo__xsl_n1366)
    , .C1 (slo__xsl_n1425), .C2 (n_0_1_129));
AOI22_X1 i_0_1_255 (.ZN (n_0_1_107), .A1 (opt_ipo_n5411), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (sgo__n1056));
OAI221_X1 i_0_1_254 (.ZN (n_0_334), .A (n_0_1_107), .B1 (n_0_1_125), .B2 (slo__n1493)
    , .C1 (slo__xsl_n1366), .C2 (n_0_1_129));
AOI22_X1 i_0_1_253 (.ZN (n_0_1_106), .A1 (sgo__n1056), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (sgo__n895));
OAI221_X1 i_0_1_252 (.ZN (n_0_333), .A (n_0_1_106), .B1 (n_0_1_125), .B2 (slo__n1828)
    , .C1 (slo__n1493), .C2 (n_0_1_129));
AOI22_X1 i_0_1_251 (.ZN (n_0_1_105), .A1 (sgo__n895), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (slo__n2107));
OAI221_X1 i_0_1_250 (.ZN (n_0_332), .A (n_0_1_105), .B1 (n_0_1_125), .B2 (slo__xsl_n4487)
    , .C1 (slo__n1828), .C2 (n_0_1_129));
AOI22_X1 i_0_1_249 (.ZN (n_0_1_104), .A1 (slo__n2107), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (opt_ipo_n5710));
OAI221_X1 i_0_1_248 (.ZN (n_0_331), .A (n_0_1_104), .B1 (n_0_1_125), .B2 (slo__n1559)
    , .C1 (slo__xsl_n4487), .C2 (n_0_1_129));
AOI22_X1 i_0_1_247 (.ZN (n_0_1_103), .A1 (opt_ipo_n5710), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (slo__n1702));
OAI221_X1 i_0_1_246 (.ZN (n_0_330), .A (n_0_1_103), .B1 (n_0_1_125), .B2 (slo__n1402)
    , .C1 (slo__n1559), .C2 (n_0_1_129));
AOI22_X1 i_0_1_245 (.ZN (n_0_1_102), .A1 (slo__n1702), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (slo__n3026));
OAI221_X1 i_0_1_244 (.ZN (n_0_329), .A (n_0_1_102), .B1 (n_0_1_125), .B2 (slo___n3458)
    , .C1 (slo__n1402), .C2 (n_0_1_129));
AOI22_X1 i_0_1_243 (.ZN (n_0_1_101), .A1 (slo__n3026), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (opt_ipo_n5465));
OAI221_X1 i_0_1_242 (.ZN (n_0_328), .A (n_0_1_101), .B1 (n_0_1_125), .B2 (opt_ipo_n5165)
    , .C1 (slo___n3458), .C2 (n_0_1_129));
AOI22_X1 i_0_1_241 (.ZN (n_0_1_100), .A1 (opt_ipo_n5465), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (opt_ipo_n5197));
OAI221_X1 i_0_1_240 (.ZN (n_0_327), .A (n_0_1_100), .B1 (n_0_1_125), .B2 (n_0_1_792)
    , .C1 (opt_ipo_n5165), .C2 (n_0_1_129));
AOI22_X1 i_0_1_239 (.ZN (n_0_1_99), .A1 (opt_ipo_n5197), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (slo__n2969));
OAI221_X1 i_0_1_238 (.ZN (n_0_326), .A (n_0_1_99), .B1 (n_0_1_125), .B2 (opt_ipo_n5794)
    , .C1 (n_0_1_792), .C2 (n_0_1_129));
AOI22_X1 i_0_1_237 (.ZN (n_0_1_98), .A1 (slo__n2969), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (CLOCK_spw__n7292));
OAI221_X1 i_0_1_236 (.ZN (n_0_325), .A (n_0_1_98), .B1 (n_0_1_125), .B2 (sgo__n874)
    , .C1 (opt_ipo_n5794), .C2 (n_0_1_129));
AOI22_X1 i_0_1_235 (.ZN (n_0_1_97), .A1 (CLOCK_spw__n7292), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (opt_ipo_n5204));
OAI221_X1 i_0_1_234 (.ZN (n_0_324), .A (n_0_1_97), .B1 (n_0_1_125), .B2 (slo__xsl_n1694)
    , .C1 (sgo__n874), .C2 (n_0_1_129));
AOI22_X1 i_0_1_233 (.ZN (n_0_1_96), .A1 (opt_ipo_n5204), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (slo__n3910));
OAI221_X1 i_0_1_232 (.ZN (n_0_323), .A (n_0_1_96), .B1 (n_0_1_125), .B2 (n_0_1_784)
    , .C1 (slo__xsl_n1694), .C2 (n_0_1_129));
AOI22_X1 i_0_1_231 (.ZN (n_0_1_95), .A1 (slo__n3910), .A2 (n_0_1_127), .B1 (drc_ipo_n56), .B2 (slo__n2805));
OAI221_X1 i_0_1_230 (.ZN (n_0_322), .A (n_0_1_95), .B1 (n_0_1_125), .B2 (sgo__n959)
    , .C1 (n_0_1_784), .C2 (n_0_1_129));
AOI22_X1 i_0_1_229 (.ZN (n_0_1_94), .A1 (slo__n2805), .A2 (slo__n2069), .B1 (drc_ipo_n56), .B2 (\A_imm_2s_complement[3] ));
OAI221_X1 i_0_1_228 (.ZN (n_0_321), .A (n_0_1_94), .B1 (n_0_1_125), .B2 (slo__xsl_n3900)
    , .C1 (sgo__n959), .C2 (n_0_1_129));
AOI22_X1 i_0_1_227 (.ZN (n_0_1_93), .A1 (\A_imm_2s_complement[3] ), .A2 (slo__n2069)
    , .B1 (drc_ipo_n56), .B2 (\A_imm_2s_complement[2] ));
OAI221_X1 i_0_1_226 (.ZN (n_0_320), .A (n_0_1_93), .B1 (n_0_1_125), .B2 (sgo__n1043)
    , .C1 (slo__xsl_n3900), .C2 (n_0_1_129));
AOI22_X1 i_0_1_225 (.ZN (n_0_1_92), .A1 (\A_imm_2s_complement[2] ), .A2 (n_0_1_127)
    , .B1 (drc_ipo_n56), .B2 (\A_imm_2s_complement[1] ));
OAI221_X1 i_0_1_224 (.ZN (n_0_319), .A (n_0_1_92), .B1 (n_0_1_125), .B2 (n_0_1_776)
    , .C1 (sgo__n1043), .C2 (n_0_1_129));
OAI21_X1 i_0_1_223 (.ZN (n_0_1_91), .A (sgo__n759), .B1 (n_0_1_124), .B2 (drc_ipo_n56));
OR2_X1 slo__sro_c2324 (.ZN (slo__sro_n2080), .A1 (n_0_1_129), .A2 (n_0_1_776));
BUF_X4 slo__c2352 (.Z (slo__n2107), .A (\A_imm_2s_complement[14] ));
AND2_X1 i_0_1_220 (.ZN (n_0_317), .A1 (n_0_1_131), .A2 (sgo__n759));
CLKBUF_X1 sgo__c831 (.Z (sgo__n850), .A (opt_ipo_n5664));
NOR4_X4 i_0_1_145 (.ZN (n_0_1_81), .A1 (\aggregated_res[14][36] ), .A2 (\aggregated_res[14][35] )
    , .A3 (\aggregated_res[14][34] ), .A4 (\aggregated_res[14][33] ));
NOR2_X1 sgo__sro_c761 (.ZN (sgo__sro_n801), .A1 (\aggregated_res[14][37] ), .A2 (\aggregated_res[14][38] ));
NAND2_X1 slo__sro_c1803 (.ZN (slo__sro_n1622), .A1 (n_0_57), .A2 (drc_ipo_n58));
NOR4_X1 i_0_1_141 (.ZN (n_0_1_77), .A1 (\aggregated_res[14][24] ), .A2 (\aggregated_res[14][22] )
    , .A3 (\aggregated_res[14][21] ), .A4 (\aggregated_res[14][16] ));
NOR4_X2 i_0_1_140 (.ZN (n_0_1_76), .A1 (\aggregated_res[14][20] ), .A2 (\aggregated_res[14][19] )
    , .A3 (\aggregated_res[14][18] ), .A4 (\aggregated_res[14][17] ));
CLKBUF_X1 sgo__c872 (.Z (sgo__n874), .A (n_0_1_788));
NOR4_X1 i_0_1_138 (.ZN (n_0_1_74), .A1 (\aggregated_res[14][28] ), .A2 (\aggregated_res[14][27] )
    , .A3 (\aggregated_res[14][26] ), .A4 (\aggregated_res[14][25] ));
AND2_X1 i_0_1_0 (.ZN (n_0_187), .A1 (n_0_812), .A2 (hfn_ipo_n46));
DLH_X2 \B_in_reg[0]  (.Q (n_0_186), .D (n_0_251), .G (n_0_283));
DLH_X2 \B_in_reg[1]  (.Q (n_0_185), .D (n_0_252), .G (n_0_283));
DLH_X1 \B_in_reg[2]  (.Q (n_0_184), .D (n_0_253), .G (n_0_283));
DLH_X1 \B_in_reg[3]  (.Q (n_0_183), .D (n_0_254), .G (n_0_283));
DLH_X1 \B_in_reg[4]  (.Q (n_0_182), .D (n_0_255), .G (n_0_283));
DLH_X1 \B_in_reg[5]  (.Q (n_0_181), .D (n_0_256), .G (n_0_283));
DLH_X1 \B_in_reg[6]  (.Q (n_0_180), .D (n_0_257), .G (n_0_283));
DLH_X1 \B_in_reg[7]  (.Q (n_0_179), .D (n_0_258), .G (n_0_283));
DLH_X1 \B_in_reg[8]  (.Q (n_0_178), .D (n_0_259), .G (n_0_283));
DLH_X1 \B_in_reg[9]  (.Q (n_0_177), .D (n_0_260), .G (n_0_283));
DLH_X1 \B_in_reg[10]  (.Q (n_0_176), .D (n_0_261), .G (n_0_283));
DLH_X1 \B_in_reg[11]  (.Q (n_0_175), .D (n_0_262), .G (n_0_283));
DLH_X1 \B_in_reg[12]  (.Q (n_0_174), .D (n_0_263), .G (n_0_283));
DLH_X1 \B_in_reg[13]  (.Q (n_0_173), .D (n_0_264), .G (n_0_283));
DLH_X1 \B_in_reg[14]  (.Q (n_0_172), .D (n_0_265), .G (n_0_283));
DLH_X1 \B_in_reg[15]  (.Q (n_0_171), .D (n_0_266), .G (n_0_283));
DLH_X1 \B_in_reg[16]  (.Q (n_0_170), .D (n_0_267), .G (n_0_283));
DLH_X1 \B_in_reg[17]  (.Q (n_0_169), .D (n_0_268), .G (n_0_283));
DLH_X1 \B_in_reg[18]  (.Q (n_0_168), .D (n_0_269), .G (n_0_283));
DLH_X1 \B_in_reg[19]  (.Q (n_0_167), .D (n_0_270), .G (n_0_283));
DLH_X1 \B_in_reg[20]  (.Q (n_0_166), .D (n_0_271), .G (n_0_283));
DLH_X1 \B_in_reg[21]  (.Q (n_0_165), .D (n_0_272), .G (n_0_283));
DLH_X1 \B_in_reg[22]  (.Q (n_0_164), .D (n_0_273), .G (n_0_283));
DLH_X1 \B_in_reg[23]  (.Q (n_0_163), .D (n_0_274), .G (n_0_283));
DLH_X1 \B_in_reg[24]  (.Q (n_0_162), .D (n_0_275), .G (n_0_283));
DLH_X1 \B_in_reg[25]  (.Q (n_0_161), .D (n_0_276), .G (n_0_283));
DLH_X1 \B_in_reg[26]  (.Q (n_0_160), .D (n_0_277), .G (n_0_283));
DLH_X1 \B_in_reg[27]  (.Q (n_0_159), .D (n_0_278), .G (n_0_283));
DLH_X1 \B_in_reg[28]  (.Q (n_0_158), .D (n_0_279), .G (n_0_283));
DLH_X1 \B_in_reg[29]  (.Q (n_0_157), .D (n_0_280), .G (n_0_283));
DLH_X1 \B_in_reg[30]  (.Q (n_0_156), .D (n_0_281), .G (n_0_283));
DLH_X1 \B_in_reg[31]  (.Q (B_in), .D (n_0_282), .G (n_0_283));
DLH_X2 \A_in_reg[0]  (.Q (n_0_155), .D (n_0_284), .G (n_0_283));
DLH_X2 \A_in_reg[1]  (.Q (n_0_154), .D (n_0_285), .G (n_0_283));
DLH_X2 \A_in_reg[2]  (.Q (n_0_153), .D (n_0_286), .G (n_0_283));
DLH_X2 \A_in_reg[3]  (.Q (n_0_152), .D (n_0_287), .G (n_0_283));
DLH_X1 \A_in_reg[4]  (.Q (n_0_151), .D (n_0_288), .G (n_0_283));
DLH_X1 \A_in_reg[5]  (.Q (n_0_150), .D (n_0_289), .G (n_0_283));
DLH_X1 \A_in_reg[6]  (.Q (n_0_149), .D (n_0_290), .G (n_0_283));
DLH_X1 \A_in_reg[7]  (.Q (n_0_148), .D (n_0_291), .G (n_0_283));
DLH_X2 \A_in_reg[8]  (.Q (n_0_147), .D (n_0_292), .G (n_0_283));
DLH_X1 \A_in_reg[9]  (.Q (n_0_146), .D (n_0_293), .G (n_0_283));
DLH_X2 \A_in_reg[10]  (.Q (n_0_145), .D (n_0_294), .G (n_0_283));
DLH_X1 \A_in_reg[11]  (.Q (n_0_144), .D (n_0_295), .G (n_0_283));
DLH_X1 \A_in_reg[12]  (.Q (n_0_143), .D (n_0_296), .G (n_0_283));
DLH_X1 \A_in_reg[13]  (.Q (n_0_142), .D (n_0_297), .G (n_0_283));
DLH_X1 \A_in_reg[14]  (.Q (n_0_141), .D (n_0_298), .G (n_0_283));
DLH_X1 \A_in_reg[15]  (.Q (n_0_140), .D (n_0_299), .G (n_0_283));
DLH_X2 \A_in_reg[16]  (.Q (n_0_139), .D (n_0_300), .G (n_0_283));
DLH_X1 \A_in_reg[17]  (.Q (n_0_138), .D (n_0_301), .G (n_0_283));
DLH_X1 \A_in_reg[18]  (.Q (n_0_137), .D (n_0_302), .G (n_0_283));
DLH_X1 \A_in_reg[19]  (.Q (n_0_136), .D (n_0_303), .G (n_0_283));
DLH_X2 \A_in_reg[20]  (.Q (n_0_135), .D (n_0_304), .G (n_0_283));
DLH_X1 \A_in_reg[21]  (.Q (n_0_134), .D (n_0_305), .G (n_0_283));
DLH_X1 \A_in_reg[22]  (.Q (n_0_133), .D (n_0_306), .G (n_0_283));
DLH_X1 \A_in_reg[23]  (.Q (n_0_132), .D (n_0_307), .G (n_0_283));
DLH_X1 \A_in_reg[24]  (.Q (n_0_131), .D (n_0_308), .G (n_0_283));
DLH_X1 \A_in_reg[25]  (.Q (n_0_130), .D (n_0_309), .G (n_0_283));
DLH_X1 \A_in_reg[26]  (.Q (n_0_129), .D (n_0_310), .G (n_0_283));
DLH_X1 \A_in_reg[27]  (.Q (n_0_128), .D (n_0_311), .G (n_0_283));
DLH_X1 \A_in_reg[28]  (.Q (n_0_127), .D (n_0_312), .G (n_0_283));
DLH_X1 \A_in_reg[29]  (.Q (n_0_126), .D (n_0_313), .G (n_0_283));
DLH_X1 \A_in_reg[30]  (.Q (n_0_125), .D (n_0_314), .G (n_0_283));
DLH_X2 \A_in_reg[31]  (.Q (sgo__n1251), .D (n_0_315), .G (n_0_283));
DLH_X1 \Res_reg[0]  (.Q (Res[0]), .D (n_0_187), .G (n_0_316));
DLH_X1 \Res_reg[1]  (.Q (Res[1]), .D (n_0_188), .G (n_0_316));
DLH_X1 \Res_reg[2]  (.Q (Res[2]), .D (n_0_189), .G (n_0_316));
DLH_X1 \Res_reg[3]  (.Q (Res[3]), .D (n_0_190), .G (n_0_316));
DLH_X1 \Res_reg[4]  (.Q (Res[4]), .D (n_0_191), .G (n_0_316));
DLH_X1 \Res_reg[5]  (.Q (Res[5]), .D (n_0_192), .G (n_0_316));
DLH_X1 \Res_reg[6]  (.Q (Res[6]), .D (n_0_193), .G (n_0_316));
DLH_X1 \Res_reg[7]  (.Q (Res[7]), .D (n_0_194), .G (n_0_316));
DLH_X1 \Res_reg[8]  (.Q (Res[8]), .D (n_0_195), .G (n_0_316));
DLH_X1 \Res_reg[9]  (.Q (Res[9]), .D (n_0_196), .G (n_0_316));
DLH_X1 \Res_reg[10]  (.Q (Res[10]), .D (n_0_197), .G (n_0_316));
DLH_X1 \Res_reg[11]  (.Q (Res[11]), .D (n_0_198), .G (n_0_316));
DLH_X1 \Res_reg[12]  (.Q (Res[12]), .D (n_0_199), .G (n_0_316));
DLH_X1 \Res_reg[13]  (.Q (Res[13]), .D (n_0_200), .G (n_0_316));
DLH_X1 \Res_reg[14]  (.Q (Res[14]), .D (n_0_201), .G (n_0_316));
DLH_X1 \Res_reg[15]  (.Q (Res[15]), .D (n_0_202), .G (n_0_316));
DLH_X1 \Res_reg[16]  (.Q (Res[16]), .D (n_0_203), .G (n_0_316));
DLH_X1 \Res_reg[17]  (.Q (Res[17]), .D (n_0_204), .G (n_0_316));
DLH_X1 \Res_reg[18]  (.Q (Res[18]), .D (n_0_205), .G (n_0_316));
DLH_X1 \Res_reg[19]  (.Q (Res[19]), .D (n_0_206), .G (n_0_316));
DLH_X1 \Res_reg[20]  (.Q (Res[20]), .D (n_0_207), .G (n_0_316));
DLH_X1 \Res_reg[21]  (.Q (Res[21]), .D (n_0_208), .G (n_0_316));
DLH_X1 \Res_reg[22]  (.Q (Res[22]), .D (n_0_209), .G (n_0_316));
DLH_X1 \Res_reg[23]  (.Q (Res[23]), .D (n_0_210), .G (n_0_316));
DLH_X1 \Res_reg[24]  (.Q (Res[24]), .D (n_0_211), .G (n_0_316));
DLH_X1 \Res_reg[25]  (.Q (Res[25]), .D (n_0_212), .G (n_0_316));
DLH_X1 \Res_reg[26]  (.Q (Res[26]), .D (n_0_213), .G (n_0_316));
DLH_X1 \Res_reg[27]  (.Q (Res[27]), .D (n_0_214), .G (n_0_316));
DLH_X1 \Res_reg[28]  (.Q (Res[28]), .D (n_0_215), .G (n_0_316));
DLH_X1 \Res_reg[29]  (.Q (Res[29]), .D (n_0_216), .G (n_0_316));
DLH_X1 \Res_reg[30]  (.Q (Res[30]), .D (n_0_217), .G (n_0_316));
DLH_X1 \Res_reg[31]  (.Q (Res[31]), .D (n_0_218), .G (n_0_316));
DLH_X1 \Res_reg[32]  (.Q (Res[32]), .D (n_0_219), .G (n_0_316));
DLH_X1 \Res_reg[33]  (.Q (Res[33]), .D (n_0_220), .G (n_0_316));
DLH_X1 \Res_reg[34]  (.Q (Res[34]), .D (n_0_221), .G (n_0_316));
DLH_X1 \Res_reg[35]  (.Q (Res[35]), .D (n_0_222), .G (n_0_316));
DLH_X1 \Res_reg[36]  (.Q (Res[36]), .D (n_0_223), .G (n_0_316));
DLH_X1 \Res_reg[37]  (.Q (Res[37]), .D (n_0_224), .G (n_0_316));
DLH_X1 \Res_reg[38]  (.Q (Res[38]), .D (n_0_225), .G (n_0_316));
DLH_X1 \Res_reg[39]  (.Q (Res[39]), .D (n_0_226), .G (n_0_316));
DLH_X1 \Res_reg[40]  (.Q (Res[40]), .D (n_0_227), .G (n_0_316));
DLH_X1 \Res_reg[41]  (.Q (Res[41]), .D (n_0_228), .G (n_0_316));
DLH_X1 \Res_reg[42]  (.Q (Res[42]), .D (n_0_229), .G (n_0_316));
DLH_X1 \Res_reg[43]  (.Q (Res[43]), .D (n_0_230), .G (n_0_316));
DLH_X1 \Res_reg[44]  (.Q (Res[44]), .D (n_0_231), .G (n_0_316));
DLH_X1 \Res_reg[45]  (.Q (Res[45]), .D (n_0_232), .G (n_0_316));
DLH_X1 \Res_reg[46]  (.Q (Res[46]), .D (n_0_233), .G (n_0_316));
DLH_X1 \Res_reg[47]  (.Q (Res[47]), .D (n_0_234), .G (n_0_316));
DLH_X1 \Res_reg[48]  (.Q (Res[48]), .D (n_0_235), .G (n_0_316));
DLH_X1 \Res_reg[49]  (.Q (Res[49]), .D (n_0_236), .G (n_0_316));
DLH_X1 \Res_reg[50]  (.Q (Res[50]), .D (n_0_237), .G (n_0_316));
DLH_X1 \Res_reg[51]  (.Q (Res[51]), .D (n_0_238), .G (n_0_316));
DLH_X1 \Res_reg[52]  (.Q (Res[52]), .D (n_0_239), .G (n_0_316));
DLH_X1 \Res_reg[53]  (.Q (Res[53]), .D (n_0_240), .G (n_0_316));
DLH_X2 \Res_reg[54]  (.Q (Res[54]), .D (n_0_241), .G (n_0_316));
DLH_X1 \Res_reg[55]  (.Q (Res[55]), .D (n_0_242), .G (n_0_316));
DLH_X1 \Res_reg[56]  (.Q (Res[56]), .D (n_0_243), .G (n_0_316));
DLH_X1 \Res_reg[57]  (.Q (Res[57]), .D (n_0_244), .G (n_0_316));
DLH_X2 \Res_reg[58]  (.Q (Res[58]), .D (n_0_245), .G (n_0_316));
DLH_X1 \Res_reg[59]  (.Q (Res[59]), .D (n_0_246), .G (n_0_316));
DLH_X1 \Res_reg[60]  (.Q (Res[60]), .D (n_0_247), .G (n_0_316));
DLH_X1 \Res_reg[61]  (.Q (Res[61]), .D (n_0_248), .G (n_0_316));
DLH_X1 \Res_reg[62]  (.Q (Res[62]), .D (n_0_249), .G (n_0_316));
DLH_X2 \Res_reg[63]  (.Q (opt_ipo_n5239), .D (n_0_250), .G (n_0_316));
datapath__0_68 i_0_6 (.p_0 ({n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, 
    n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, 
    n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, 
    n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, 
    n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, 
    n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, 
    n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, uc_503})
    , .\aggregated_res[14]  ({\aggregated_res[14][63] , \aggregated_res[14][62] , 
    \aggregated_res[14][61] , \aggregated_res[14][60] , \aggregated_res[14][59] , 
    \aggregated_res[14][58] , \aggregated_res[14][57] , \aggregated_res[14][56] , 
    \aggregated_res[14][55] , \aggregated_res[14][54] , \aggregated_res[14][53] , 
    \aggregated_res[14][52] , \aggregated_res[14][51] , \aggregated_res[14][50] , 
    \aggregated_res[14][49] , \aggregated_res[14][48] , \aggregated_res[14][47] , 
    \aggregated_res[14][46] , \aggregated_res[14][45] , \aggregated_res[14][44] , 
    \aggregated_res[14][43] , \aggregated_res[14][42] , \aggregated_res[14][41] , 
    \aggregated_res[14][40] , \aggregated_res[14][39] , \aggregated_res[14][38] , 
    \aggregated_res[14][37] , \aggregated_res[14][36] , \aggregated_res[14][35] , 
    \aggregated_res[14][34] , \aggregated_res[14][33] , \aggregated_res[14][32] , 
    \aggregated_res[14][31] , \aggregated_res[14][30] , \aggregated_res[14][29] , 
    \aggregated_res[14][28] , \aggregated_res[14][27] , \aggregated_res[14][26] , 
    \aggregated_res[14][25] , \aggregated_res[14][24] , \aggregated_res[14][23] , 
    \aggregated_res[14][22] , \aggregated_res[14][21] , \aggregated_res[14][20] , 
    \aggregated_res[14][19] , \aggregated_res[14][18] , \aggregated_res[14][17] , 
    \aggregated_res[14][16] , \aggregated_res[14][15] , \aggregated_res[14][14] , 
    \aggregated_res[14][13] , \aggregated_res[14][12] , \aggregated_res[14][11] , 
    \aggregated_res[14][10] , \aggregated_res[14][9] , \aggregated_res[14][8] , \aggregated_res[14][7] , 
    \aggregated_res[14][6] , \aggregated_res[14][5] , \aggregated_res[14][4] , \aggregated_res[14][3] , 
    \aggregated_res[14][2] , n_0_813, n_0_812}));
datapath__0_67 i_0_5 (.\aggregated_res[14]  ({\aggregated_res[14][63] , \aggregated_res[14][62] , 
    \aggregated_res[14][61] , \aggregated_res[14][60] , \aggregated_res[14][59] , 
    \aggregated_res[14][58] , \aggregated_res[14][57] , \aggregated_res[14][56] , 
    \aggregated_res[14][55] , \aggregated_res[14][54] , \aggregated_res[14][53] , 
    \aggregated_res[14][52] , \aggregated_res[14][51] , \aggregated_res[14][50] , 
    \aggregated_res[14][49] , \aggregated_res[14][48] , \aggregated_res[14][47] , 
    \aggregated_res[14][46] , \aggregated_res[14][45] , \aggregated_res[14][44] , 
    \aggregated_res[14][43] , \aggregated_res[14][42] , \aggregated_res[14][41] , 
    \aggregated_res[14][40] , \aggregated_res[14][39] , \aggregated_res[14][38] , 
    \aggregated_res[14][37] , \aggregated_res[14][36] , \aggregated_res[14][35] , 
    \aggregated_res[14][34] , \aggregated_res[14][33] , \aggregated_res[14][32] , 
    \aggregated_res[14][31] , \aggregated_res[14][30] , \aggregated_res[14][29] , 
    \aggregated_res[14][28] , \aggregated_res[14][27] , \aggregated_res[14][26] , 
    \aggregated_res[14][25] , \aggregated_res[14][24] , \aggregated_res[14][23] , 
    \aggregated_res[14][22] , \aggregated_res[14][21] , \aggregated_res[14][20] , 
    \aggregated_res[14][19] , \aggregated_res[14][18] , \aggregated_res[14][17] , 
    \aggregated_res[14][16] , \aggregated_res[14][15] , \aggregated_res[14][14] , 
    \aggregated_res[14][13] , \aggregated_res[14][12] , \aggregated_res[14][11] , 
    \aggregated_res[14][10] , \aggregated_res[14][9] , \aggregated_res[14][8] , \aggregated_res[14][7] , 
    \aggregated_res[14][6] , \aggregated_res[14][5] , \aggregated_res[14][4] , \aggregated_res[14][3] , 
    \aggregated_res[14][2] , uc_501, uc_502}), .p_0 ({uc_3, uc_4, uc_5, uc_6, uc_7, 
    uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, 
    uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, 
    uc_31, n_0_811, n_0_810, n_0_809, n_0_808, sgo__sro_n1289, n_0_806, n_0_805, 
    n_0_804, n_0_803, n_0_802, n_0_801, n_0_800, n_0_799, n_0_798, n_0_797, n_0_796, 
    n_0_795, n_0_794, n_0_793, n_0_792, n_0_791, n_0_790, n_0_789, n_0_788, n_0_787, 
    n_0_786, n_0_785, n_0_784, n_0_783, n_0_782, n_0_781, n_0_780, n_0_779, uc_32, 
    uc_33}), .p_10 ({uc_313, uc_314, uc_315, uc_316, uc_317, uc_318, uc_319, uc_320, 
    uc_321, n_0_481, n_0_480, n_0_479, n_0_478, n_0_477, n_0_476, n_0_475, n_0_474, 
    n_0_473, n_0_472, n_0_471, n_0_470, n_0_469, n_0_468, n_0_467, n_0_466, n_0_465, 
    n_0_464, n_0_463, n_0_462, n_0_461, n_0_460, n_0_459, n_0_458, n_0_457, n_0_456, 
    n_0_455, n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, uc_322, uc_323, 
    uc_324, uc_325, uc_326, uc_327, uc_328, uc_329, uc_330, uc_331, uc_332, uc_333, 
    uc_334, uc_335, uc_336, uc_337, uc_338, uc_339, uc_340, uc_341, uc_342, uc_343})
    , .p_11 ({uc_344, uc_345, uc_346, uc_347, uc_348, uc_349, uc_350, n_0_448, n_0_447, 
    n_0_446, n_0_445, n_0_444, n_0_443, n_0_442, n_0_441, n_0_440, n_0_439, n_0_438, 
    n_0_437, n_0_436, n_0_435, n_0_434, n_0_433, n_0_432, n_0_431, n_0_430, n_0_429, 
    n_0_428, n_0_427, n_0_426, n_0_425, n_0_424, n_0_423, n_0_422, n_0_421, n_0_420, 
    n_0_419, n_0_418, n_0_417, n_0_416, uc_351, uc_352, uc_353, uc_354, uc_355, uc_356, 
    uc_357, uc_358, uc_359, uc_360, uc_361, uc_362, uc_363, uc_364, uc_365, uc_366, 
    uc_367, uc_368, uc_369, uc_370, uc_371, uc_372, uc_373, uc_374}), .p_12 ({uc_375, 
    uc_376, uc_377, uc_378, uc_379, n_0_415, n_0_414, n_0_413, n_0_412, n_0_411, 
    n_0_410, n_0_409, n_0_408, n_0_407, n_0_406, n_0_405, n_0_404, n_0_403, n_0_402, 
    n_0_401, n_0_400, n_0_399, n_0_398, n_0_397, n_0_396, n_0_395, n_0_394, n_0_393, 
    n_0_392, n_0_391, n_0_390, n_0_389, n_0_388, n_0_387, n_0_386, n_0_385, n_0_384, 
    n_0_383, uc_380, uc_381, uc_382, uc_383, uc_384, uc_385, uc_386, uc_387, uc_388, 
    uc_389, uc_390, uc_391, uc_392, uc_393, uc_394, uc_395, uc_396, uc_397, uc_398, 
    uc_399, uc_400, uc_401, uc_402, uc_403, uc_404, uc_405}), .p_13 ({uc_406, uc_407, 
    uc_408, n_0_382, n_0_381, n_0_380, n_0_379, n_0_378, n_0_377, n_0_376, n_0_375, 
    n_0_374, n_0_373, n_0_372, n_0_371, n_0_370, n_0_369, n_0_368, n_0_367, n_0_366, 
    n_0_365, n_0_364, n_0_363, n_0_362, n_0_361, n_0_360, n_0_359, n_0_358, n_0_357, 
    n_0_356, n_0_355, n_0_354, n_0_353, n_0_352, n_0_351, n_0_350, uc_409, uc_410, 
    uc_411, uc_412, uc_413, uc_414, uc_415, uc_416, uc_417, uc_418, uc_419, uc_420, 
    uc_421, uc_422, uc_423, uc_424, uc_425, uc_426, uc_427, uc_428, uc_429, uc_430, 
    uc_431, uc_432, uc_433, uc_434, uc_435, uc_436}), .p_14 ({uc_437, n_0_349, n_0_348, 
    n_0_347, n_0_346, n_0_345, n_0_344, n_0_343, n_0_342, n_0_341, n_0_340, n_0_339, 
    n_0_338, n_0_337, n_0_336, n_0_335, n_0_334, n_0_333, n_0_332, n_0_331, n_0_330, 
    n_0_329, n_0_328, n_0_327, n_0_326, n_0_325, n_0_324, n_0_323, n_0_322, n_0_321, 
    n_0_320, n_0_319, slo__sro_n2079, n_0_317, uc_438, uc_439, uc_440, uc_441, uc_442, 
    uc_443, uc_444, uc_445, uc_446, uc_447, uc_448, uc_449, uc_450, uc_451, uc_452, 
    uc_453, uc_454, uc_455, uc_456, uc_457, uc_458, uc_459, uc_460, uc_461, uc_462, 
    uc_463, uc_464, uc_465, uc_466, uc_467}), .p_15 ({uc_468, uc_469, uc_470, uc_471, 
    uc_472, uc_473, uc_474, uc_475, uc_476, uc_477, uc_478, uc_479, uc_480, uc_481, 
    uc_482, uc_483, uc_484, uc_485, uc_486, uc_487, uc_488, uc_489, uc_490, uc_491, 
    uc_492, uc_493, uc_494, uc_495, uc_496, uc_497, uc_498, n_0_844, n_0_843, n_0_842, 
    n_0_841, n_0_840, n_0_839, n_0_838, n_0_837, n_0_836, slo__sro_n3406, n_0_834, 
    n_0_833, n_0_832, n_0_831, n_0_830, n_0_829, CLOCK_slo__sro_n6808, n_0_827, n_0_826, 
    n_0_825, n_0_824, n_0_823, n_0_822, n_0_821, n_0_820, n_0_819, n_0_818, n_0_817, 
    n_0_816, n_0_815, n_0_814, uc_499, uc_500}), .p_1 ({uc_34, uc_35, uc_36, uc_37, 
    uc_38, uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, 
    uc_49, uc_50, uc_51, uc_52, uc_53, uc_54, uc_55, uc_56, uc_57, uc_58, uc_59, 
    uc_60, n_0_778, n_0_777, n_0_776, n_0_775, n_0_774, n_0_773, n_0_772, n_0_771, 
    n_0_770, n_0_769, n_0_768, n_0_767, n_0_766, n_0_765, CLOCK_slo__sro_n6740, n_0_763, 
    n_0_762, n_0_761, n_0_760, n_0_759, n_0_758, n_0_757, n_0_756, n_0_755, n_0_754, 
    n_0_753, n_0_752, n_0_751, n_0_750, n_0_749, n_0_748, n_0_747, n_0_746, uc_61, 
    uc_62, uc_63, uc_64}), .p_2 ({uc_65, uc_66, uc_67, uc_68, uc_69, uc_70, uc_71, 
    uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, uc_79, uc_80, uc_81, uc_82, 
    uc_83, uc_84, uc_85, uc_86, uc_87, uc_88, uc_89, n_0_745, n_0_744, n_0_743, n_0_742, 
    n_0_741, n_0_740, n_0_739, n_0_738, n_0_737, n_0_736, n_0_735, n_0_734, n_0_733, 
    n_0_732, n_0_731, n_0_730, n_0_729, n_0_728, n_0_727, n_0_726, n_0_725, n_0_724, 
    n_0_723, n_0_722, n_0_721, n_0_720, n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
    n_0_714, n_0_713, uc_90, uc_91, uc_92, uc_93, uc_94, uc_95}), .p_3 ({uc_96, uc_97, 
    uc_98, uc_99, uc_100, uc_101, uc_102, uc_103, uc_104, uc_105, uc_106, uc_107, 
    uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, uc_114, uc_115, uc_116, uc_117, 
    uc_118, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, n_0_706, n_0_705, 
    n_0_704, n_0_703, n_0_702, n_0_701, n_0_700, n_0_699, n_0_698, n_0_697, n_0_696, 
    n_0_695, n_0_694, n_0_693, n_0_692, n_0_691, slo__sro_n1594, n_0_689, n_0_688, 
    n_0_687, n_0_686, n_0_685, n_0_684, n_0_683, n_0_682, n_0_681, n_0_680, uc_119, 
    uc_120, uc_121, uc_122, uc_123, uc_124, uc_125, uc_126}), .p_4 ({uc_127, uc_128, 
    uc_129, uc_130, uc_131, uc_132, uc_133, uc_134, uc_135, uc_136, uc_137, uc_138, 
    uc_139, uc_140, uc_141, uc_142, uc_143, uc_144, uc_145, uc_146, uc_147, n_0_679, 
    n_0_678, n_0_677, n_0_676, n_0_675, n_0_674, n_0_673, n_0_672, n_0_671, n_0_670, 
    n_0_669, n_0_668, n_0_667, n_0_666, n_0_665, n_0_664, n_0_663, n_0_662, n_0_661, 
    n_0_660, n_0_659, n_0_658, n_0_657, n_0_656, n_0_655, n_0_654, n_0_653, n_0_652, 
    n_0_651, n_0_650, n_0_649, n_0_648, n_0_647, uc_148, uc_149, uc_150, uc_151, 
    uc_152, uc_153, uc_154, uc_155, uc_156, uc_157}), .p_5 ({uc_158, uc_159, uc_160, 
    uc_161, uc_162, uc_163, uc_164, uc_165, uc_166, uc_167, uc_168, uc_169, uc_170, 
    uc_171, uc_172, uc_173, uc_174, uc_175, uc_176, n_0_646, n_0_645, n_0_644, n_0_643, 
    n_0_642, n_0_641, n_0_640, n_0_639, n_0_638, n_0_637, n_0_636, n_0_635, n_0_634, 
    n_0_633, n_0_632, n_0_631, n_0_630, n_0_629, n_0_628, n_0_627, n_0_626, n_0_625, 
    n_0_624, n_0_623, n_0_622, n_0_621, n_0_620, n_0_619, n_0_618, n_0_617, n_0_616, 
    n_0_615, n_0_614, uc_177, uc_178, uc_179, uc_180, uc_181, uc_182, uc_183, uc_184, 
    uc_185, uc_186, uc_187, uc_188}), .p_6 ({uc_189, uc_190, uc_191, uc_192, uc_193, 
    uc_194, uc_195, uc_196, uc_197, uc_198, uc_199, uc_200, uc_201, uc_202, uc_203, 
    uc_204, uc_205, n_0_613, n_0_612, n_0_611, n_0_610, n_0_609, n_0_608, n_0_607, 
    n_0_606, n_0_605, n_0_604, n_0_603, n_0_602, n_0_601, n_0_600, n_0_599, n_0_598, 
    n_0_597, n_0_596, n_0_595, n_0_594, n_0_593, n_0_592, n_0_591, n_0_590, n_0_589, 
    n_0_588, n_0_587, n_0_586, n_0_585, n_0_584, n_0_583, n_0_582, n_0_581, uc_206, 
    uc_207, uc_208, uc_209, uc_210, uc_211, uc_212, uc_213, uc_214, uc_215, uc_216, 
    uc_217, uc_218, uc_219}), .p_7 ({uc_220, uc_221, uc_222, uc_223, uc_224, uc_225, 
    uc_226, uc_227, uc_228, uc_229, uc_230, uc_231, uc_232, uc_233, uc_234, n_0_580, 
    n_0_579, n_0_578, n_0_577, n_0_576, n_0_575, n_0_574, n_0_573, n_0_572, n_0_571, 
    n_0_570, n_0_569, n_0_568, n_0_567, n_0_566, n_0_565, n_0_564, n_0_563, n_0_562, 
    n_0_561, n_0_560, n_0_559, n_0_558, n_0_557, n_0_556, n_0_555, n_0_554, n_0_553, 
    n_0_552, n_0_551, n_0_550, n_0_549, n_0_548, uc_235, uc_236, uc_237, uc_238, 
    uc_239, uc_240, uc_241, uc_242, uc_243, uc_244, uc_245, uc_246, uc_247, uc_248, 
    uc_249, uc_250}), .p_8 ({uc_251, uc_252, uc_253, uc_254, uc_255, uc_256, uc_257, 
    uc_258, uc_259, uc_260, uc_261, uc_262, uc_263, n_0_547, n_0_546, n_0_545, n_0_544, 
    n_0_543, n_0_542, n_0_541, n_0_540, n_0_539, n_0_538, n_0_537, n_0_536, n_0_535, 
    n_0_534, n_0_533, n_0_532, n_0_531, n_0_530, n_0_529, n_0_528, n_0_527, n_0_526, 
    n_0_525, n_0_524, n_0_523, n_0_522, n_0_521, n_0_520, n_0_519, n_0_518, n_0_517, 
    n_0_516, n_0_515, uc_264, uc_265, uc_266, uc_267, uc_268, uc_269, uc_270, uc_271, 
    uc_272, uc_273, uc_274, uc_275, uc_276, uc_277, uc_278, uc_279, uc_280, uc_281})
    , .p_9 ({uc_282, uc_283, uc_284, uc_285, uc_286, uc_287, uc_288, uc_289, uc_290, 
    uc_291, uc_292, n_0_514, n_0_513, n_0_512, n_0_511, n_0_510, n_0_509, n_0_508, 
    n_0_507, n_0_506, n_0_505, n_0_504, n_0_503, n_0_502, n_0_501, n_0_500, n_0_499, 
    n_0_498, n_0_497, n_0_496, n_0_495, n_0_494, n_0_493, n_0_492, n_0_491, n_0_490, 
    n_0_489, n_0_488, n_0_487, n_0_486, n_0_485, n_0_484, n_0_483, n_0_482, uc_293, 
    uc_294, uc_295, uc_296, uc_297, uc_298, uc_299, uc_300, uc_301, uc_302, uc_303, 
    uc_304, uc_305, uc_306, uc_307, uc_308, uc_309, uc_310, uc_311, uc_312}));
datapath__0_1 i_0_3 (.p_0 ({n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, 
    n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, 
    n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, 
    n_0_34, n_0_33, n_0_32, n_0_31, uc_2}), .B_in ({drc_ipo_n58, n_0_156, n_0_157, 
    n_0_158, n_0_159, n_0_160, n_0_161, n_0_162, n_0_163, n_0_164, n_0_165, n_0_166, 
    n_0_167, n_0_168, n_0_169, n_0_170, n_0_171, n_0_172, n_0_173, n_0_174, n_0_175, 
    n_0_176, n_0_177, n_0_178, n_0_179, n_0_180, n_0_181, n_0_182, n_0_183, n_0_184, 
    n_0_185, n_0_186}));
datapath__0_0 i_0_2 (.A_imm_2s_complement ({\A_imm_2s_complement[31] , \A_imm_2s_complement[30] , 
    \A_imm_2s_complement[29] , \A_imm_2s_complement[28] , \A_imm_2s_complement[27] , 
    \A_imm_2s_complement[26] , \A_imm_2s_complement[25] , \A_imm_2s_complement[24] , 
    \A_imm_2s_complement[23] , \A_imm_2s_complement[22] , \A_imm_2s_complement[21] , 
    \A_imm_2s_complement[20] , \A_imm_2s_complement[19] , \A_imm_2s_complement[18] , 
    \A_imm_2s_complement[17] , \A_imm_2s_complement[16] , \A_imm_2s_complement[15] , 
    \A_imm_2s_complement[14] , \A_imm_2s_complement[13] , \A_imm_2s_complement[12] , 
    \A_imm_2s_complement[11] , \A_imm_2s_complement[10] , \A_imm_2s_complement[9] , 
    \A_imm_2s_complement[8] , \A_imm_2s_complement[7] , \A_imm_2s_complement[6] , 
    \A_imm_2s_complement[5] , \A_imm_2s_complement[4] , \A_imm_2s_complement[3] , 
    \A_imm_2s_complement[2] , \A_imm_2s_complement[1] , uc_1}), .A_imm ({\A_imm[31] , 
    \A_imm[30] , \A_imm[29] , \A_imm[28] , \A_imm[27] , n_0_1_826, sgo__n880, \A_imm[24] , 
    \A_imm[23] , \A_imm[22] , opt_ipo_n5146, n_0_1_814, n_0_1_812, \A_imm[18] , opt_ipo_n5191, 
    \A_imm[16] , opt_ipo_n5417, \A_imm[14] , \A_imm[13] , \A_imm[12] , n_0_1_796, 
    n_0_1_794, \A_imm[9] , opt_ipo_n5795, \A_imm[7] , spw__n7741, slo__sro_n3368, 
    \A_imm[4] , \A_imm[3] , \A_imm[2] , \A_imm[1] , sgo__n759}), .opt_ipoPP_2 (opt_ipo_n5145)
    , .opt_ipoPP_3 (opt_ipo_n5165), .opt_ipoPP_6 (opt_ipo_n5195), .opt_ipoPP_7 (opt_ipo_n5196)
    , .opt_ipoPP_8 (opt_ipo_n5208), .opt_ipoPP_12 (opt_ipo_n5297), .opt_ipoPP_13 (opt_ipo_n5303)
    , .opt_ipoPP_14 (opt_ipo_n5362), .opt_ipoPP_15 (sgo__n880), .opt_ipoPP_17 (opt_ipo_n5415)
    , .opt_ipoPP_20 (\A_imm[14] ), .opt_ipoPP_21 (n_0_1_796), .opt_ipoPP_22 (opt_ipo_n5794));
datapath i_0_0 (.p_0 ({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, 
    n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, 
    n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, 
    n_0_1, n_0_0, uc_0}), .A_in ({A_in, n_0_125, n_0_126, n_0_127, n_0_128, n_0_129, 
    n_0_130, n_0_131, n_0_132, n_0_133, n_0_134, n_0_135, n_0_136, n_0_137, n_0_138, 
    n_0_139, n_0_140, opt_ipo_n5712, n_0_142, n_0_143, n_0_144, n_0_145, n_0_146, 
    n_0_147, n_0_148, opt_ipo_n5703, n_0_150, n_0_151, n_0_152, n_0_153, n_0_154, 
    drc_ipo_n59}), .opt_ipoPP_1 (n_0_134), .opt_ipoPP_13 (opt_ipo_n5702), .opt_ipoPP_14 (opt_ipo_n5711));
BUF_X16 hfn_ipo_c44 (.Z (hfn_ipo_n44), .A (n_0_1_752));
CLKBUF_X1 hfn_ipo_c45 (.Z (hfn_ipo_n45), .A (n_0_1_970));
BUF_X8 drc_ipo_c58 (.Z (drc_ipo_n58), .A (B_in));
BUF_X16 hfn_ipo_c41 (.Z (hfn_ipo_n41), .A (A_in));
CLKBUF_X3 opt_ipo_c5719 (.Z (opt_ipo_n5135), .A (sgo__n850));
BUF_X4 drc_ipo_c52 (.Z (drc_ipo_n52), .A (n_0_1_513));
INV_X8 opt_ipo_c5780 (.ZN (opt_ipo_n5196), .A (n_0_1_814));
BUF_X8 drc_ipo_c50 (.Z (drc_ipo_n50), .A (n_0_1_212));
BUF_X8 drc_ipo_c59 (.Z (drc_ipo_n59), .A (n_0_155));
BUF_X4 drc_ipo_c56 (.Z (drc_ipo_n56), .A (n_0_1_123));
CLKBUF_X1 sph__c8608 (.Z (sph__n7810), .A (sph__n7809));
BUF_X8 drc_ipo_c54 (.Z (drc_ipo_n54), .A (n_0_1_427));
BUF_X16 drc_ipo_c53 (.Z (drc_ipo_n53), .A (n_0_1_470));
BUF_X16 drc_ipo_c48 (.Z (drc_ipo_n48), .A (n_0_1_298));
BUF_X4 sgo__c600 (.Z (sgo__n678), .A (\A_imm_2s_complement[28] ));
BUF_X16 hfn_ipo_c46 (.Z (hfn_ipo_n46), .A (n_0_1_970));
BUF_X2 sgo__c672 (.Z (sgo__n731), .A (\A_imm_2s_complement[31] ));
BUF_X4 slo__c5515 (.Z (slo__n4931), .A (n_0_1_920));
NAND2_X4 sgo__sro_c724 (.ZN (sgo__sro_n772), .A1 (drc_ipo_n54), .A2 (\A_imm_2s_complement[2] ));
NAND2_X1 sgo__sro_c725 (.ZN (sgo__sro_n771), .A1 (sgo__n1053), .A2 (n_0_1_429));
INV_X1 sgo__sro_c681 (.ZN (sgo__sro_n741), .A (slo__sro_n3170));
NOR2_X1 sgo__sro_c624 (.ZN (sgo__sro_n697), .A1 (\aggregated_res[14][41] ), .A2 (\aggregated_res[14][42] ));
NAND2_X1 CLOCK_slo__sro_c7554 (.ZN (CLOCK_slo__sro_n6808), .A1 (n_0_1_953), .A2 (CLOCK_slo__sro_n6809));
BUF_X2 spw__L2_c8529 (.Z (spw__n7730), .A (spw__n7729));
NOR2_X2 sgo__sro_c683 (.ZN (sgo__sro_n739), .A1 (n_0_1_877), .A2 (n_0_1_871));
BUF_X8 sgo__c957 (.Z (sgo__n943), .A (\A_imm_2s_complement[26] ));
INV_X1 sgo__sro_c637 (.ZN (sgo__sro_n705), .A (\aggregated_res[14][29] ));
NOR2_X1 sgo__sro_c638 (.ZN (sgo__sro_n704), .A1 (\aggregated_res[14][30] ), .A2 (\aggregated_res[14][23] ));
NAND2_X1 sgo__sro_c639 (.ZN (sgo__sro_n703), .A1 (sgo__sro_n704), .A2 (sgo__sro_n705));
NOR2_X4 sgo__sro_c640 (.ZN (sgo__sro_n702), .A1 (\aggregated_res[14][63] ), .A2 (sgo__sro_n703));
AOI21_X2 sgo__sro_c727 (.ZN (sgo__sro_n769), .A (sgo__sro_n770), .B1 (n_0_1_430), .B2 (\A_imm_2s_complement[3] ));
BUF_X4 sgo__c734 (.Z (sgo__n779), .A (n_0_1_430));
CLKBUF_X1 CLOCK_slh__c7890 (.Z (CLOCK_slh__n7180), .A (CLOCK_slh__n7179));
CLKBUF_X1 CLOCK_slh__c7913 (.Z (CLOCK_slh__n7206), .A (CLOCK_slh__n7202));
AND2_X1 sgo__sro_c660 (.ZN (sgo__sro_n722), .A1 (n_0_1_74), .A2 (n_0_1_77));
CLKBUF_X1 CLOCK_slh__c7911 (.Z (CLOCK_slh__n7201), .A (CLOCK_slh__n7200));
INV_X2 sgo__sro_c662 (.ZN (sgo__sro_n720), .A (CLOCK_slo__mro_n6798));
NAND2_X2 sgo__sro_c663 (.ZN (sgo__sro_n719), .A1 (sgo__sro_n720), .A2 (n_0_1_81));
NOR4_X2 sgo__c716 (.ZN (n_0_1_876), .A1 (\aggregated_res[14][53] ), .A2 (\aggregated_res[14][54] )
    , .A3 (\aggregated_res[14][51] ), .A4 (\aggregated_res[14][52] ));
NOR2_X1 sgo__sro_c762 (.ZN (sgo__sro_n800), .A1 (\aggregated_res[14][46] ), .A2 (\aggregated_res[14][40] ));
AND2_X2 sgo__sro_c763 (.ZN (sgo__sro_n799), .A1 (sgo__sro_n800), .A2 (sgo__sro_n801));
BUF_X4 opt_ipo_c5746 (.Z (opt_ipo_n5162), .A (\A_imm_2s_complement[16] ));
BUF_X8 sgo__c814 (.Z (sgo__n836), .A (\A_imm_2s_complement[22] ));
BUF_X4 sgo__c1058 (.Z (sgo__n1009), .A (\A_imm_2s_complement[21] ));
NAND3_X2 sgo__sro_c776 (.ZN (sgo__sro_n809), .A1 (slo__sro_n1605), .A2 (sgo__sro_n811), .A3 (sgo__sro_n799));
BUF_X32 sgo__c1358 (.Z (A_in), .A (sgo__n1251));
INV_X8 opt_ipo_c5729 (.ZN (opt_ipo_n5145), .A (opt_ipo_n5664));
BUF_X2 spw__L1_c8576 (.Z (spw__n7777), .A (n_0_1_599));
INV_X1 sgo__sro_c904 (.ZN (sgo__sro_n909), .A (opt_ipo_n5278));
INV_X1 sgo__sro_c905 (.ZN (sgo__sro_n908), .A (\A_imm_2s_complement[15] ));
NAND2_X1 sgo__sro_c906 (.ZN (sgo__sro_n907), .A1 (opt_ipo_n5415), .A2 (n_0_1_687));
OAI21_X1 sgo__sro_c907 (.ZN (sgo__sro_n906), .A (sgo__sro_n907), .B1 (sgo__sro_n908), .B2 (sgo__sro_n909));
AOI21_X2 sgo__sro_c908 (.ZN (sgo__sro_n905), .A (sgo__sro_n906), .B1 (\A_imm_2s_complement[16] ), .B2 (opt_ipo_n5679));
BUF_X4 opt_ipo_c5749 (.Z (opt_ipo_n5165), .A (n_0_1_794));
CLKBUF_X2 sgo__c983 (.Z (sgo__n959), .A (slo__n3345));
BUF_X1 sgo__c986 (.Z (sgo__n962), .A (\A_imm[4] ));
AND2_X4 sgo__c973 (.ZN (sgo__sro_n811), .A1 (sgo__sro_n702), .A2 (n_0_1_76));
CLKBUF_X3 sgo__c1110 (.Z (sgo__n1043), .A (slo__xsl_n4322));
NAND2_X1 sgo__sro_c1283 (.ZN (sgo__sro_n1195), .A1 (opt_ipo_n5303), .A2 (opt_ipo_n5423));
CLKBUF_X1 CLOCK_slh__c7906 (.Z (CLOCK_slh__n7196), .A (CLOCK_slh__n7195));
BUF_X1 sgo__c1120 (.Z (sgo__n1053), .A (\A_imm[2] ));
BUF_X2 sgo__c1123 (.Z (sgo__n1056), .A (\A_imm_2s_complement[16] ));
OAI21_X1 sgo__sro_c1284 (.ZN (sgo__sro_n1194), .A (sgo__sro_n1195), .B1 (opt_ipo_n5374), .B2 (sgo__sro_n1197));
BUF_X32 opt_ipo_c6234 (.Z (opt_ipo_n5679), .A (n_0_1_688));
AOI21_X2 sgo__sro_c1285 (.ZN (n_0_1_544), .A (sgo__sro_n1194), .B1 (opt_ipo_n5785), .B2 (slo___n2464));
CLKBUF_X2 sgo__c1345 (.Z (sgo__n1238), .A (n_0_1_822));
BUF_X8 sgo__c1348 (.Z (sgo__n1241), .A (\A_imm_2s_complement[29] ));
INV_X1 sgo__sro_c1302 (.ZN (sgo__sro_n1210), .A (n_0_1_897));
INV_X1 sgo__sro_c1303 (.ZN (sgo__sro_n1209), .A (n_0_1_902));
NAND2_X1 sgo__sro_c1304 (.ZN (sgo__sro_n1208), .A1 (sgo__sro_n1210), .A2 (sgo__sro_n1209));
NOR3_X4 sgo__sro_c1305 (.ZN (n_0_1_894), .A1 (sgo__sro_n809), .A2 (sgo__sro_n719), .A3 (sgo__sro_n1208));
INV_X4 sgo__c1447 (.ZN (sgo__n1325), .A (sgo__n1324));
INV_X8 CLOCK_slo__mro_c7451 (.ZN (n_0_1_344), .A (CLOCK_slo__mro_n6730));
OR2_X1 sgo__sro_c1407 (.ZN (sgo__sro_n1290), .A1 (slo__xsl_n1669), .A2 (n_0_1_729));
NAND3_X1 sgo__sro_c1408 (.ZN (sgo__sro_n1289), .A1 (n_0_1_939), .A2 (n_0_1_940), .A3 (sgo__sro_n1290));
BUF_X4 sgo__c1324 (.Z (sgo__n1223), .A (n_0_1_767));
BUF_X1 spw__L1_c1_c8538 (.Z (\A_imm[6] ), .A (spw__n7741));
BUF_X8 sgo__c1463 (.Z (sgo__n1339), .A (\A_imm_2s_complement[25] ));
AND2_X4 sgo__sro_c1384 (.ZN (sgo__sro_n1270), .A1 (n_0_1_889), .A2 (n_0_1_892));
NAND3_X4 sgo__sro_c1385 (.ZN (n_0_1_888), .A1 (n_0_1_891), .A2 (n_0_1_890), .A3 (sgo__sro_n1270));
AOI222_X1 slo__sro_c2758 (.ZN (slo__sro_n2477), .A1 (opt_ipo_n5438), .A2 (\A_imm_2s_complement[8] )
    , .B1 (\A_imm_2s_complement[7] ), .B2 (opt_ipo_n5258), .C1 (opt_ipo_n5423), .C2 (slo__n1788));
NAND3_X2 sgo__sro_c1391 (.ZN (sgo__sro_n1273), .A1 (n_0_1_894), .A2 (n_0_1_882), .A3 (n_0_1_907));
NOR2_X4 sgo__sro_c1392 (.ZN (sgo__sro_n1272), .A1 (slo__sro_n1908), .A2 (sgo__sro_n1273));
INV_X4 opt_ipo_c6350 (.ZN (opt_ipo_n5795), .A (n_0_1_790));
INV_X4 opt_ipo_c6340 (.ZN (opt_ipo_n5785), .A (\A_imm_2s_complement[20] ));
INV_X1 slo__xsl_c1498 (.ZN (slo__xsl_n1367), .A (n_0_1_808));
INV_X2 slo__xsl_c1499 (.ZN (slo__xsl_n1366), .A (slo__xsl_n1367));
INV_X2 slo__c1508 (.ZN (slo__n1376), .A (n_0_1_767));
BUF_X2 slo__c1722 (.Z (slo__n1550), .A (\A_imm_2s_complement[24] ));
CLKBUF_X3 slo__c1620 (.Z (spd__n7595), .A (n_0_1_301));
CLKBUF_X2 slo__c1731 (.Z (slo__n1559), .A (n_0_1_800));
INV_X1 slo__xsl_c1564 (.ZN (slo__xsl_n1426), .A (n_0_1_810));
INV_X4 slo__xsl_c1565 (.ZN (slo__xsl_n1425), .A (slo__xsl_n1426));
OR2_X1 slo__sro_c1600 (.ZN (slo__sro_n1459), .A1 (slo__n1588), .A2 (n_0_1_609));
CLKBUF_X2 slo__c1541 (.Z (slo__n1402), .A (n_0_1_798));
OR2_X4 slo__sro_c1601 (.ZN (slo__sro_n1458), .A1 (opt_ipo_n5315), .A2 (slo__sro_n1459));
CLKBUF_X1 slo__c1641 (.Z (slo__n1493), .A (n_0_1_806));
INV_X1 slo__c1755 (.ZN (slo__n1581), .A (slo__n1580));
INV_X8 slo__c1756 (.ZN (n_0_1_600), .A (slo__n1581));
NOR2_X1 slo__sro_c1769 (.ZN (slo__sro_n1596), .A1 (n_0_1_600), .A2 (opt_ipo_n5165));
INV_X1 slo__sro_c1770 (.ZN (slo__sro_n1595), .A (slo__sro_n1596));
NAND2_X1 slo__sro_c1771 (.ZN (slo__sro_n1594), .A1 (slo__sro_n1595), .A2 (n_0_1_577));
INV_X1 slo__sro_c1802 (.ZN (slo__sro_n1623), .A (drc_ipo_n58));
INV_X1 slo__sro_c1786 (.ZN (slo__sro_n1608), .A (\aggregated_res[14][39] ));
INV_X1 slo__sro_c1787 (.ZN (slo__sro_n1607), .A (n_0_812));
NAND2_X1 slo__sro_c1788 (.ZN (slo__sro_n1606), .A1 (slo__sro_n1608), .A2 (slo__sro_n1607));
NOR2_X2 slo__sro_c1789 (.ZN (slo__sro_n1605), .A1 (\aggregated_res[14][45] ), .A2 (slo__sro_n1606));
NAND2_X1 slo__sro_c1804 (.ZN (slo__sro_n1621), .A1 (n_0_159), .A2 (slo__sro_n1623));
NAND2_X2 slo__sro_c1805 (.ZN (n_0_1_220), .A1 (slo__sro_n1622), .A2 (slo__sro_n1621));
INV_X1 slo__c1814 (.ZN (n_0_1_172), .A (slo__n1627));
INV_X1 slo__xsl_c1885 (.ZN (slo__xsl_n1695), .A (spw__n7686));
INV_X1 slo__xsl_c1832 (.ZN (slo__xsl_n1642), .A (n_0_1_818));
INV_X2 slo__xsl_c1833 (.ZN (slo__xsl_n1641), .A (slo__xsl_n1642));
INV_X2 slo__xsl_c1886 (.ZN (slo__xsl_n1694), .A (slo__xsl_n1695));
BUF_X2 slo__c1893 (.Z (slo__n1702), .A (\A_imm_2s_complement[12] ));
INV_X1 slo__xsl_c1860 (.ZN (slo__xsl_n1670), .A (n_0_1_830));
INV_X2 slo__xsl_c1861 (.ZN (slo__xsl_n1669), .A (slo__xsl_n1670));
INV_X1 slo__sro_c1943 (.ZN (slo__sro_n1749), .A (\A_imm[29] ));
INV_X1 slo__sro_c1944 (.ZN (slo__sro_n1748), .A (n_0_1_730));
NOR2_X1 slo__sro_c1945 (.ZN (slo__sro_n1747), .A1 (slo__sro_n1749), .A2 (slo__sro_n1748));
CLKBUF_X1 CLOCK_slh__c7871 (.Z (CLOCK_slh__n7168), .A (CLOCK_slh__n7160));
INV_X1 slo__xsl_c1933 (.ZN (slo__xsl_n1737), .A (n_0_1_832));
INV_X2 slo__xsl_c1934 (.ZN (slo__xsl_n1736), .A (slo__xsl_n1737));
AOI21_X1 slo__sro_c1946 (.ZN (slo__sro_n1746), .A (slo__sro_n1747), .B1 (\A_imm_2s_complement[30] ), .B2 (n_0_1_731));
CLKBUF_X2 slo__c2008 (.Z (slo__n1801), .A (\A_imm[3] ));
BUF_X2 slo__c1962 (.Z (slo__n1762), .A (n_0_1_473));
INV_X1 slo__xsl_c2112 (.ZN (slo__xsl_n1890), .A (opt_ipo_n5208));
INV_X2 slo__xsl_c2113 (.ZN (slo__xsl_n1889), .A (slo__xsl_n1890));
CLKBUF_X1 slo__c2019 (.Z (slo__n1812), .A (n_0_1_820));
CLKBUF_X2 slo__c2035 (.Z (slo__n1828), .A (slo__xsl_n4785));
CLKBUF_X1 slo__c2120 (.Z (slo__n1897), .A (opt_ipo_n5209));
NAND3_X2 slo__sro_c2130 (.ZN (slo__sro_n1908), .A1 (sgo__sro_n741), .A2 (sgo__sro_n739), .A3 (n_0_1_876));
NOR2_X1 slo__mro_c2073 (.ZN (slo__mro_n1861), .A1 (n_0_1_519), .A2 (slo__n2885));
BUF_X4 slo__mro_c2074 (.Z (slo__mro_n1860), .A (slo__mro_n1861));
BUF_X4 slo__c2162 (.Z (slo__n1936), .A (n_0_1_215));
INV_X1 slo__xsl_c2196 (.ZN (slo__xsl_n1964), .A (n_0_1_478));
INV_X4 slo__xsl_c2197 (.ZN (slo__xsl_n1963), .A (slo__xsl_n1964));
CLKBUF_X1 CLOCK_slh__c7918 (.Z (sph__n7808), .A (CLOCK_slh__n7207));
CLKBUF_X1 CLOCK_slh__c7917 (.Z (CLOCK_slh__n7207), .A (CLOCK_slh__n7206));
BUF_X8 opt_ipo_c6329 (.Z (opt_ipo_n5774), .A (n_0_1_558));
INV_X1 slo__xsl_c2249 (.ZN (slo__xsl_n2011), .A (sgo__n880));
INV_X2 slo__xsl_c2250 (.ZN (slo__xsl_n2010), .A (slo__xsl_n2011));
BUF_X8 slo__c2314 (.Z (slo__n2069), .A (n_0_1_127));
NAND2_X1 slo__mro_c2320 (.ZN (slo__mro_n2075), .A1 (n_0_1_127), .A2 (\A_imm_2s_complement[1] ));
NAND3_X1 slo__sro_c2325 (.ZN (slo__sro_n2079), .A1 (n_0_1_91), .A2 (slo__mro_n2075), .A3 (slo__sro_n2080));
CLKBUF_X1 CLOCK_slh__c7907 (.Z (CLOCK_slh__n7200), .A (CLOCK_slh__n7196));
BUF_X1 spw__L2_c8577 (.Z (spw__n7778), .A (spw__n7777));
INV_X1 opt_ipo_c5748 (.ZN (opt_ipo_n5164), .A (opt_ipo_n5165));
BUF_X8 spd__c8396 (.Z (slo__n1475), .A (spd__n7595));
OR2_X1 slo__sro_c2400 (.ZN (slo__sro_n2150), .A1 (n_0_1_394), .A2 (n_0_1_351));
NOR2_X4 slo__sro_c2401 (.ZN (slo__sro_n2149), .A1 (slo__n3799), .A2 (slo__sro_n2150));
CLKBUF_X2 slo__c2474 (.Z (slo__n2216), .A (\A_imm[24] ));
INV_X2 slo__c2491 (.ZN (slo__n2235), .A (n_0_1_767));
CLKBUF_X3 slo___L1_c2500 (.Z (slo___n2244), .A (n_0_1_472));
NOR2_X2 slo__c2488 (.ZN (slo__n2232), .A1 (sgo__sro_n1272), .A2 (n_0_1_908));
CLKBUF_X3 slo___L2_c2501 (.Z (slo___n2245), .A (slo___n2244));
NAND2_X1 CLOCK_slo__sro_c7459 (.ZN (CLOCK_slo__sro_n6735), .A1 (drc_ipo_n58), .A2 (n_0_49));
CLKBUF_X1 slo___L1_c2503 (.Z (slo___n2247), .A (n_0_1_472));
CLKBUF_X1 slo___L1_c2504 (.Z (slo___n2248), .A (n_0_1_472));
AOI222_X1 slo__sro_c2593 (.ZN (slo__sro_n2333), .A1 (n_0_1_687), .A2 (slo__n1801)
    , .B1 (opt_ipo_n5280), .B2 (\A_imm_2s_complement[3] ), .C1 (n_0_1_688), .C2 (\A_imm_2s_complement[4] ));
INV_X4 opt_ipo_c5775 (.ZN (opt_ipo_n5191), .A (slo__n3399));
INV_X1 slo__c2799 (.ZN (slo__n2517), .A (slo__n2400));
AOI222_X1 slo__sro_c2818 (.ZN (n_0_1_137), .A1 (n_0_1_168), .A2 (\A_imm_2s_complement[3] )
    , .B1 (n_0_1_170), .B2 (sgo__n1053), .C1 (n_0_1_167), .C2 (\A_imm_2s_complement[2] ));
INV_X4 slo__c2811 (.ZN (slo__n2528), .A (\aggregated_res[14][56] ));
XNOR2_X2 slo__c3181 (.ZN (slo__n2871), .A (n_0_1_522), .B (n_0_1_480));
NAND2_X4 slo__c2666 (.ZN (slo__n2400), .A1 (slo__n2232), .A2 (hfn_ipo_n46));
BUF_X4 slo__c3112 (.Z (slo__n2805), .A (\A_imm_2s_complement[4] ));
NAND2_X4 CLOCK_slo__sro_c7461 (.ZN (n_0_1_394), .A1 (CLOCK_slo__sro_n6735), .A2 (CLOCK_slo__sro_n6734));
CLKBUF_X1 CLOCK_slh__c7865 (.Z (CLOCK_slh__n7158), .A (enable));
CLKBUF_X1 slo__c3067 (.Z (slo__n2762), .A (n_0_1_828));
OR2_X2 slo__sro_c2861 (.ZN (slo__sro_n2570), .A1 (n_0_1_436), .A2 (n_0_1_435));
INV_X8 slo__sro_c2862 (.ZN (n_0_1_429), .A (slo__sro_n2570));
CLKBUF_X1 slo__c3225 (.Z (slo__n2915), .A (\A_imm[18] ));
CLKBUF_X1 CLOCK_slh__c7879 (.Z (CLOCK_slh__n7169), .A (CLOCK_slh__n7168));
CLKBUF_X1 CLOCK_slh__c7901 (.Z (CLOCK_slh__n7194), .A (CLOCK_slh__n7190));
BUF_X4 slo__c3278 (.Z (slo__n2969), .A (\A_imm_2s_complement[8] ));
AOI222_X1 slo__sro_c3295 (.ZN (slo__sro_n2992), .A1 (\A_imm_2s_complement[26] ), .A2 (slo___n2464)
    , .B1 (\A_imm_2s_complement[25] ), .B2 (opt_ipo_n5258), .C1 (opt_ipo_n5774), .C2 (opt_ipo_n5362));
BUF_X1 slo__c3195 (.Z (slo__n2885), .A (slo__n3640));
INV_X4 slo__c3336 (.ZN (slo__n3030), .A (slo__sro_n1458));
MUX2_X2 slo__sro_c3268 (.Z (slo__sro_n2959), .A (n_0_176), .B (n_0_40), .S (drc_ipo_n58));
CLKBUF_X1 CLOCK_slh__c7869 (.Z (CLOCK_slh__n7159), .A (CLOCK_slh__n7158));
BUF_X8 opt_ipo_c6265 (.Z (opt_ipo_n5710), .A (\A_imm_2s_complement[13] ));
INV_X2 opt_ipo_c6267 (.ZN (opt_ipo_n5712), .A (n_0_141));
BUF_X4 slo___L1_c3424 (.Z (slo___n3116), .A (n_0_1_387));
BUF_X2 spw__L1_c2_c8540 (.Z (spw__n7740), .A (spw__n7741));
CLKBUF_X1 slo__c3319 (.Z (slo__n3016), .A (\A_imm[1] ));
NAND3_X1 slo__sro_c3481 (.ZN (slo__sro_n3170), .A1 (n_0_1_838), .A2 (n_0_1_869), .A3 (n_0_1_870));
AOI222_X1 slo__sro_c3557 (.ZN (slo__sro_n3243), .A1 (\A_imm_2s_complement[28] ), .A2 (slo__n4931)
    , .B1 (\A_imm_2s_complement[27] ), .B2 (spw__n7778), .C1 (\A_imm[27] ), .C2 (opt_ipo_n5311));
AOI222_X1 slo__sro_c3636 (.ZN (slo__sro_n3317), .A1 (opt_ipo_n5151), .A2 (\A_imm_2s_complement[5] )
    , .B1 (slo__n3614), .B2 (\A_imm_2s_complement[4] ), .C1 (opt_ipo_n5312), .C2 (sgo__n962));
OR2_X4 slo__c3620 (.ZN (slo__n3307), .A1 (n_0_1_608), .A2 (n_0_1_607));
MUX2_X2 slo__c3445 (.Z (slo__n3134), .A (n_0_169), .B (n_0_47), .S (drc_ipo_n58));
MUX2_X2 slo__c3518 (.Z (slo__n3204), .A (n_0_165), .B (n_0_51), .S (drc_ipo_n58));
INV_X1 slo__sro_c3688 (.ZN (slo__sro_n3369), .A (slo__sro_n3370));
NOR2_X1 slo__sro_c3689 (.ZN (slo__sro_n3368), .A1 (n_0_1_968), .A2 (slo__sro_n3369));
CLKBUF_X1 CLOCK_slh__c7870 (.Z (CLOCK_slh__n7160), .A (CLOCK_slh__n7159));
AOI21_X4 slo__c3716 (.ZN (slo__n3399), .A (n_0_1_809), .B1 (n_0_16), .B2 (hfn_ipo_n41));
CLKBUF_X2 slo__c3719 (.Z (slo__n3402), .A (opt_ipo_n5191));
OR2_X1 slo__sro_c3723 (.ZN (slo__sro_n3407), .A1 (slo__n1812), .A2 (n_0_1_772));
NAND2_X1 slo__sro_c3724 (.ZN (slo__sro_n3406), .A1 (n_0_1_761), .A2 (slo__sro_n3407));
CLKBUF_X3 opt_ipo_c6219 (.Z (opt_ipo_n5664), .A (opt_ipo_n5146));
NAND2_X1 CLOCK_slo__sro_c7460 (.ZN (CLOCK_slo__sro_n6734), .A1 (n_0_167), .A2 (CLOCK_slo__sro_n6736));
INV_X1 CLOCK_slo__sro_c7458 (.ZN (CLOCK_slo__sro_n6736), .A (drc_ipo_n58));
CLKBUF_X1 slo___L1_c3784 (.Z (slo___n3458), .A (n_0_1_796));
INV_X1 opt_ipo_c6266 (.ZN (opt_ipo_n5711), .A (opt_ipo_n5712));
BUF_X4 slo___L1_c3815 (.Z (slo___n3489), .A (n_0_1_566));
BUF_X4 opt_ipo_c6241 (.Z (opt_ipo_n5686), .A (n_0_1_429));
BUF_X4 opt_ipo_c5687 (.Z (opt_ipo_n5103), .A (n_0_1_165));
INV_X2 opt_ipo_c5691 (.ZN (opt_ipo_n5107), .A (opt_ipo_n5108));
INV_X2 opt_ipo_c5692 (.ZN (opt_ipo_n5108), .A (n_0_1_220));
CLKBUF_X1 CTS_L1_c_tid1_6457 (.Z (CTS_n_tid1_5915), .A (clk));
CLKBUF_X1 slo___L1_c3822 (.Z (slo___n3496), .A (n_0_1_566));
BUF_X8 CLOCK_sgo__c7115 (.Z (CLOCK_sgo__n6468), .A (n_0_1_214));
CLKBUF_X2 slo__c3879 (.Z (slo__n3547), .A (\A_imm[16] ));
INV_X2 slo__c3945 (.ZN (slo__n3614), .A (slo__sro_n1458));
XNOR2_X1 slo__c3848 (.ZN (slo__n3522), .A (n_0_1_565), .B (n_0_1_521));
BUF_X2 slo__c3948 (.Z (slo__n3617), .A (\A_imm_2s_complement[7] ));
MUX2_X1 slo__c3930 (.Z (slo__n3595), .A (n_0_176), .B (n_0_40), .S (drc_ipo_n58));
XNOR2_X2 slo__c4031 (.ZN (slo__n3691), .A (slo__sro_n2959), .B (opt_ipo_n5315));
OR2_X2 slo__sro_c3918 (.ZN (slo__sro_n3584), .A1 (n_0_1_565), .A2 (n_0_1_607));
NOR2_X4 slo__sro_c3919 (.ZN (slo__n4197), .A1 (slo__n3595), .A2 (slo__sro_n3584));
INV_X4 opt_ipo_c5779 (.ZN (opt_ipo_n5195), .A (opt_ipo_n5196));
MUX2_X2 slo__c3974 (.Z (slo__n3640), .A (n_0_173), .B (n_0_43), .S (drc_ipo_n58));
BUF_X4 opt_ipo_c5743 (.Z (opt_ipo_n5159), .A (n_0_1_386));
NAND2_X1 slo__sro_c4025 (.ZN (slo__sro_n3685), .A1 (slo__n3204), .A2 (n_0_1_308));
INV_X1 opt_ipo_c6257 (.ZN (opt_ipo_n5702), .A (opt_ipo_n5703));
BUF_X4 opt_ipo_c6274 (.Z (opt_ipo_n5719), .A (n_0_1_384));
BUF_X8 opt_ipo_c5709 (.Z (opt_ipo_n5125), .A (n_0_1_255));
NAND2_X2 slo__sro_c4157 (.ZN (slo__sro_n3808), .A1 (slo__n2871), .A2 (slo__xsl_n1963));
INV_X4 slo__sro_c4158 (.ZN (n_0_1_473), .A (slo__sro_n3808));
INV_X1 slo__sro_c4076 (.ZN (slo__sro_n3736), .A (n_0_1_868));
INV_X1 slo__sro_c4077 (.ZN (slo__sro_n3735), .A (drc_ipo_n58));
NAND2_X1 slo__sro_c4078 (.ZN (slo__sro_n3734), .A1 (slo__sro_n3736), .A2 (slo__sro_n3735));
NAND2_X1 slo__sro_c4079 (.ZN (n_0_1_174), .A1 (n_0_1_177), .A2 (slo__sro_n3734));
BUF_X4 CLOCK_sgo__c7050 (.Z (CLOCK_sgo__n6410), .A (n_0_1_168));
INV_X1 slo__c4148 (.ZN (slo__n3799), .A (slo__n3204));
BUF_X4 slo__c4275 (.Z (slo__n3910), .A (\A_imm_2s_complement[5] ));
AND2_X2 slo__c4209 (.ZN (n_0_1_920), .A1 (slo__n3840), .A2 (opt_ipo_n5314));
CLKBUF_X1 CLOCK_spw__L1_c8100 (.Z (CLOCK_spw__n7299), .A (n_0_1_782));
XNOR2_X1 slo__c4196 (.ZN (slo__n3840), .A (n_0_1_651), .B (n_0_1_609));
INV_X1 slo__xsl_c4262 (.ZN (slo__xsl_n3901), .A (sgo__n1116));
INV_X4 slo__xsl_c4263 (.ZN (slo__xsl_n3900), .A (slo__xsl_n3901));
NAND2_X2 slo__sro_c4555 (.ZN (slo__sro_n4175), .A1 (n_0_39), .A2 (drc_ipo_n58));
NAND2_X1 slo__sro_c4556 (.ZN (slo__sro_n4174), .A1 (n_0_177), .A2 (slo__sro_n4176));
NAND2_X4 slo__sro_c4557 (.ZN (n_0_1_607), .A1 (slo__sro_n4175), .A2 (slo__sro_n4174));
INV_X1 slo__xsl_c4616 (.ZN (slo__xsl_n4224), .A (n_0_1_306));
INV_X4 slo__xsl_c4617 (.ZN (slo__xsl_n4223), .A (slo__xsl_n4224));
INV_X1 slo__xsl_c4740 (.ZN (slo__xsl_n4323), .A (n_0_1_778));
INV_X1 slo__xsl_c4741 (.ZN (slo__xsl_n4322), .A (slo__xsl_n4323));
CLKBUF_X1 spw__L1_c8485 (.Z (spw__n7686), .A (n_0_1_786));
BUF_X2 CLOCK_spw__L1_c8130 (.Z (CLOCK_spw__n7329), .A (drc_ipo_n52));
BUF_X1 CLOCK_spw__L2_c8123 (.Z (CLOCK_spw__n7322), .A (CLOCK_spw__n7320));
BUF_X4 opt_ipo_c5736 (.Z (opt_ipo_n5152), .A (slo__n1588));
INV_X1 slo__xsl_c5348 (.ZN (slo__xsl_n4786), .A (opt_ipo_n5416));
INV_X1 slo__xsl_c4945 (.ZN (slo__xsl_n4488), .A (CLOCK_spw__n7303));
INV_X2 slo__xsl_c4946 (.ZN (slo__xsl_n4487), .A (slo__xsl_n4488));
INV_X1 slo__xsl_c5349 (.ZN (slo__xsl_n4785), .A (slo__xsl_n4786));
BUF_X2 opt_ipo_c5781 (.Z (opt_ipo_n5197), .A (opt_ipo_n5198));
BUF_X16 slo__c5421 (.Z (sgo__n734), .A (slo__n4849));
INV_X4 opt_ipo_c5782 (.ZN (opt_ipo_n5198), .A (\A_imm_2s_complement[9] ));
CLKBUF_X1 sph__c8609 (.Z (CLOCK_slh_n7157), .A (sph__n7810));
INV_X4 CLOCK_opt_ipo_c6423 (.ZN (CLOCK_opt_ipo_n5880), .A (\A_imm_2s_complement[17] ));
CLKBUF_X2 opt_ipo_c5788 (.Z (opt_ipo_n5204), .A (opt_ipo_n5205));
INV_X8 opt_ipo_c5789 (.ZN (opt_ipo_n5205), .A (\A_imm_2s_complement[6] ));
BUF_X8 CLOCK_spw__L1_c8145 (.Z (CLOCK_spw__n7344), .A (n_0_1_645));
INV_X1 opt_ipo_c5792 (.ZN (opt_ipo_n5208), .A (opt_ipo_n5209));
INV_X1 opt_ipo_c5793 (.ZN (opt_ipo_n5209), .A (n_0_1_826));
CLKBUF_X1 CLOCK_slh__c7891 (.Z (CLOCK_slh__n7188), .A (CLOCK_slh__n7180));
INV_X2 opt_ipo_c5807 (.ZN (opt_ipo_n5223), .A (n_0_45));
BUF_X8 opt_ipo_c5808 (.Z (opt_ipo_n5224), .A (n_0_1_300));
BUF_X4 opt_ipo_c5814 (.Z (opt_ipo_n5230), .A (n_0_1_213));
CLKBUF_X1 CLOCK_spw__L1_c8104 (.Z (CLOCK_spw__n7303), .A (sgo__n681));
BUF_X4 opt_ipo_c5820 (.Z (Res[63]), .A (opt_ipo_n5239));
BUF_X8 opt_ipo_c5839 (.Z (opt_ipo_n5258), .A (slo__n4197));
BUF_X8 opt_ipo_c5859 (.Z (opt_ipo_n5278), .A (opt_ipo_n5280));
INV_X4 opt_ipo_c5861 (.ZN (opt_ipo_n5280), .A (n_0_1_930));
BUF_X8 opt_ipo_c5866 (.Z (opt_ipo_n5285), .A (slo__n1762));
BUF_X2 CLOCK_spw__L1_c8121 (.Z (CLOCK_spw__n7320), .A (n_0_1_385));
NAND2_X1 CLOCK_slo__sro_c7470 (.ZN (CLOCK_slo__sro_n6741), .A1 (CLOCK_slo__sro_n6742), .A2 (CLOCK_slo__sro_n6743));
CLKBUF_X1 CLOCK_slh__c7881 (.Z (CLOCK_slh__n7178), .A (CLOCK_slh__n7170));
INV_X4 opt_ipo_c5878 (.ZN (opt_ipo_n5297), .A (n_0_1_796));
CLKBUF_X1 CLOCK_slh__c7899 (.Z (CLOCK_slh__n7189), .A (CLOCK_slh__n7188));
BUF_X1 CLOCK_spw__L1_c8092 (.Z (CLOCK_spw__n7291), .A (slo__n3617));
INV_X4 opt_ipo_c5884 (.ZN (opt_ipo_n5303), .A (opt_ipo_n5307));
BUF_X4 opt_ipo_c5888 (.Z (opt_ipo_n5307), .A (n_0_1_812));
CLKBUF_X3 opt_ipo_c5892 (.Z (opt_ipo_n5311), .A (opt_ipo_n5312));
INV_X8 opt_ipo_c5893 (.ZN (opt_ipo_n5312), .A (slo__n3307));
INV_X1 opt_ipo_c5895 (.ZN (opt_ipo_n5314), .A (opt_ipo_n5315));
INV_X4 opt_ipo_c5896 (.ZN (opt_ipo_n5315), .A (n_0_1_607));
BUF_X4 CLOCK_spw__L2_c8122 (.Z (CLOCK_spw__n7321), .A (CLOCK_spw__n7320));
BUF_X4 opt_ipo_c5913 (.Z (opt_ipo_n5332), .A (slo__sro_n2149));
BUF_X8 opt_ipo_c5920 (.Z (opt_ipo_n5339), .A (opt_ipo_n5785));
BUF_X2 opt_ipo_c5939 (.Z (opt_ipo_n5358), .A (sgo__n844));
INV_X2 opt_ipo_c5943 (.ZN (opt_ipo_n5362), .A (sgo__n880));
BUF_X4 CLOCK_spw__L1_c8093 (.Z (CLOCK_spw__n7292), .A (slo__n3617));
INV_X8 opt_ipo_c5954 (.ZN (opt_ipo_n5373), .A (opt_ipo_n5374));
INV_X8 opt_ipo_c5955 (.ZN (opt_ipo_n5374), .A (\A_imm_2s_complement[19] ));
BUF_X8 opt_ipo_c5966 (.Z (opt_ipo_n5385), .A (n_0_1_170));
BUF_X8 opt_ipo_c5974 (.Z (opt_ipo_n5393), .A (n_0_1_642));
BUF_X16 opt_ipo_c5976 (.Z (opt_ipo_n5395), .A (n_0_1_644));
BUF_X1 opt_ipo_c5979 (.Z (opt_ipo_n5398), .A (n_0_1_650));
BUF_X8 opt_ipo_c5992 (.Z (opt_ipo_n5411), .A (CLOCK_opt_ipo_n5880));
INV_X4 opt_ipo_c5996 (.ZN (opt_ipo_n5415), .A (opt_ipo_n5416));
INV_X1 opt_ipo_c5997 (.ZN (opt_ipo_n5416), .A (opt_ipo_n5417));
INV_X2 opt_ipo_c5998 (.ZN (opt_ipo_n5417), .A (n_0_1_804));
BUF_X8 opt_ipo_c6000 (.Z (opt_ipo_n5419), .A (drc_ipo_n54));
BUF_X4 opt_ipo_c6004 (.Z (opt_ipo_n5423), .A (n_0_1_558));
BUF_X8 opt_ipo_c6014 (.Z (opt_ipo_n5433), .A (drc_ipo_n50));
BUF_X4 opt_ipo_c6019 (.Z (opt_ipo_n5438), .A (n_0_1_559));
CLKBUF_X1 CLOCK_slh__c7889 (.Z (CLOCK_slh__n7179), .A (CLOCK_slh__n7178));
CLKBUF_X3 opt_ipo_c6040 (.Z (opt_ipo_n5459), .A (slo__n3016));
CLKBUF_X3 opt_ipo_c6046 (.Z (opt_ipo_n5465), .A (opt_ipo_n5466));
INV_X8 opt_ipo_c6047 (.ZN (opt_ipo_n5466), .A (\A_imm_2s_complement[10] ));
INV_X2 opt_ipo_c6085 (.ZN (OVF), .A (opt_ipo_n5506));

endmodule //boothAlgoR4


