
// 	Thu Dec 22 19:36:37 2022
//	vlsi
//	192.168.126.129

module datapath__0_3 (opt_ipoPP_2, opt_ipoPP_6, opt_ipoPP_7, Res_imm, p_0);

output [63:0] p_0;
input [63:0] Res_imm;
input opt_ipoPP_2;
input opt_ipoPP_6;
input opt_ipoPP_7;
wire n_80;
wire n_66;
wire n_79;
wire n_63;
wire n_64;
wire n_5;
wire n_48;
wire n_3;
wire n_4;
wire n_41;
wire n_2;
wire n_94;
wire n_92;
wire n_95;
wire n_93;
wire n_103;
wire n_101;
wire n_105;
wire n_104;
wire n_113;
wire n_109;
wire n_120;
wire n_114;
wire n_128;
wire n_123;
wire n_135;
wire n_98;
wire n_137;
wire n_89;
wire n_90;
wire n_87;
wire n_88;
wire n_85;
wire n_83;
wire n_84;
wire n_23;
wire n_82;
wire n_21;
wire n_22;
wire n_19;
wire n_20;
wire n_31;
wire n_18;
wire n_29;
wire n_30;
wire n_27;
wire n_28;
wire n_78;
wire n_24;
wire n_25;
wire n_37;
wire n_77;
wire n_33;
wire n_76;
wire n_32;
wire n_74;
wire n_75;
wire n_70;
wire n_71;
wire n_68;
wire n_69;
wire n_43;
wire n_45;
wire n_49;
wire n_131;
wire n_61;
wire n_46;
wire n_26;
wire n_145;
wire n_42;
wire n_194;
wire n_60;
wire n_52;
wire n_171;
wire n_116;
wire n_50;
wire n_51;
wire n_55;
wire n_57;
wire n_53;
wire n_54;
wire n_56;
wire n_58;
wire n_65;
wire n_59;
wire n_144;
wire n_62;
wire n_204;
wire n_200;
wire n_184;
wire sgo__sro_n49;
wire sgo__sro_n31;
wire n_147;
wire n_142;
wire n_164;
wire n_150;
wire n_156;
wire n_151;
wire n_157;
wire n_159;
wire sgo__n77;
wire n_165;
wire n_155;
wire n_149;
wire n_160;
wire n_161;
wire n_158;
wire n_154;
wire n_162;
wire n_167;
wire n_163;
wire n_185;
wire n_13;
wire n_207;
wire n_205;
wire n_168;
wire n_202;
wire n_177;
wire n_175;
wire n_176;
wire n_181;
wire n_179;
wire n_180;
wire n_201;
wire n_182;
wire n_199;
wire n_209;
wire n_211;
wire n_210;
wire n_47;
wire n_146;
wire n_73;
wire n_36;
wire n_44;
wire n_140;
wire n_172;
wire n_72;
wire n_186;
wire n_190;
wire n_170;
wire n_215;
wire n_214;
wire n_148;
wire n_192;
wire n_174;
wire n_16;
wire n_198;
wire n_218;
wire n_15;
wire n_1;
wire n_14;
wire n_6;
wire n_7;
wire n_195;
wire n_212;
wire n_8;
wire n_9;
wire n_10;
wire n_17;
wire n_188;
wire n_11;
wire n_12;
wire n_216;
wire n_187;
wire n_39;
wire n_40;
wire n_96;
wire n_97;
wire n_99;
wire n_100;
wire n_102;
wire n_106;
wire n_107;
wire n_108;
wire n_112;
wire n_110;
wire n_111;
wire n_115;
wire n_117;
wire n_118;
wire n_119;
wire n_121;
wire n_122;
wire n_125;
wire n_124;
wire n_126;
wire n_127;
wire n_129;
wire n_133;
wire n_134;
wire n_136;
wire n_138;
wire n_139;
wire sgo__sro_n50;
wire n_153;
wire n_166;
wire n_189;
wire n_197;
wire sgo__sro_n32;
wire n_193;
wire n_203;
wire n_206;
wire n_213;


INV_X2 sgo__sro_c38 (.ZN (sgo__sro_n31), .A (sgo__sro_n32));
OR4_X2 i_272 (.ZN (n_216), .A1 (Res_imm[25]), .A2 (Res_imm[24]), .A3 (Res_imm[27]), .A4 (Res_imm[26]));
INV_X1 i_271 (.ZN (n_215), .A (Res_imm[39]));
INV_X1 i_270 (.ZN (n_214), .A (Res_imm[38]));
INV_X1 i_269 (.ZN (n_213), .A (n_193));
NAND2_X1 i_268 (.ZN (n_212), .A1 (n_197), .A2 (n_42));
NOR4_X1 i_267 (.ZN (n_211), .A1 (n_213), .A2 (n_212), .A3 (Res_imm[39]), .A4 (Res_imm[38]));
AND2_X1 i_266 (.ZN (n_210), .A1 (n_190), .A2 (n_186));
NOR3_X2 i_265 (.ZN (n_207), .A1 (Res_imm[46]), .A2 (Res_imm[44]), .A3 (Res_imm[45]));
INV_X1 i_264 (.ZN (n_206), .A (Res_imm[58]));
NAND3_X1 i_263 (.ZN (n_205), .A1 (n_154), .A2 (n_153), .A3 (n_206));
NOR4_X4 i_262 (.ZN (n_204), .A1 (Res_imm[51]), .A2 (Res_imm[50]), .A3 (Res_imm[49]), .A4 (Res_imm[48]));
NOR3_X1 i_261 (.ZN (n_203), .A1 (Res_imm[59]), .A2 (n_205), .A3 (Res_imm[47]));
AND3_X2 i_260 (.ZN (n_202), .A1 (n_160), .A2 (n_203), .A3 (n_204));
INV_X1 i_259 (.ZN (n_201), .A (Res_imm[62]));
NOR2_X1 i_258 (.ZN (n_200), .A1 (Res_imm[61]), .A2 (Res_imm[60]));
AND2_X1 i_257 (.ZN (n_199), .A1 (n_201), .A2 (n_200));
INV_X1 i_256 (.ZN (n_198), .A (Res_imm[32]));
INV_X1 i_255 (.ZN (n_197), .A (Res_imm[31]));
INV_X1 i_253 (.ZN (n_195), .A (Res_imm[29]));
INV_X1 i_252 (.ZN (n_194), .A (Res_imm[28]));
NOR2_X1 i_251 (.ZN (n_193), .A1 (Res_imm[29]), .A2 (Res_imm[28]));
NAND3_X1 i_250 (.ZN (n_192), .A1 (n_197), .A2 (n_42), .A3 (n_193));
NOR3_X4 i_248 (.ZN (n_190), .A1 (Res_imm[35]), .A2 (Res_imm[33]), .A3 (Res_imm[34]));
INV_X1 i_247 (.ZN (n_189), .A (n_190));
NOR3_X2 i_246 (.ZN (n_188), .A1 (Res_imm[39]), .A2 (Res_imm[38]), .A3 (n_189));
OR2_X1 i_245 (.ZN (n_187), .A1 (Res_imm[36]), .A2 (Res_imm[32]));
NOR2_X1 i_244 (.ZN (n_186), .A1 (Res_imm[37]), .A2 (n_187));
AND3_X1 i_243 (.ZN (n_185), .A1 (n_148), .A2 (n_188), .A3 (n_186));
INV_X1 i_242 (.ZN (n_184), .A (Res_imm[42]));
INV_X1 sgo__sro_c63 (.ZN (sgo__sro_n49), .A (sgo__sro_n50));
AOI21_X1 sgo__sro_c64 (.ZN (p_0[53]), .A (sgo__sro_n49), .B1 (n_65), .B2 (n_144));
NOR4_X4 i_239 (.ZN (n_171), .A1 (Res_imm[43]), .A2 (Res_imm[42]), .A3 (Res_imm[41]), .A4 (Res_imm[40]));
INV_X1 i_238 (.ZN (n_166), .A (n_171));
NOR2_X2 i_237 (.ZN (n_165), .A1 (Res_imm[47]), .A2 (n_166));
NOR3_X1 i_236 (.ZN (n_164), .A1 (Res_imm[54]), .A2 (opt_ipoPP_7), .A3 (Res_imm[53]));
NOR4_X4 i_235 (.ZN (n_160), .A1 (Res_imm[54]), .A2 (Res_imm[53]), .A3 (Res_imm[52]), .A4 (Res_imm[55]));
AND2_X1 i_234 (.ZN (n_159), .A1 (n_153), .A2 (n_160));
INV_X1 i_233 (.ZN (n_154), .A (Res_imm[57]));
INV_X1 i_232 (.ZN (n_153), .A (Res_imm[56]));
NOR2_X1 i_231 (.ZN (n_149), .A1 (opt_ipoPP_6), .A2 (Res_imm[56]));
NOR2_X1 i_230 (.ZN (n_144), .A1 (Res_imm[53]), .A2 (opt_ipoPP_7));
NAND3_X2 sgo__sro_c37 (.ZN (sgo__sro_n32), .A1 (n_185), .A2 (n_13), .A3 (n_207));
INV_X1 i_226 (.ZN (n_139), .A (n_135));
NOR3_X1 i_225 (.ZN (n_138), .A1 (Res_imm[25]), .A2 (n_139), .A3 (Res_imm[26]));
INV_X1 i_224 (.ZN (n_137), .A (n_138));
AOI21_X1 i_223 (.ZN (p_0[26]), .A (n_138), .B1 (Res_imm[26]), .B2 (n_134));
INV_X1 i_222 (.ZN (n_136), .A (Res_imm[25]));
NOR2_X1 i_221 (.ZN (n_135), .A1 (n_98), .A2 (Res_imm[24]));
NAND2_X1 i_220 (.ZN (n_134), .A1 (n_136), .A2 (n_135));
OAI21_X1 i_219 (.ZN (n_133), .A (n_134), .B1 (n_136), .B2 (n_135));
INV_X1 i_218 (.ZN (p_0[25]), .A (n_133));
NAND2_X2 sgo__sro_c39 (.ZN (n_163), .A1 (n_165), .A2 (sgo__sro_n31));
NOR4_X4 i_216 (.ZN (n_131), .A1 (Res_imm[23]), .A2 (Res_imm[22]), .A3 (Res_imm[21]), .A4 (n_123));
AOI21_X1 i_214 (.ZN (p_0[23]), .A (n_131), .B1 (Res_imm[23]), .B2 (n_127));
INV_X1 i_213 (.ZN (n_129), .A (Res_imm[22]));
NOR2_X1 i_212 (.ZN (n_128), .A1 (n_123), .A2 (Res_imm[21]));
NAND2_X1 i_211 (.ZN (n_127), .A1 (n_129), .A2 (n_128));
OAI21_X1 i_210 (.ZN (n_126), .A (n_127), .B1 (n_129), .B2 (n_128));
INV_X1 i_209 (.ZN (p_0[22]), .A (n_126));
INV_X1 i_208 (.ZN (n_125), .A (Res_imm[20]));
INV_X1 i_207 (.ZN (n_124), .A (Res_imm[18]));
NAND4_X4 i_206 (.ZN (n_123), .A1 (n_125), .A2 (n_115), .A3 (n_121), .A4 (n_124));
OAI21_X1 i_205 (.ZN (n_122), .A (n_123), .B1 (n_125), .B2 (n_118));
INV_X1 i_204 (.ZN (p_0[20]), .A (n_122));
INV_X1 i_203 (.ZN (n_121), .A (Res_imm[19]));
NOR2_X1 i_202 (.ZN (n_120), .A1 (n_114), .A2 (Res_imm[18]));
INV_X1 i_201 (.ZN (n_119), .A (n_120));
NOR2_X1 i_200 (.ZN (n_118), .A1 (Res_imm[19]), .A2 (n_119));
AOI21_X1 i_199 (.ZN (p_0[19]), .A (n_118), .B1 (Res_imm[19]), .B2 (n_119));
INV_X1 i_198 (.ZN (n_117), .A (Res_imm[16]));
NAND3_X2 i_197 (.ZN (n_116), .A1 (n_112), .A2 (n_110), .A3 (n_117));
NOR2_X2 i_196 (.ZN (n_115), .A1 (Res_imm[17]), .A2 (n_116));
INV_X1 i_195 (.ZN (n_114), .A (n_115));
AOI21_X1 i_194 (.ZN (p_0[17]), .A (n_115), .B1 (Res_imm[17]), .B2 (n_116));
INV_X1 i_193 (.ZN (n_112), .A (n_108));
INV_X1 i_192 (.ZN (n_111), .A (n_107));
NOR2_X1 i_191 (.ZN (n_110), .A1 (Res_imm[15]), .A2 (n_101));
NAND2_X1 i_190 (.ZN (n_109), .A1 (n_112), .A2 (n_110));
AOI22_X1 i_189 (.ZN (p_0[15]), .A1 (n_112), .A2 (n_110), .B1 (Res_imm[15]), .B2 (n_111));
OR3_X1 i_188 (.ZN (n_108), .A1 (Res_imm[14]), .A2 (Res_imm[12]), .A3 (Res_imm[13]));
AOI21_X1 i_187 (.ZN (p_0[14]), .A (n_107), .B1 (Res_imm[14]), .B2 (n_106));
NOR2_X1 i_186 (.ZN (n_107), .A1 (n_106), .A2 (Res_imm[14]));
INV_X1 i_185 (.ZN (n_106), .A (n_105));
NOR2_X1 i_184 (.ZN (n_105), .A1 (n_104), .A2 (Res_imm[13]));
INV_X1 i_183 (.ZN (n_104), .A (n_103));
NOR2_X1 i_182 (.ZN (n_103), .A1 (n_101), .A2 (Res_imm[12]));
INV_X1 i_181 (.ZN (n_102), .A (Res_imm[11]));
NAND3_X1 i_180 (.ZN (n_101), .A1 (n_39), .A2 (n_99), .A3 (n_102));
OAI21_X1 i_179 (.ZN (n_100), .A (n_101), .B1 (n_102), .B2 (n_97));
INV_X1 i_178 (.ZN (p_0[11]), .A (n_100));
NOR3_X1 i_177 (.ZN (n_99), .A1 (Res_imm[10]), .A2 (Res_imm[8]), .A3 (Res_imm[9]));
AOI21_X1 i_176 (.ZN (p_0[10]), .A (n_97), .B1 (Res_imm[10]), .B2 (n_96));
NOR2_X1 i_175 (.ZN (n_97), .A1 (n_96), .A2 (Res_imm[10]));
INV_X1 i_174 (.ZN (n_96), .A (n_95));
NOR2_X1 i_173 (.ZN (n_95), .A1 (n_93), .A2 (Res_imm[9]));
INV_X1 i_172 (.ZN (n_94), .A (n_93));
OR2_X1 i_171 (.ZN (n_93), .A1 (n_92), .A2 (Res_imm[8]));
INV_X1 i_170 (.ZN (n_92), .A (n_39));
NOR2_X1 i_169 (.ZN (n_80), .A1 (Res_imm[1]), .A2 (Res_imm[0]));
INV_X1 i_168 (.ZN (n_79), .A (n_80));
NOR2_X1 i_167 (.ZN (n_66), .A1 (Res_imm[2]), .A2 (n_79));
INV_X1 i_166 (.ZN (n_64), .A (n_66));
NOR2_X1 i_165 (.ZN (n_63), .A1 (Res_imm[3]), .A2 (n_64));
INV_X1 i_164 (.ZN (n_48), .A (n_63));
NOR4_X1 i_163 (.ZN (n_41), .A1 (Res_imm[6]), .A2 (Res_imm[5]), .A3 (Res_imm[4]), .A4 (n_48));
INV_X1 i_162 (.ZN (n_40), .A (n_41));
NOR2_X1 i_161 (.ZN (n_39), .A1 (Res_imm[7]), .A2 (n_40));
AOI21_X1 i_160 (.ZN (p_0[7]), .A (n_39), .B1 (Res_imm[7]), .B2 (n_40));
INV_X1 i_335 (.ZN (n_17), .A (Res_imm[45]));
INV_X1 i_334 (.ZN (n_16), .A (Res_imm[44]));
INV_X1 i_159 (.ZN (n_15), .A (Res_imm[37]));
INV_X1 i_158 (.ZN (n_14), .A (n_187));
NAND3_X1 i_156 (.ZN (n_12), .A1 (n_15), .A2 (n_14), .A3 (n_13));
INV_X1 i_155 (.ZN (n_11), .A (n_12));
NAND3_X2 i_154 (.ZN (n_77), .A1 (n_148), .A2 (n_188), .A3 (n_11));
INV_X32 sgo__c104 (.ZN (n_13), .A (sgo__n77));
NAND4_X1 i_303 (.ZN (n_71), .A1 (n_78), .A2 (n_17), .A3 (n_16), .A4 (n_171));
NAND2_X1 i_302 (.ZN (n_10), .A1 (n_171), .A2 (n_16));
OAI21_X1 i_301 (.ZN (n_9), .A (Res_imm[45]), .B1 (n_10), .B2 (n_77));
NAND2_X1 i_300 (.ZN (n_8), .A1 (n_9), .A2 (n_71));
INV_X1 i_297 (.ZN (p_0[45]), .A (n_8));
INV_X1 i_153 (.ZN (n_142), .A (n_212));
NAND3_X4 i_152 (.ZN (n_7), .A1 (n_13), .A2 (n_194), .A3 (n_195));
INV_X4 i_151 (.ZN (n_87), .A (n_7));
NAND2_X1 i_150 (.ZN (n_6), .A1 (n_87), .A2 (n_142));
INV_X1 i_149 (.ZN (n_1), .A (n_6));
NAND3_X1 i_148 (.ZN (n_28), .A1 (n_1), .A2 (n_190), .A3 (n_14));
INV_X1 i_147 (.ZN (n_29), .A (n_28));
NAND2_X1 i_146 (.ZN (n_147), .A1 (n_29), .A2 (n_15));
XNOR2_X1 i_145 (.ZN (n_218), .A (n_147), .B (Res_imm[38]));
INV_X1 i_131 (.ZN (p_0[38]), .A (n_218));
NAND4_X1 i_130 (.ZN (n_30), .A1 (n_190), .A2 (n_198), .A3 (n_142), .A4 (n_87));
INV_X1 i_129 (.ZN (n_31), .A (n_30));
NAND3_X1 i_229 (.ZN (n_174), .A1 (n_78), .A2 (n_16), .A3 (n_171));
INV_X1 i_228 (.ZN (n_74), .A (n_174));
INV_X1 i_127 (.ZN (n_172), .A (opt_ipoPP_2));
INV_X1 i_126 (.ZN (n_170), .A (Res_imm[40]));
INV_X1 i_125 (.ZN (n_148), .A (n_192));
NAND4_X1 i_124 (.ZN (n_146), .A1 (n_170), .A2 (n_215), .A3 (n_214), .A4 (n_148));
INV_X1 i_123 (.ZN (n_140), .A (n_146));
NAND3_X1 i_122 (.ZN (n_73), .A1 (n_186), .A2 (n_13), .A3 (n_190));
INV_X1 i_121 (.ZN (n_72), .A (n_73));
NAND3_X1 i_120 (.ZN (n_47), .A1 (n_140), .A2 (n_172), .A3 (n_72));
OAI21_X1 i_119 (.ZN (n_44), .A (opt_ipoPP_2), .B1 (n_146), .B2 (n_73));
NAND2_X1 i_118 (.ZN (n_36), .A1 (n_44), .A2 (n_47));
INV_X1 i_117 (.ZN (p_0[41]), .A (n_36));
NOR2_X1 i_116 (.ZN (n_37), .A1 (n_146), .A2 (n_73));
AND4_X2 sgo__c80 (.ZN (n_209), .A1 (n_210), .A2 (n_13), .A3 (n_211), .A4 (n_207));
OR2_X4 sgo__c102 (.ZN (sgo__n77), .A1 (n_216), .A2 (n_98));
NAND4_X1 i_108 (.ZN (n_182), .A1 (n_209), .A2 (n_171), .A3 (n_202), .A4 (n_199));
INV_X1 i_107 (.ZN (n_181), .A (n_182));
NAND2_X1 i_106 (.ZN (n_180), .A1 (n_201), .A2 (Res_imm[63]));
NAND4_X1 i_105 (.ZN (n_179), .A1 (n_209), .A2 (n_200), .A3 (n_202), .A4 (n_171));
OAI22_X1 i_104 (.ZN (p_0[63]), .A1 (n_179), .A2 (n_180), .B1 (n_181), .B2 (Res_imm[63]));
AOI21_X1 i_103 (.ZN (p_0[62]), .A (n_181), .B1 (n_179), .B2 (Res_imm[62]));
NAND2_X1 sgo__sro_c62 (.ZN (sgo__sro_n50), .A1 (Res_imm[53]), .A2 (n_60));
NAND2_X1 i_101 (.ZN (n_69), .A1 (n_209), .A2 (n_171));
INV_X1 i_100 (.ZN (n_70), .A (n_69));
AOI21_X1 i_99 (.ZN (n_177), .A (n_46), .B1 (n_70), .B2 (n_202));
NAND4_X1 i_98 (.ZN (n_176), .A1 (n_209), .A2 (n_46), .A3 (n_202), .A4 (n_171));
INV_X1 i_97 (.ZN (n_175), .A (n_176));
NOR2_X1 i_96 (.ZN (p_0[60]), .A1 (n_177), .A2 (n_175));
NAND4_X1 i_95 (.ZN (n_168), .A1 (n_78), .A2 (n_171), .A3 (n_207), .A4 (n_202));
INV_X1 i_94 (.ZN (n_61), .A (n_168));
INV_X1 i_93 (.ZN (n_167), .A (n_205));
INV_X4 i_91 (.ZN (n_68), .A (n_163));
NAND4_X2 i_90 (.ZN (n_162), .A1 (n_68), .A2 (n_160), .A3 (n_204), .A4 (n_167));
AOI21_X1 i_89 (.ZN (p_0[59]), .A (n_61), .B1 (n_162), .B2 (Res_imm[59]));
INV_X1 i_88 (.ZN (n_161), .A (n_162));
NAND4_X1 i_87 (.ZN (n_158), .A1 (n_68), .A2 (n_154), .A3 (n_204), .A4 (n_159));
AOI21_X1 i_86 (.ZN (p_0[58]), .A (n_161), .B1 (n_158), .B2 (Res_imm[58]));
NAND4_X1 i_82 (.ZN (n_157), .A1 (n_209), .A2 (n_160), .A3 (n_204), .A4 (n_165));
INV_X1 i_80 (.ZN (n_156), .A (n_157));
NAND3_X1 i_79 (.ZN (n_155), .A1 (n_68), .A2 (n_204), .A3 (n_159));
AOI22_X1 i_78 (.ZN (p_0[57]), .A1 (n_155), .A2 (opt_ipoPP_6), .B1 (n_156), .B2 (n_149));
NAND3_X1 i_77 (.ZN (n_49), .A1 (n_209), .A2 (n_204), .A3 (n_165));
AOI22_X1 i_73 (.ZN (p_0[56]), .A1 (n_157), .A2 (Res_imm[56]), .B1 (n_65), .B2 (n_159));
NAND3_X1 i_72 (.ZN (n_151), .A1 (n_68), .A2 (n_164), .A3 (n_204));
AOI21_X1 i_71 (.ZN (p_0[55]), .A (n_156), .B1 (n_151), .B2 (Res_imm[55]));
NAND2_X1 i_70 (.ZN (n_150), .A1 (n_65), .A2 (n_144));
AOI22_X1 i_69 (.ZN (p_0[54]), .A1 (n_65), .A2 (n_164), .B1 (Res_imm[54]), .B2 (n_150));
NAND2_X4 i_68 (.ZN (n_82), .A1 (n_87), .A2 (n_142));
INV_X1 i_67 (.ZN (n_27), .A (n_147));
NOR2_X1 i_66 (.ZN (n_25), .A1 (n_147), .A2 (Res_imm[38]));
NAND3_X1 i_64 (.ZN (n_145), .A1 (n_184), .A2 (n_172), .A3 (n_170));
AOI22_X1 i_62 (.ZN (p_0[61]), .A1 (n_61), .A2 (n_200), .B1 (Res_imm[61]), .B2 (n_26));
INV_X2 i_61 (.ZN (n_65), .A (n_49));
INV_X1 i_60 (.ZN (n_62), .A (opt_ipoPP_7));
NAND3_X1 i_59 (.ZN (n_60), .A1 (n_68), .A2 (n_62), .A3 (n_204));
INV_X1 i_144 (.ZN (n_59), .A (Res_imm[50]));
INV_X1 i_143 (.ZN (n_58), .A (Res_imm[49]));
INV_X1 i_142 (.ZN (n_57), .A (Res_imm[48]));
NAND4_X2 i_141 (.ZN (n_56), .A1 (n_68), .A2 (n_59), .A3 (n_58), .A4 (n_57));
AOI21_X1 i_140 (.ZN (p_0[51]), .A (n_65), .B1 (n_56), .B2 (Res_imm[51]));
NAND3_X1 i_139 (.ZN (n_55), .A1 (n_68), .A2 (n_58), .A3 (n_57));
NAND2_X1 i_138 (.ZN (n_54), .A1 (n_55), .A2 (Res_imm[50]));
NAND2_X1 i_137 (.ZN (n_53), .A1 (n_54), .A2 (n_56));
INV_X1 i_136 (.ZN (p_0[50]), .A (n_53));
NAND2_X1 i_135 (.ZN (n_52), .A1 (n_68), .A2 (n_57));
NAND2_X1 i_134 (.ZN (n_51), .A1 (n_52), .A2 (Res_imm[49]));
NAND2_X1 i_133 (.ZN (n_50), .A1 (n_51), .A2 (n_55));
INV_X1 i_132 (.ZN (p_0[49]), .A (n_50));
INV_X1 i_57 (.ZN (n_113), .A (n_116));
NAND2_X1 i_113 (.ZN (n_75), .A1 (n_78), .A2 (n_171));
INV_X1 i_112 (.ZN (n_43), .A (n_52));
INV_X1 i_55 (.ZN (n_45), .A (n_60));
INV_X1 i_54 (.ZN (n_46), .A (Res_imm[60]));
INV_X1 i_53 (.ZN (n_42), .A (Res_imm[30]));
NAND2_X1 i_52 (.ZN (n_88), .A1 (n_13), .A2 (n_194));
INV_X1 i_51 (.ZN (n_89), .A (n_88));
INV_X1 i_50 (.ZN (n_90), .A (n_13));
NAND2_X1 i_49 (.ZN (n_84), .A1 (n_87), .A2 (n_42));
INV_X1 i_48 (.ZN (n_85), .A (n_84));
INV_X1 i_47 (.ZN (n_83), .A (n_82));
INV_X2 i_46 (.ZN (n_78), .A (n_77));
NAND2_X1 i_44 (.ZN (n_26), .A1 (n_61), .A2 (n_46));
INV_X1 i_43 (.ZN (n_98), .A (n_131));
INV_X1 i_65 (.ZN (n_76), .A (n_75));
AOI21_X1 i_41 (.ZN (p_0[52]), .A (n_45), .B1 (opt_ipoPP_7), .B2 (n_49));
AOI21_X1 i_85 (.ZN (p_0[48]), .A (n_43), .B1 (Res_imm[48]), .B2 (n_163));
AOI21_X1 i_84 (.ZN (p_0[47]), .A (n_68), .B1 (Res_imm[47]), .B2 (n_69));
AOI21_X1 i_83 (.ZN (p_0[46]), .A (n_70), .B1 (Res_imm[46]), .B2 (n_71));
AOI21_X1 i_81 (.ZN (p_0[44]), .A (n_74), .B1 (Res_imm[44]), .B2 (n_75));
NOR2_X1 i_39 (.ZN (n_33), .A1 (n_145), .A2 (n_77));
INV_X1 i_75 (.ZN (n_32), .A (n_33));
AOI21_X1 i_74 (.ZN (p_0[43]), .A (n_76), .B1 (Res_imm[43]), .B2 (n_32));
AOI21_X1 i_37 (.ZN (p_0[42]), .A (n_33), .B1 (Res_imm[42]), .B2 (n_47));
AOI21_X1 i_36 (.ZN (p_0[40]), .A (n_37), .B1 (Res_imm[40]), .B2 (n_77));
INV_X1 i_35 (.ZN (n_24), .A (n_25));
AOI21_X1 i_34 (.ZN (p_0[39]), .A (n_78), .B1 (Res_imm[39]), .B2 (n_24));
AOI21_X1 i_33 (.ZN (p_0[37]), .A (n_27), .B1 (Res_imm[37]), .B2 (n_28));
AOI21_X1 i_32 (.ZN (p_0[36]), .A (n_29), .B1 (Res_imm[36]), .B2 (n_30));
NOR2_X2 i_31 (.ZN (n_23), .A1 (Res_imm[32]), .A2 (n_82));
INV_X1 i_30 (.ZN (n_22), .A (n_23));
NOR2_X4 i_29 (.ZN (n_21), .A1 (Res_imm[33]), .A2 (n_22));
INV_X2 i_28 (.ZN (n_20), .A (n_21));
NOR2_X2 i_27 (.ZN (n_19), .A1 (Res_imm[34]), .A2 (n_20));
INV_X1 i_26 (.ZN (n_18), .A (n_19));
AOI21_X1 i_25 (.ZN (p_0[35]), .A (n_31), .B1 (Res_imm[35]), .B2 (n_18));
AOI21_X1 i_22 (.ZN (p_0[34]), .A (n_19), .B1 (Res_imm[34]), .B2 (n_20));
AOI21_X1 i_21 (.ZN (p_0[33]), .A (n_21), .B1 (Res_imm[33]), .B2 (n_22));
AOI21_X1 i_20 (.ZN (p_0[32]), .A (n_23), .B1 (Res_imm[32]), .B2 (n_82));
AOI21_X1 i_19 (.ZN (p_0[31]), .A (n_83), .B1 (Res_imm[31]), .B2 (n_84));
AOI21_X1 i_18 (.ZN (p_0[30]), .A (n_85), .B1 (Res_imm[30]), .B2 (n_7));
AOI21_X1 i_17 (.ZN (p_0[29]), .A (n_87), .B1 (Res_imm[29]), .B2 (n_88));
AOI21_X1 i_16 (.ZN (p_0[28]), .A (n_89), .B1 (Res_imm[28]), .B2 (n_90));
AOI21_X1 i_15 (.ZN (p_0[27]), .A (n_13), .B1 (Res_imm[27]), .B2 (n_137));
AOI21_X1 i_14 (.ZN (p_0[24]), .A (n_135), .B1 (Res_imm[24]), .B2 (n_98));
AOI21_X1 i_38 (.ZN (p_0[21]), .A (n_128), .B1 (Res_imm[21]), .B2 (n_123));
AOI21_X1 i_13 (.ZN (p_0[18]), .A (n_120), .B1 (Res_imm[18]), .B2 (n_114));
AOI21_X1 i_12 (.ZN (p_0[16]), .A (n_113), .B1 (Res_imm[16]), .B2 (n_109));
AOI21_X1 i_24 (.ZN (p_0[13]), .A (n_105), .B1 (Res_imm[13]), .B2 (n_104));
AOI21_X1 i_23 (.ZN (p_0[12]), .A (n_103), .B1 (Res_imm[12]), .B2 (n_101));
AOI21_X1 i_11 (.ZN (p_0[9]), .A (n_95), .B1 (Res_imm[9]), .B2 (n_93));
AOI21_X1 i_10 (.ZN (p_0[8]), .A (n_94), .B1 (Res_imm[8]), .B2 (n_92));
NOR2_X1 i_9 (.ZN (n_5), .A1 (Res_imm[4]), .A2 (n_48));
INV_X1 i_8 (.ZN (n_4), .A (n_5));
NOR2_X1 i_7 (.ZN (n_3), .A1 (Res_imm[5]), .A2 (n_4));
INV_X1 i_6 (.ZN (n_2), .A (n_3));
AOI21_X1 i_5 (.ZN (p_0[6]), .A (n_41), .B1 (Res_imm[6]), .B2 (n_2));
AOI21_X1 i_4 (.ZN (p_0[5]), .A (n_3), .B1 (Res_imm[5]), .B2 (n_4));
AOI21_X1 i_3 (.ZN (p_0[4]), .A (n_5), .B1 (Res_imm[4]), .B2 (n_48));
AOI21_X1 i_2 (.ZN (p_0[3]), .A (n_63), .B1 (Res_imm[3]), .B2 (n_64));
AOI21_X1 i_1 (.ZN (p_0[2]), .A (n_66), .B1 (Res_imm[2]), .B2 (n_79));
AOI21_X1 i_0 (.ZN (p_0[1]), .A (n_80), .B1 (Res_imm[1]), .B2 (Res_imm[0]));

endmodule //datapath__0_3

module datapath__0_2 (opt_ipoPP_0, B_imm, A_imm, Res_imm);

output [63:0] Res_imm;
input [31:0] A_imm;
input [31:0] B_imm;
input opt_ipoPP_0;
wire n_0;
wire n_1;
wire n_2;
wire n_1271;
wire n_6740;
wire n_6836;
wire n_4366;
wire n_3554;
wire n_3;
wire n_1265;
wire n_1270;
wire n_1268;
wire n_1264;
wire n_4;
wire n_1273;
wire n_1272;
wire n_1262;
wire n_5;
wire n_1281;
wire n_1280;
wire n_1260;
wire n_6;
wire n_1288;
wire n_1287;
wire n_1258;
wire n_7;
wire n_1297;
wire n_1296;
wire n_8;
wire n_1256;
wire n_1306;
wire n_1253;
wire n_9;
wire n_1251;
wire n_1315;
wire n_1314;
wire n_1250;
wire n_10;
wire n_1324;
wire n_1328;
wire n_11;
wire n_1249;
wire n_1339;
wire n_1334;
wire n_1248;
wire n_12;
wire n_13;
wire n_1449;
wire n_1246;
wire n_14;
wire n_16;
wire n_15;
wire n_1491;
wire n_17;
wire n_1530;
wire n_1488;
wire n_18;
wire n_1244;
wire n_19;
wire n_1537;
wire n_1535;
wire n_20;
wire n_21;
wire n_22;
wire n_1238;
wire n_1594;
wire n_1534;
wire n_24;
wire n_23;
wire n_1243;
wire n_1233;
wire n_1240;
wire n_26;
wire n_25;
wire n_1235;
wire n_1718;
wire n_1229;
wire n_1226;
wire n_27;
wire n_39;
wire n_36;
wire n_28;
wire n_34;
wire n_29;
wire n_30;
wire n_40;
wire n_1144;
wire n_33;
wire n_31;
wire n_42;
wire n_1128;
wire n_44;
wire n_32;
wire n_41;
wire n_35;
wire n_37;
wire n_1795;
wire n_38;
wire n_1141;
wire n_1146;
wire n_1140;
wire n_1153;
wire n_1162;
wire n_1145;
wire n_43;
wire n_1161;
wire n_1185;
wire n_1133;
wire n_1129;
wire n_45;
wire n_1223;
wire n_1222;
wire n_92;
wire n_46;
wire n_47;
wire n_1116;
wire n_2105;
wire n_48;
wire n_56;
wire n_49;
wire n_50;
wire n_59;
wire n_2215;
wire n_51;
wire n_52;
wire n_55;
wire n_61;
wire n_2328;
wire n_53;
wire n_54;
wire n_64;
wire n_60;
wire n_57;
wire n_58;
wire n_1117;
wire n_2217;
wire n_62;
wire n_63;
wire n_2329;
wire n_2339;
wire n_2333;
wire n_1121;
wire n_90;
wire n_65;
wire n_2631;
wire n_74;
wire n_66;
wire n_72;
wire n_67;
wire n_75;
wire n_2769;
wire n_71;
wire n_68;
wire n_2928;
wire n_1104;
wire n_69;
wire n_70;
wire n_78;
wire n_77;
wire n_76;
wire n_73;
wire n_2774;
wire n_2636;
wire n_2633;
wire n_2931;
wire n_2923;
wire n_2775;
wire n_2771;
wire n_3077;
wire n_1105;
wire n_88;
wire n_79;
wire n_1013;
wire n_1060;
wire n_80;
wire n_82;
wire n_81;
wire n_93;
wire n_1009;
wire n_87;
wire n_1012;
wire n_85;
wire n_83;
wire n_96;
wire n_95;
wire n_97;
wire n_84;
wire n_94;
wire n_86;
wire n_89;
wire n_1102;
wire n_91;
wire n_1119;
wire n_1114;
wire n_2323;
wire n_2104;
wire n_1138;
wire n_1131;
wire n_1124;
wire n_1024;
wire n_1020;
wire n_1038;
wire n_1023;
wire n_1019;
wire n_1005;
wire n_1037;
wire n_1002;
wire n_98;
wire n_1000;
wire n_3992;
wire n_99;
wire n_104;
wire n_100;
wire n_4252;
wire n_4217;
wire n_103;
wire n_101;
wire n_3986;
wire n_4229;
wire n_108;
wire n_102;
wire n_107;
wire n_106;
wire n_105;
wire n_3984;
wire n_4222;
wire n_109;
wire n_163;
wire n_5724;
wire n_993;
wire n_110;
wire n_111;
wire n_119;
wire n_990;
wire n_5689;
wire n_112;
wire n_118;
wire n_985;
wire n_5658;
wire n_115;
wire n_113;
wire n_117;
wire n_988;
wire n_114;
wire n_982;
wire n_116;
wire n_5666;
wire n_122;
wire n_121;
wire n_120;
wire CLOCK_opt_ipo_n363;
wire n_124;
wire n_139;
wire n_7465;
wire n_976;
wire n_133;
wire n_141;
wire n_127;
wire n_125;
wire n_129;
wire n_126;
wire n_972;
wire n_6943;
wire n_128;
wire n_145;
wire n_977;
wire n_130;
wire n_6936;
wire n_131;
wire n_135;
wire n_132;
wire n_144;
wire n_971;
wire n_146;
wire n_134;
wire n_143;
wire n_136;
wire n_137;
wire n_138;
wire n_980;
wire n_140;
wire n_142;
wire n_6964;
wire n_147;
wire n_148;
wire n_162;
wire n_961;
wire n_5505;
wire n_154;
wire n_166;
wire n_151;
wire n_149;
wire n_153;
wire n_5112;
wire n_150;
wire n_170;
wire n_5121;
wire n_152;
wire n_964;
wire n_155;
wire n_156;
wire n_158;
wire n_157;
wire n_169;
wire n_159;
wire n_171;
wire n_168;
wire n_160;
wire n_161;
wire n_164;
wire n_165;
wire n_3981;
wire n_967;
wire n_6934;
wire n_167;
wire n_954;
wire n_5139;
wire n_959;
wire n_958;
wire n_172;
wire n_173;
wire n_951;
wire n_855;
wire n_589;
wire n_174;
wire n_184;
wire n_761;
wire n_594;
wire n_183;
wire n_176;
wire n_177;
wire n_593;
wire n_678;
wire n_178;
wire n_181;
wire n_179;
wire n_180;
wire n_182;
wire n_600;
wire n_588;
wire n_186;
wire n_185;
wire n_187;
wire n_586;
wire n_521;
wire n_203;
wire n_188;
wire n_202;
wire n_200;
wire n_189;
wire n_192;
wire n_190;
wire n_191;
wire n_193;
wire n_261;
wire n_355;
wire n_263;
wire n_363;
wire n_195;
wire n_194;
wire n_206;
wire n_197;
wire n_199;
wire n_196;
wire n_205;
wire n_198;
wire n_264;
wire n_201;
wire n_204;
wire n_526;
wire n_523;
wire n_258;
wire n_379;
wire CLOCK_opt_ipo_n452;
wire n_229;
wire n_227;
wire n_208;
wire n_211;
wire n_209;
wire n_210;
wire n_212;
wire n_256;
wire n_251;
wire n_273;
wire n_269;
wire n_214;
wire n_213;
wire n_224;
wire n_216;
wire n_218;
wire n_217;
wire n_215;
wire n_291;
wire n_249;
wire n_220;
wire n_219;
wire n_233;
wire n_222;
wire n_226;
wire n_221;
wire n_232;
wire n_223;
wire n_254;
wire n_225;
wire n_228;
wire n_230;
wire n_231;
wire n_257;
wire n_353;
wire n_250;
wire n_319;
wire n_234;
wire n_244;
wire n_235;
wire n_236;
wire n_242;
wire n_8975;
wire n_239;
wire n_238;
wire n_241;
wire n_240;
wire n_9027;
wire n_9026;
wire n_8976;
wire n_243;
wire n_9025;
wire n_245;
wire n_266;
wire n_246;
wire n_267;
wire n_247;
wire n_255;
wire n_248;
wire n_316;
wire n_293;
wire n_322;
wire n_320;
wire n_253;
wire n_280;
wire n_252;
wire n_274;
wire n_286;
wire n_289;
wire n_271;
wire n_270;
wire n_265;
wire n_259;
wire n_407;
wire n_380;
wire n_260;
wire n_262;
wire n_365;
wire n_378;
wire n_558;
wire n_360;
wire n_357;
wire n_268;
wire n_430;
wire n_431;
wire n_408;
wire n_272;
wire n_275;
wire n_279;
wire n_278;
wire n_276;
wire n_277;
wire n_301;
wire n_306;
wire n_305;
wire n_281;
wire n_284;
wire n_282;
wire n_283;
wire n_486;
wire n_454;
wire n_487;
wire n_285;
wire n_326;
wire n_329;
wire n_330;
wire n_287;
wire n_288;
wire n_298;
wire n_299;
wire n_295;
wire n_290;
wire n_315;
wire n_292;
wire n_294;
wire n_297;
wire n_296;
wire n_335;
wire n_333;
wire n_324;
wire n_300;
wire n_313;
wire n_304;
wire n_302;
wire n_441;
wire n_303;
wire n_442;
wire n_433;
wire n_309;
wire n_307;
wire n_507;
wire n_308;
wire n_519;
wire n_504;
wire n_310;
wire n_342;
wire n_311;
wire n_312;
wire n_341;
wire n_344;
wire n_314;
wire n_8984;
wire n_8983;
wire n_8986;
wire n_323;
wire n_317;
wire n_318;
wire n_345;
wire n_346;
wire n_321;
wire n_8979;
wire n_9009;
wire n_9008;
wire n_334;
wire n_325;
wire n_327;
wire n_328;
wire n_8990;
wire n_8992;
wire n_8989;
wire n_331;
wire n_9003;
wire n_9005;
wire n_436;
wire n_437;
wire n_332;
wire n_435;
wire n_337;
wire n_340;
wire n_336;
wire n_339;
wire n_338;
wire n_9000;
wire n_9002;
wire n_8999;
wire n_446;
wire n_447;
wire n_343;
wire n_445;
wire n_350;
wire n_347;
wire n_348;
wire n_349;
wire n_9017;
wire n_9019;
wire n_9016;
wire n_351;
wire n_8981;
wire n_352;
wire n_8995;
wire n_8996;
wire n_354;
wire n_359;
wire n_356;
wire n_358;
wire n_371;
wire n_366;
wire n_370;
wire n_381;
wire n_361;
wire n_362;
wire n_385;
wire n_384;
wire n_364;
wire n_369;
wire n_367;
wire n_389;
wire n_368;
wire n_391;
wire n_392;
wire n_373;
wire n_376;
wire n_372;
wire n_374;
wire n_375;
wire n_533;
wire n_532;
wire n_529;
wire n_399;
wire n_377;
wire n_401;
wire n_402;
wire n_527;
wire n_559;
wire n_382;
wire n_383;
wire n_410;
wire n_412;
wire n_413;
wire n_386;
wire n_397;
wire n_387;
wire n_388;
wire n_390;
wire n_571;
wire n_570;
wire n_563;
wire n_395;
wire n_393;
wire n_541;
wire n_394;
wire n_540;
wire n_537;
wire n_396;
wire n_416;
wire n_419;
wire n_418;
wire n_398;
wire n_400;
wire n_474;
wire n_475;
wire n_473;
wire n_405;
wire n_403;
wire n_581;
wire n_575;
wire n_404;
wire n_582;
wire n_566;
wire n_564;
wire n_406;
wire n_568;
wire n_428;
wire n_409;
wire n_411;
wire n_456;
wire n_469;
wire n_468;
wire n_425;
wire n_414;
wire n_415;
wire n_498;
wire n_417;
wire n_499;
wire n_497;
wire n_420;
wire n_423;
wire n_421;
wire n_422;
wire n_465;
wire n_467;
wire n_464;
wire n_547;
wire n_424;
wire n_550;
wire n_545;
wire n_426;
wire n_489;
wire n_492;
wire n_427;
wire n_493;
wire n_429;
wire n_452;
wire n_432;
wire n_439;
wire n_434;
wire n_9038;
wire n_8794;
wire n_9004;
wire n_8972;
wire n_438;
wire n_440;
wire n_449;
wire n_443;
wire n_444;
wire n_9020;
wire n_9021;
wire n_8974;
wire n_9037;
wire n_448;
wire n_450;
wire n_451;
wire n_459;
wire n_462;
wire n_458;
wire n_453;
wire n_485;
wire n_455;
wire n_457;
wire n_461;
wire n_479;
wire n_460;
wire n_8994;
wire n_8993;
wire n_478;
wire n_480;
wire n_463;
wire n_466;
wire n_7912;
wire n_470;
wire n_483;
wire n_471;
wire n_472;
wire n_476;
wire n_481;
wire n_477;
wire n_8821;
wire n_482;
wire n_555;
wire n_554;
wire n_556;
wire n_484;
wire n_517;
wire n_518;
wire n_515;
wire n_502;
wire n_488;
wire n_490;
wire n_511;
wire n_491;
wire n_512;
wire n_510;
wire n_494;
wire n_495;
wire n_496;
wire n_501;
wire n_578;
wire n_500;
wire n_8907;
wire n_577;
wire n_579;
wire n_503;
wire n_506;
wire n_505;
wire n_508;
wire n_513;
wire n_509;
wire n_9006;
wire n_8948;
wire n_516;
wire n_514;
wire n_520;
wire n_525;
wire n_522;
wire n_636;
wire n_524;
wire n_606;
wire n_635;
wire n_557;
wire n_528;
wire n_531;
wire n_530;
wire n_663;
wire n_662;
wire n_641;
wire n_536;
wire n_534;
wire n_535;
wire n_631;
wire n_618;
wire n_628;
wire n_539;
wire n_669;
wire n_677;
wire n_538;
wire n_668;
wire n_542;
wire n_552;
wire n_543;
wire n_544;
wire n_546;
wire n_548;
wire n_549;
wire n_673;
wire n_672;
wire n_674;
wire n_551;
wire n_553;
wire n_8767;
wire n_560;
wire n_562;
wire n_613;
wire n_561;
wire n_608;
wire n_612;
wire n_569;
wire n_565;
wire n_621;
wire n_626;
wire n_622;
wire n_567;
wire n_643;
wire n_650;
wire n_574;
wire n_572;
wire n_653;
wire n_573;
wire n_652;
wire n_642;
wire n_580;
wire n_576;
wire n_8958;
wire n_584;
wire n_583;
wire n_585;
wire n_657;
wire n_656;
wire n_658;
wire n_587;
wire n_598;
wire n_591;
wire n_597;
wire n_603;
wire n_601;
wire n_858;
wire n_860;
wire n_590;
wire n_856;
wire n_5175;
wire n_592;
wire n_596;
wire n_680;
wire n_685;
wire n_682;
wire n_595;
wire n_763;
wire n_765;
wire n_768;
wire n_599;
wire n_602;
wire n_717;
wire n_686;
wire n_720;
wire n_605;
wire n_604;
wire n_607;
wire n_634;
wire n_611;
wire n_609;
wire n_743;
wire n_723;
wire n_610;
wire n_744;
wire n_617;
wire n_614;
wire n_615;
wire n_713;
wire n_696;
wire n_616;
wire n_712;
wire n_627;
wire n_619;
wire n_620;
wire n_623;
wire n_624;
wire n_625;
wire n_701;
wire n_700;
wire n_702;
wire n_629;
wire n_630;
wire n_632;
wire n_750;
wire n_633;
wire n_751;
wire n_758;
wire n_707;
wire n_705;
wire n_698;
wire n_640;
wire n_637;
wire n_638;
wire n_691;
wire n_687;
wire n_639;
wire n_692;
wire n_661;
wire n_651;
wire n_646;
wire n_644;
wire n_649;
wire n_648;
wire n_645;
wire n_756;
wire n_755;
wire n_757;
wire n_647;
wire n_8906;
wire n_654;
wire n_659;
wire n_655;
wire n_730;
wire n_725;
wire n_660;
wire n_729;
wire n_666;
wire n_664;
wire n_665;
wire n_732;
wire n_733;
wire n_724;
wire n_667;
wire n_670;
wire n_675;
wire n_671;
wire n_8957;
wire n_676;
wire n_738;
wire n_739;
wire n_736;
wire n_679;
wire n_681;
wire n_771;
wire n_817;
wire n_770;
wire n_684;
wire n_683;
wire n_689;
wire n_688;
wire n_792;
wire n_774;
wire n_775;
wire n_690;
wire n_695;
wire n_693;
wire n_694;
wire n_846;
wire n_826;
wire n_847;
wire n_711;
wire n_697;
wire n_703;
wire n_699;
wire n_704;
wire n_706;
wire n_708;
wire n_709;
wire n_788;
wire n_789;
wire n_710;
wire n_787;
wire n_714;
wire n_715;
wire n_835;
wire n_833;
wire n_827;
wire n_782;
wire n_716;
wire n_781;
wire n_785;
wire n_718;
wire n_719;
wire n_721;
wire n_821;
wire n_722;
wire n_819;
wire n_853;
wire n_742;
wire n_731;
wire n_728;
wire n_726;
wire n_727;
wire n_830;
wire n_829;
wire n_831;
wire n_8893;
wire n_8859;
wire n_734;
wire n_741;
wire n_735;
wire n_737;
wire n_839;
wire n_740;
wire n_840;
wire n_838;
wire n_810;
wire n_811;
wire n_808;
wire n_745;
wire n_748;
wire n_746;
wire n_795;
wire n_747;
wire n_794;
wire n_806;
wire n_749;
wire n_753;
wire n_752;
wire n_754;
wire n_8860;
wire n_799;
wire n_760;
wire n_759;
wire n_798;
wire n_800;
wire n_762;
wire n_764;
wire n_903;
wire n_861;
wire n_904;
wire n_767;
wire n_766;
wire n_769;
wire n_814;
wire n_772;
wire n_773;
wire n_779;
wire n_776;
wire n_777;
wire n_944;
wire n_778;
wire n_940;
wire n_946;
wire n_780;
wire n_783;
wire n_912;
wire n_913;
wire n_784;
wire n_911;
wire n_786;
wire n_790;
wire n_893;
wire n_791;
wire n_892;
wire n_894;
wire n_793;
wire n_803;
wire n_796;
wire n_797;
wire n_880;
wire n_802;
wire n_801;
wire n_879;
wire n_881;
wire n_804;
wire n_896;
wire n_805;
wire n_890;
wire n_897;
wire n_807;
wire n_809;
wire n_922;
wire n_813;
wire n_812;
wire n_921;
wire n_923;
wire n_815;
wire n_816;
wire n_868;
wire n_866;
wire n_863;
wire n_818;
wire n_852;
wire n_820;
wire n_887;
wire n_823;
wire n_825;
wire n_822;
wire n_886;
wire n_824;
wire n_873;
wire n_845;
wire n_832;
wire n_828;
wire n_8525;
wire n_834;
wire n_842;
wire n_836;
wire n_837;
wire n_841;
wire n_843;
wire n_844;
wire n_928;
wire n_926;
wire n_931;
wire n_850;
wire n_848;
wire n_876;
wire n_884;
wire n_849;
wire n_875;
wire n_917;
wire n_851;
wire n_918;
wire n_909;
wire n_854;
wire n_935;
wire n_936;
wire n_908;
wire n_857;
wire n_5171;
wire n_5173;
wire n_859;
wire n_862;
wire n_865;
wire n_864;
wire n_5217;
wire n_5246;
wire n_5216;
wire n_867;
wire n_870;
wire n_872;
wire n_869;
wire n_5338;
wire n_871;
wire n_5321;
wire n_5335;
wire n_885;
wire n_874;
wire n_882;
wire n_877;
wire n_878;
wire n_5231;
wire n_883;
wire n_5235;
wire n_5229;
wire n_889;
wire n_902;
wire n_5226;
wire n_888;
wire n_901;
wire n_895;
wire n_891;
wire n_8423;
wire n_898;
wire n_5242;
wire n_900;
wire n_899;
wire n_5241;
wire n_5243;
wire n_5225;
wire n_5223;
wire n_907;
wire n_905;
wire n_906;
wire n_5273;
wire n_5368;
wire n_5271;
wire n_934;
wire n_916;
wire n_910;
wire n_8956;
wire n_8892;
wire n_914;
wire n_5328;
wire n_5329;
wire n_915;
wire n_5327;
wire n_924;
wire n_919;
wire n_920;
wire n_925;
wire n_927;
wire n_929;
wire n_5262;
wire n_5263;
wire n_930;
wire n_5261;
wire n_5349;
wire n_933;
wire n_932;
wire n_5348;
wire n_5350;
wire n_939;
wire n_937;
wire n_938;
wire n_5249;
wire n_5248;
wire n_5265;
wire n_943;
wire n_941;
wire n_5324;
wire n_942;
wire n_5323;
wire n_5333;
wire n_945;
wire n_948;
wire n_950;
wire n_5345;
wire n_947;
wire n_5255;
wire n_5259;
wire n_949;
wire n_5253;
wire n_5344;
wire n_5358;
wire n_952;
wire n_995;
wire n_3980;
wire n_953;
wire n_957;
wire n_960;
wire n_966;
wire n_956;
wire n_5137;
wire n_955;
wire n_5140;
wire n_5168;
wire n_5172;
wire n_5122;
wire n_5130;
wire n_5135;
wire n_5138;
wire n_962;
wire n_963;
wire n_5506;
wire n_5509;
wire n_5655;
wire n_7200;
wire n_965;
wire n_5114;
wire n_5116;
wire n_968;
wire n_6935;
wire n_969;
wire n_970;
wire n_974;
wire n_979;
wire n_7000;
wire n_6997;
wire n_6965;
wire n_6975;
wire n_6963;
wire n_6961;
wire n_973;
wire n_6954;
wire n_6941;
wire n_6952;
wire n_975;
wire n_7733;
wire n_7467;
wire n_7737;
wire n_978;
wire n_6938;
wire n_6939;
wire n_6942;
wire n_981;
wire n_989;
wire n_5668;
wire n_983;
wire n_5688;
wire n_984;
wire n_7470;
wire n_7476;
wire n_7475;
wire n_5660;
wire n_987;
wire n_986;
wire n_5669;
wire n_5678;
wire n_5675;
wire n_5665;
wire n_992;
wire n_991;
wire n_5690;
wire n_6089;
wire n_5692;
wire n_5695;
wire n_5726;
wire n_994;
wire n_6009;
wire n_6010;
wire n_997;
wire n_999;
wire n_1001;
wire n_3998;
wire n_3993;
wire n_3996;
wire n_1003;
wire n_1015;
wire n_1004;
wire n_1011;
wire n_1007;
wire n_1010;
wire n_1006;
wire n_1008;
wire n_1028;
wire n_1025;
wire n_1062;
wire n_1058;
wire n_1018;
wire n_1014;
wire n_3081;
wire n_1063;
wire n_1061;
wire n_1101;
wire n_1016;
wire n_1017;
wire n_1022;
wire n_1021;
wire n_1039;
wire n_1054;
wire n_1057;
wire n_1027;
wire n_1026;
wire n_1029;
wire n_1031;
wire n_1036;
wire n_1030;
wire n_1092;
wire n_1070;
wire n_1094;
wire n_1032;
wire n_1043;
wire n_1033;
wire n_1045;
wire n_1044;
wire n_4015;
wire n_1035;
wire n_1034;
wire n_4021;
wire n_4209;
wire n_4097;
wire n_4024;
wire n_1042;
wire n_1041;
wire n_1040;
wire n_4016;
wire n_4022;
wire n_1049;
wire n_1047;
wire n_1083;
wire n_1046;
wire n_1048;
wire n_1086;
wire n_1076;
wire n_1050;
wire n_1053;
wire n_1051;
wire n_1052;
wire n_4394;
wire n_4392;
wire n_4313;
wire n_1055;
wire n_1056;
wire n_4006;
wire n_4007;
wire n_4001;
wire n_1059;
wire n_4214;
wire n_4216;
wire n_4000;
wire n_3082;
wire n_1064;
wire n_1066;
wire n_1069;
wire n_3112;
wire n_3088;
wire n_1065;
wire n_3115;
wire n_1068;
wire n_1067;
wire n_1071;
wire n_1074;
wire n_1073;
wire n_1072;
wire n_1088;
wire n_1087;
wire n_3124;
wire n_1075;
wire n_1078;
wire n_1077;
wire n_4320;
wire n_4319;
wire n_4316;
wire n_4315;
wire n_1079;
wire n_1080;
wire n_1081;
wire n_1082;
wire n_4432;
wire n_4474;
wire n_4473;
wire n_1084;
wire n_1085;
wire n_3128;
wire n_3122;
wire n_1089;
wire n_1091;
wire n_1090;
wire n_4670;
wire n_4730;
wire n_4728;
wire n_4669;
wire n_1093;
wire n_1100;
wire n_1097;
wire n_1095;
wire n_3103;
wire n_1096;
wire n_3106;
wire n_3098;
wire n_1098;
wire n_1099;
wire n_4025;
wire n_4026;
wire n_4034;
wire n_1112;
wire n_1134;
wire n_1107;
wire n_1103;
wire n_2932;
wire n_3135;
wire n_2930;
wire n_1106;
wire n_3079;
wire n_1108;
wire n_1111;
wire n_1109;
wire n_2635;
wire n_1110;
wire n_2929;
wire n_1113;
wire n_1122;
wire n_2325;
wire n_1115;
wire n_2218;
wire n_2212;
wire n_2106;
wire n_1118;
wire n_2216;
wire n_1120;
wire n_1123;
wire n_1125;
wire n_1127;
wire n_1126;
wire n_1186;
wire n_1130;
wire n_1132;
wire n_1187;
wire n_1221;
wire n_1219;
wire n_1136;
wire n_1137;
wire n_1156;
wire n_1139;
wire n_1143;
wire n_1142;
wire n_1147;
wire n_1149;
wire n_1152;
wire n_1900;
wire n_1894;
wire n_1148;
wire n_1898;
wire n_1150;
wire n_1151;
wire n_1173;
wire n_1172;
wire n_1165;
wire n_1155;
wire n_1154;
wire n_1163;
wire n_1182;
wire n_1181;
wire n_1184;
wire n_1157;
wire n_1158;
wire n_1160;
wire n_1159;
wire n_1164;
wire n_1166;
wire n_1169;
wire n_1167;
wire n_1168;
wire n_1205;
wire n_1200;
wire n_1207;
wire n_1170;
wire n_1171;
wire n_1210;
wire n_1209;
wire n_1212;
wire n_1958;
wire n_1175;
wire n_1177;
wire n_2022;
wire n_1180;
wire n_1174;
wire n_1176;
wire n_2021;
wire n_2019;
wire n_2133;
wire n_1179;
wire n_1178;
wire n_2139;
wire n_2140;
wire n_2143;
wire n_2176;
wire n_2141;
wire n_2134;
wire n_1189;
wire n_1196;
wire n_1198;
wire n_1183;
wire n_1188;
wire n_1195;
wire n_1193;
wire n_1190;
wire n_2121;
wire n_1192;
wire n_1191;
wire n_2125;
wire n_2126;
wire n_2132;
wire n_2127;
wire n_1194;
wire n_1214;
wire n_1197;
wire n_1199;
wire n_1213;
wire n_1201;
wire n_1204;
wire n_1202;
wire n_1203;
wire n_2290;
wire n_2289;
wire n_2255;
wire n_1211;
wire n_1206;
wire n_1208;
wire n_2377;
wire n_2410;
wire n_2409;
wire n_1956;
wire n_1954;
wire n_1215;
wire n_1218;
wire n_1216;
wire n_2253;
wire n_1217;
wire n_2249;
wire n_2251;
wire n_2252;
wire n_1220;
wire n_2111;
wire n_2109;
wire n_2112;
wire n_2114;
wire n_2108;
wire n_2107;
wire n_2210;
wire n_2207;
wire n_1225;
wire n_1224;
wire n_1717;
wire n_1227;
wire n_1228;
wire n_1230;
wire n_1796;
wire n_1720;
wire n_1232;
wire n_1231;
wire n_1797;
wire n_1897;
wire n_1892;
wire n_1719;
wire n_1234;
wire n_1242;
wire n_1598;
wire n_1236;
wire n_1237;
wire n_1239;
wire n_1593;
wire n_1595;
wire n_1241;
wire n_1788;
wire n_1793;
wire n_1721;
wire n_1490;
wire n_1245;
wire n_1247;
wire n_1450;
wire n_1487;
wire n_1333;
wire n_1327;
wire n_1313;
wire n_1252;
wire n_1254;
wire n_1255;
wire n_1309;
wire n_1307;
wire n_1310;
wire n_1394;
wire n_1257;
wire n_1259;
wire n_1261;
wire n_1263;
wire n_1267;
wire n_1445;
wire n_1266;
wire n_1269;
wire n_6584;
wire n_1274;
wire n_1277;
wire n_1275;
wire n_1276;
wire n_1360;
wire n_1358;
wire n_1359;
wire n_1278;
wire n_1279;
wire n_1444;
wire n_1446;
wire n_1282;
wire n_1285;
wire n_1283;
wire n_1284;
wire n_1355;
wire n_1353;
wire n_1354;
wire n_1286;
wire n_1434;
wire n_1443;
wire n_1291;
wire n_1305;
wire n_1295;
wire n_1290;
wire n_1289;
wire n_1423;
wire n_1294;
wire n_1349;
wire n_1347;
wire n_1351;
wire n_1292;
wire n_1293;
wire n_1425;
wire n_1433;
wire n_1424;
wire n_1312;
wire n_1301;
wire n_1299;
wire n_1304;
wire n_1303;
wire n_1298;
wire n_1346;
wire n_1362;
wire n_1300;
wire n_1361;
wire n_1302;
wire n_1345;
wire n_1415;
wire n_1414;
wire n_1308;
wire n_1344;
wire n_1371;
wire n_1370;
wire n_1343;
wire n_1311;
wire n_1395;
wire n_1396;
wire n_1413;
wire n_1317;
wire n_1319;
wire n_1323;
wire n_1322;
wire n_1321;
wire n_1316;
wire n_1318;
wire n_1342;
wire n_1380;
wire n_1382;
wire n_1320;
wire n_1390;
wire n_1392;
wire n_1389;
wire n_1393;
wire n_1325;
wire n_1340;
wire n_1326;
wire n_1330;
wire n_1329;
wire n_1332;
wire n_1335;
wire n_1457;
wire n_1462;
wire n_1461;
wire n_1331;
wire n_1459;
wire n_1458;
wire n_1341;
wire n_1336;
wire n_1448;
wire n_1337;
wire n_1338;
wire n_1453;
wire n_1451;
wire n_1455;
wire n_1447;
wire n_1348;
wire n_1409;
wire n_1411;
wire n_1408;
wire n_1350;
wire n_8429;
wire n_1352;
wire n_1357;
wire n_1356;
wire n_6678;
wire n_6677;
wire n_3718;
wire n_1363;
wire n_1365;
wire n_1367;
wire n_1429;
wire n_1364;
wire n_1426;
wire n_1431;
wire n_1366;
wire n_1406;
wire n_1405;
wire n_1412;
wire n_1369;
wire n_1368;
wire n_1375;
wire n_1373;
wire n_1377;
wire n_1418;
wire n_1374;
wire n_1372;
wire n_1417;
wire n_1376;
wire n_1379;
wire n_1478;
wire n_1378;
wire n_1481;
wire n_1482;
wire n_1381;
wire n_1388;
wire n_1386;
wire n_1383;
wire n_1385;
wire n_1401;
wire n_1398;
wire n_1384;
wire n_1403;
wire n_1387;
wire n_1574;
wire n_1563;
wire n_1562;
wire n_1391;
wire n_1466;
wire n_1472;
wire n_1470;
wire n_1465;
wire n_1397;
wire n_1400;
wire n_1399;
wire n_1566;
wire n_1573;
wire n_1565;
wire n_1402;
wire n_8232;
wire n_1404;
wire n_1407;
wire n_1410;
wire n_6817;
wire n_1416;
wire n_1421;
wire n_1420;
wire n_1419;
wire n_1572;
wire n_1571;
wire n_1569;
wire n_1422;
wire n_1570;
wire n_1427;
wire n_1428;
wire n_1430;
wire n_8293;
wire n_1432;
wire n_1440;
wire n_1442;
wire n_1439;
wire n_1437;
wire n_1435;
wire n_1436;
wire n_1441;
wire n_1438;
wire n_1452;
wire n_1498;
wire n_1496;
wire n_1499;
wire n_1501;
wire n_1454;
wire n_1456;
wire n_1504;
wire n_1510;
wire n_1509;
wire n_1460;
wire n_1506;
wire n_1505;
wire n_1485;
wire n_1464;
wire n_1484;
wire n_1483;
wire n_1463;
wire n_1467;
wire n_1469;
wire n_1517;
wire n_1521;
wire n_1468;
wire n_1520;
wire n_1518;
wire n_1522;
wire n_1471;
wire n_1474;
wire n_1480;
wire n_1473;
wire n_1476;
wire n_1475;
wire n_1650;
wire n_1649;
wire n_1647;
wire n_1477;
wire n_1646;
wire n_1479;
wire n_1654;
wire n_1655;
wire n_1653;
wire n_8573;
wire n_1559;
wire n_1576;
wire n_1575;
wire n_1486;
wire n_1560;
wire n_1526;
wire n_1528;
wire n_1493;
wire n_1489;
wire n_1494;
wire n_1529;
wire n_1492;
wire n_1495;
wire n_1497;
wire n_1554;
wire n_1552;
wire n_1556;
wire n_1555;
wire n_1551;
wire n_1503;
wire n_1500;
wire n_1525;
wire n_1523;
wire n_1502;
wire n_1524;
wire n_1656;
wire n_1645;
wire n_1644;
wire n_1507;
wire n_1508;
wire n_1516;
wire n_1514;
wire n_1512;
wire n_1515;
wire n_1511;
wire n_1513;
wire n_1637;
wire n_1641;
wire n_1642;
wire n_1639;
wire n_1638;
wire n_1519;
wire n_1760;
wire n_1761;
wire n_1759;
wire n_1632;
wire n_1634;
wire n_1628;
wire n_1527;
wire n_1542;
wire n_1548;
wire n_1546;
wire n_1544;
wire n_1543;
wire n_1531;
wire n_1539;
wire n_1533;
wire n_1532;
wire n_1540;
wire n_1590;
wire n_1588;
wire n_1604;
wire n_1536;
wire n_1592;
wire n_1538;
wire n_1541;
wire n_1616;
wire n_1621;
wire n_1620;
wire n_1545;
wire n_1547;
wire n_1550;
wire n_1587;
wire n_1585;
wire n_1549;
wire n_1586;
wire n_1553;
wire n_1696;
wire n_1701;
wire n_1702;
wire n_1698;
wire n_1697;
wire n_1558;
wire n_1582;
wire n_1581;
wire n_1557;
wire n_1580;
wire n_1561;
wire n_1564;
wire n_1567;
wire n_1568;
wire n_7691;
wire n_6577;
wire n_8947;
wire n_1578;
wire n_1579;
wire n_8347;
wire n_1577;
wire n_1756;
wire n_1755;
wire n_1753;
wire n_1752;
wire n_1754;
wire n_1757;
wire n_1762;
wire n_1751;
wire n_1750;
wire n_1583;
wire n_1584;
wire n_1695;
wire n_1685;
wire n_1708;
wire n_1589;
wire n_1607;
wire n_1591;
wire n_1609;
wire n_1608;
wire n_1613;
wire n_1612;
wire n_1605;
wire n_1662;
wire n_1665;
wire n_1597;
wire n_1596;
wire n_1599;
wire n_1601;
wire n_1603;
wire n_1600;
wire n_1670;
wire n_1663;
wire n_1671;
wire n_1602;
wire n_1725;
wire n_1723;
wire n_1726;
wire n_1729;
wire n_1722;
wire n_1606;
wire n_1679;
wire n_1683;
wire n_1688;
wire n_1610;
wire n_1611;
wire n_1658;
wire n_1615;
wire n_1660;
wire n_1657;
wire n_1614;
wire n_1617;
wire n_1619;
wire n_1618;
wire n_1747;
wire n_1763;
wire n_1766;
wire n_1748;
wire n_1627;
wire n_1624;
wire n_1623;
wire n_1626;
wire n_1622;
wire n_1846;
wire n_1844;
wire n_1845;
wire n_1625;
wire n_1630;
wire n_1629;
wire n_1851;
wire n_1850;
wire n_1849;
wire n_1631;
wire n_1633;
wire n_1636;
wire n_1643;
wire n_1635;
wire n_1856;
wire n_1855;
wire n_1854;
wire n_1640;
wire n_8645;
wire n_1648;
wire n_1652;
wire n_1651;
wire n_8511;
wire n_8644;
wire n_1659;
wire n_1745;
wire n_1775;
wire n_1774;
wire n_1661;
wire n_1664;
wire n_1666;
wire n_1667;
wire n_1669;
wire n_1668;
wire n_1733;
wire n_1737;
wire n_1739;
wire n_1732;
wire n_1673;
wire n_1678;
wire n_1676;
wire n_1672;
wire n_1677;
wire n_1674;
wire n_1675;
wire n_1858;
wire n_1857;
wire n_1823;
wire n_1681;
wire n_1680;
wire n_1829;
wire n_1833;
wire n_1825;
wire n_1682;
wire n_1827;
wire n_1826;
wire n_1684;
wire n_1691;
wire n_1690;
wire n_1687;
wire n_1686;
wire n_1716;
wire n_1714;
wire n_1709;
wire n_1710;
wire n_1693;
wire n_1689;
wire n_1861;
wire n_1867;
wire n_1864;
wire n_1862;
wire n_1866;
wire n_1692;
wire n_1694;
wire n_1707;
wire n_1700;
wire n_1842;
wire n_1841;
wire n_1840;
wire n_1699;
wire n_1704;
wire n_1703;
wire n_1706;
wire n_1705;
wire n_1878;
wire n_1880;
wire n_1877;
wire n_1713;
wire n_1837;
wire n_1836;
wire n_1835;
wire n_1711;
wire n_1712;
wire n_1831;
wire n_1715;
wire n_1881;
wire n_1875;
wire n_1874;
wire n_1794;
wire n_1728;
wire n_1724;
wire n_1813;
wire n_1820;
wire n_1819;
wire n_1814;
wire n_1727;
wire n_1731;
wire n_1784;
wire n_1787;
wire n_1730;
wire n_1735;
wire n_1734;
wire n_1920;
wire n_1925;
wire n_1924;
wire n_1736;
wire n_1922;
wire n_1921;
wire n_1738;
wire n_1744;
wire n_1741;
wire n_1740;
wire n_1743;
wire n_2055;
wire n_2053;
wire n_2045;
wire n_1742;
wire n_2046;
wire n_1746;
wire n_1749;
wire n_1758;
wire n_1765;
wire n_1764;
wire n_1767;
wire n_1773;
wire n_1771;
wire n_1769;
wire n_1768;
wire n_2089;
wire n_2088;
wire n_2087;
wire n_1770;
wire n_1772;
wire n_2071;
wire n_2070;
wire n_2069;
wire n_1782;
wire n_1778;
wire n_1781;
wire n_1777;
wire n_1780;
wire n_1776;
wire n_2066;
wire n_2064;
wire n_2062;
wire n_1779;
wire n_2061;
wire n_2051;
wire n_2050;
wire n_2048;
wire n_1783;
wire n_2049;
wire n_1785;
wire n_1786;
wire n_1917;
wire n_1916;
wire n_1911;
wire n_1789;
wire n_1790;
wire n_1804;
wire n_1807;
wire n_1792;
wire n_1791;
wire n_1903;
wire n_1908;
wire n_1907;
wire n_1802;
wire n_1798;
wire n_1803;
wire n_1799;
wire n_1800;
wire n_1801;
wire n_1806;
wire n_1805;
wire n_1808;
wire n_1810;
wire n_1811;
wire n_2032;
wire n_2037;
wire n_1809;
wire n_2042;
wire n_2075;
wire n_2098;
wire n_2096;
wire n_2040;
wire n_2038;
wire n_2033;
wire n_1812;
wire n_1815;
wire n_1818;
wire n_1816;
wire n_1817;
wire n_2073;
wire n_2043;
wire n_1822;
wire n_1891;
wire n_1889;
wire n_1821;
wire n_1888;
wire n_1824;
wire n_2084;
wire n_2083;
wire n_2082;
wire n_1828;
wire n_1832;
wire n_1830;
wire n_1834;
wire n_1839;
wire n_1843;
wire n_1838;
wire n_8880;
wire n_1848;
wire n_1847;
wire n_8849;
wire n_1853;
wire n_1852;
wire n_1860;
wire n_1885;
wire n_1883;
wire n_1882;
wire n_1859;
wire n_1863;
wire n_1991;
wire n_1992;
wire n_1989;
wire n_1865;
wire n_1872;
wire n_1870;
wire n_1868;
wire n_1871;
wire n_1869;
wire n_2170;
wire n_2169;
wire n_2167;
wire n_1873;
wire n_1876;
wire n_1879;
wire n_8751;
wire n_1884;
wire n_1887;
wire n_2080;
wire n_1886;
wire n_2078;
wire n_2276;
wire n_2079;
wire n_1890;
wire n_1967;
wire n_1973;
wire n_1971;
wire n_1966;
wire n_1893;
wire n_1896;
wire n_1895;
wire n_2099;
wire n_2020;
wire n_2016;
wire n_1899;
wire n_1950;
wire n_1901;
wire n_1949;
wire n_1902;
wire n_1904;
wire n_1906;
wire n_1905;
wire n_1965;
wire n_1980;
wire n_1979;
wire n_1964;
wire n_1910;
wire n_1945;
wire n_1909;
wire n_1944;
wire n_1912;
wire n_1915;
wire n_1913;
wire n_1914;
wire n_1996;
wire n_1994;
wire n_1983;
wire n_1937;
wire n_1919;
wire n_1918;
wire n_1936;
wire n_2005;
wire n_2004;
wire n_2002;
wire n_2003;
wire n_1923;
wire n_2001;
wire n_1934;
wire n_1933;
wire n_1929;
wire n_1927;
wire n_1932;
wire n_1926;
wire n_1928;
wire n_2165;
wire n_2164;
wire n_2171;
wire n_1931;
wire n_1930;
wire n_1993;
wire n_1987;
wire n_1985;
wire n_1935;
wire n_1986;
wire n_1939;
wire n_1938;
wire n_1941;
wire n_2162;
wire n_2158;
wire n_1940;
wire n_2160;
wire n_2159;
wire n_2173;
wire n_1942;
wire n_1943;
wire n_1947;
wire n_1946;
wire n_2151;
wire n_2150;
wire n_2148;
wire n_2146;
wire n_1948;
wire n_2145;
wire n_1955;
wire n_1951;
wire n_1952;
wire n_1953;
wire n_1957;
wire n_1963;
wire n_2013;
wire n_2012;
wire n_1959;
wire n_1961;
wire n_1962;
wire n_1960;
wire n_2385;
wire n_2384;
wire n_2379;
wire n_1969;
wire n_1968;
wire n_2199;
wire n_2193;
wire n_2191;
wire n_1970;
wire n_2192;
wire n_1972;
wire n_1976;
wire n_1974;
wire n_7913;
wire n_1975;
wire n_2273;
wire n_2272;
wire n_2279;
wire n_1978;
wire n_1977;
wire n_2007;
wire n_1982;
wire n_1981;
wire n_2006;
wire n_1984;
wire n_1990;
wire n_1988;
wire n_1995;
wire n_1998;
wire n_1997;
wire n_2000;
wire n_2399;
wire n_2398;
wire n_2396;
wire n_1999;
wire n_2397;
wire n_8795;
wire n_2008;
wire n_2011;
wire n_2009;
wire n_2010;
wire n_2297;
wire n_2299;
wire n_2294;
wire n_2302;
wire n_2300;
wire n_2293;
wire n_2014;
wire n_2015;
wire n_2017;
wire n_2018;
wire n_2024;
wire n_2031;
wire n_2023;
wire n_2029;
wire n_2025;
wire n_2027;
wire n_2026;
wire n_2261;
wire n_2256;
wire n_2028;
wire n_2286;
wire n_2285;
wire n_2262;
wire n_2269;
wire n_2030;
wire n_2260;
wire n_2034;
wire n_2036;
wire n_2035;
wire n_2182;
wire n_2181;
wire n_2179;
wire n_2039;
wire n_2095;
wire n_2041;
wire n_2044;
wire n_2047;
wire n_2052;
wire n_2060;
wire n_2054;
wire n_2057;
wire n_2058;
wire n_2059;
wire n_2056;
wire n_2198;
wire n_2197;
wire n_2195;
wire n_2063;
wire n_2065;
wire n_2068;
wire n_2072;
wire n_2067;
wire n_8926;
wire n_2074;
wire n_2093;
wire n_2092;
wire n_2076;
wire n_2091;
wire n_2077;
wire n_2277;
wire n_2278;
wire n_2275;
wire n_2081;
wire n_2086;
wire n_2085;
wire n_2090;
wire n_2283;
wire n_2282;
wire n_2281;
wire n_2094;
wire n_2264;
wire n_2270;
wire n_2097;
wire n_2268;
wire n_2263;
wire n_2100;
wire n_2103;
wire n_2101;
wire n_2102;
wire n_2174;
wire n_2144;
wire n_2113;
wire n_2235;
wire n_2243;
wire n_2110;
wire n_2241;
wire n_2242;
wire n_2236;
wire n_2120;
wire n_2116;
wire n_2118;
wire n_2119;
wire n_2115;
wire n_2365;
wire n_2117;
wire n_2373;
wire n_2371;
wire n_2372;
wire n_2366;
wire n_2123;
wire n_2122;
wire n_2375;
wire n_2421;
wire n_2418;
wire n_2124;
wire n_2128;
wire n_2130;
wire n_2131;
wire n_2493;
wire n_2129;
wire n_2498;
wire n_2500;
wire n_2499;
wire n_2496;
wire n_2494;
wire n_2135;
wire n_2137;
wire n_2423;
wire n_2136;
wire n_2443;
wire n_2445;
wire n_2138;
wire n_2444;
wire n_2203;
wire n_2142;
wire n_2149;
wire n_2147;
wire n_2430;
wire n_2429;
wire n_2427;
wire n_2157;
wire n_2154;
wire n_2153;
wire n_2152;
wire n_2156;
wire n_2402;
wire n_2401;
wire n_2394;
wire n_2393;
wire n_2155;
wire n_2400;
wire n_2163;
wire n_2172;
wire n_2407;
wire n_2406;
wire n_2405;
wire n_2161;
wire n_2168;
wire n_2166;
wire n_2175;
wire n_2178;
wire n_2200;
wire n_2201;
wire n_2177;
wire n_2180;
wire n_2189;
wire n_2185;
wire n_2184;
wire n_2188;
wire n_2183;
wire n_2442;
wire n_2441;
wire n_2440;
wire n_2186;
wire n_2187;
wire n_2190;
wire n_2194;
wire n_2196;
wire n_2424;
wire n_2434;
wire n_2431;
wire n_2202;
wire n_2425;
wire n_2205;
wire n_2204;
wire n_2504;
wire n_2503;
wire n_2206;
wire n_2208;
wire n_2209;
wire n_2227;
wire n_2226;
wire n_2211;
wire n_2221;
wire n_2225;
wire n_2214;
wire n_2213;
wire n_2219;
wire n_2319;
wire n_2322;
wire n_2470;
wire n_2473;
wire n_2348;
wire n_2341;
wire n_2220;
wire n_2222;
wire n_2223;
wire n_2224;
wire n_2351;
wire n_2356;
wire n_2359;
wire n_2364;
wire n_2357;
wire n_2229;
wire n_2234;
wire n_2233;
wire n_2228;
wire n_2230;
wire n_2232;
wire n_2231;
wire n_2521;
wire n_2491;
wire n_2574;
wire n_2573;
wire n_2490;
wire n_2237;
wire n_2240;
wire n_2238;
wire n_2239;
wire n_2518;
wire n_2492;
wire n_2248;
wire n_2244;
wire n_2245;
wire n_2247;
wire n_2246;
wire n_2578;
wire n_2584;
wire n_2583;
wire n_2577;
wire n_2250;
wire n_2520;
wire n_2560;
wire n_2563;
wire n_2254;
wire n_2315;
wire n_2259;
wire n_2257;
wire n_2258;
wire n_2535;
wire n_2534;
wire n_2532;
wire n_2284;
wire n_2266;
wire n_2265;
wire n_2556;
wire n_2555;
wire n_2554;
wire n_2267;
wire n_2271;
wire n_2280;
wire n_2274;
wire n_2557;
wire n_2552;
wire n_2551;
wire n_2287;
wire n_2288;
wire n_2292;
wire n_2312;
wire n_2311;
wire n_2291;
wire n_2310;
wire n_2296;
wire n_2295;
wire n_2546;
wire n_2547;
wire n_2544;
wire n_2298;
wire n_8973;
wire n_2301;
wire n_2305;
wire n_2304;
wire n_2303;
wire n_2307;
wire n_2541;
wire n_2540;
wire n_2306;
wire n_2309;
wire n_2308;
wire n_2542;
wire n_2537;
wire n_2536;
wire n_2530;
wire n_2313;
wire n_2314;
wire n_2538;
wire n_2317;
wire n_2316;
wire n_2588;
wire n_2601;
wire n_2603;
wire n_2318;
wire n_2320;
wire n_2321;
wire n_2346;
wire n_2342;
wire n_2324;
wire n_2327;
wire n_2765;
wire n_2637;
wire n_2768;
wire n_2330;
wire n_2332;
wire n_2331;
wire n_2334;
wire n_2336;
wire n_2338;
wire n_2335;
wire n_2478;
wire n_2471;
wire n_2477;
wire n_2337;
wire n_2642;
wire n_2639;
wire n_2644;
wire n_2646;
wire n_2638;
wire n_2469;
wire n_2340;
wire n_2343;
wire n_2345;
wire n_2344;
wire n_2481;
wire n_2487;
wire n_2486;
wire n_2482;
wire n_2347;
wire n_2350;
wire n_2466;
wire n_2468;
wire n_2349;
wire n_2352;
wire n_2354;
wire n_2353;
wire n_2661;
wire n_2659;
wire n_2662;
wire n_2664;
wire n_2355;
wire n_2363;
wire n_2358;
wire n_2360;
wire n_2362;
wire n_2361;
wire n_2699;
wire n_2678;
wire n_2711;
wire n_2707;
wire n_2677;
wire n_2367;
wire n_2370;
wire n_2368;
wire n_2369;
wire n_2697;
wire n_2679;
wire n_2374;
wire n_2461;
wire n_2408;
wire n_2376;
wire n_2378;
wire n_2381;
wire n_2380;
wire n_2600;
wire n_2599;
wire n_2598;
wire n_2382;
wire n_2383;
wire n_2392;
wire n_2387;
wire n_2391;
wire n_2386;
wire n_2390;
wire n_2388;
wire n_2389;
wire n_2696;
wire n_2695;
wire n_2694;
wire n_2395;
wire n_8971;
wire n_2404;
wire n_2403;
wire n_2413;
wire n_2416;
wire n_2417;
wire n_2412;
wire n_2415;
wire n_2411;
wire n_2691;
wire n_2690;
wire n_2689;
wire n_2414;
wire n_2589;
wire n_2593;
wire n_2596;
wire n_2595;
wire n_2594;
wire n_2591;
wire n_2590;
wire n_2420;
wire n_2419;
wire n_2422;
wire n_2459;
wire n_2455;
wire n_2433;
wire n_2428;
wire n_2426;
wire n_2432;
wire n_2437;
wire n_2436;
wire n_2439;
wire n_2435;
wire n_2729;
wire n_2728;
wire n_2726;
wire n_2438;
wire n_8752;
wire n_2448;
wire n_2453;
wire n_2452;
wire n_2447;
wire n_2446;
wire n_2451;
wire n_2740;
wire n_2739;
wire n_2738;
wire n_2449;
wire n_2450;
wire n_2731;
wire n_2724;
wire n_2722;
wire n_2454;
wire n_2723;
wire n_2457;
wire n_2683;
wire n_2456;
wire n_2680;
wire n_2458;
wire n_2686;
wire n_2685;
wire n_2688;
wire n_2460;
wire n_2682;
wire n_2462;
wire n_2463;
wire n_2465;
wire n_2464;
wire n_2732;
wire n_2717;
wire n_2741;
wire n_2744;
wire n_2716;
wire n_2467;
wire n_2658;
wire n_2674;
wire n_2672;
wire n_2657;
wire n_2472;
wire n_2476;
wire n_2474;
wire n_2475;
wire n_2649;
wire n_2654;
wire n_2653;
wire n_2651;
wire n_2650;
wire n_2480;
wire n_2627;
wire n_2626;
wire n_2479;
wire n_2625;
wire n_2485;
wire n_2483;
wire n_2484;
wire n_2796;
wire n_2805;
wire n_2803;
wire n_2798;
wire n_2797;
wire n_2489;
wire n_2619;
wire n_2617;
wire n_2488;
wire n_2616;
wire n_2495;
wire n_2718;
wire n_2720;
wire n_2497;
wire n_2502;
wire n_2516;
wire n_2515;
wire n_2501;
wire n_2514;
wire n_2511;
wire n_2507;
wire n_2510;
wire n_2506;
wire n_2509;
wire n_2505;
wire n_2873;
wire n_2872;
wire n_2871;
wire n_2508;
wire n_2830;
wire n_2829;
wire n_2828;
wire n_2512;
wire n_2513;
wire n_2825;
wire n_2824;
wire n_2822;
wire n_2823;
wire n_2517;
wire n_2821;
wire n_2523;
wire n_2519;
wire n_2526;
wire n_2528;
wire n_2522;
wire n_2527;
wire n_2524;
wire n_2525;
wire n_2833;
wire n_2831;
wire n_2820;
wire n_2559;
wire n_2529;
wire n_2531;
wire n_2533;
wire n_8829;
wire n_2550;
wire n_2539;
wire n_2549;
wire n_2543;
wire n_2545;
wire n_2548;
wire n_2553;
wire n_8927;
wire n_2558;
wire n_2561;
wire n_2562;
wire n_2571;
wire n_2564;
wire n_2572;
wire n_2570;
wire n_2565;
wire n_2567;
wire n_2566;
wire n_2889;
wire n_2888;
wire n_2890;
wire n_2569;
wire n_2568;
wire n_2868;
wire n_2867;
wire n_2866;
wire n_2614;
wire n_2576;
wire n_2615;
wire n_2613;
wire n_2575;
wire n_2579;
wire n_2581;
wire n_2580;
wire n_2852;
wire n_2848;
wire n_2846;
wire n_2851;
wire n_2845;
wire n_2582;
wire n_2586;
wire n_2608;
wire n_2585;
wire n_2607;
wire n_2587;
wire n_2862;
wire n_2861;
wire n_2859;
wire n_2860;
wire n_2592;
wire n_2858;
wire n_2597;
wire n_8908;
wire n_2602;
wire n_2604;
wire n_2606;
wire n_2605;
wire n_2863;
wire n_2857;
wire n_2856;
wire n_2610;
wire n_2609;
wire n_2892;
wire n_2887;
wire n_2891;
wire n_2611;
wire n_2612;
wire n_2621;
wire n_2622;
wire n_2838;
wire n_2623;
wire n_2837;
wire n_2818;
wire n_2618;
wire n_2817;
wire n_2875;
wire n_2874;
wire n_2620;
wire n_2624;
wire n_2841;
wire n_2840;
wire n_2844;
wire n_2795;
wire n_2814;
wire n_2813;
wire n_2628;
wire n_2630;
wire n_2632;
wire n_2926;
wire n_2634;
wire n_2924;
wire n_2645;
wire n_2787;
wire n_2640;
wire n_2641;
wire n_2791;
wire n_2912;
wire n_2794;
wire n_2792;
wire n_2643;
wire n_2648;
wire n_2763;
wire n_2762;
wire n_2647;
wire n_2761;
wire n_2955;
wire n_2960;
wire n_2959;
wire n_2652;
wire n_2656;
wire n_2756;
wire n_2655;
wire n_2755;
wire n_2660;
wire n_2881;
wire n_2880;
wire n_2884;
wire n_2878;
wire n_2879;
wire n_2668;
wire n_2666;
wire n_2663;
wire n_2671;
wire n_2669;
wire n_2670;
wire n_2665;
wire n_2977;
wire n_2667;
wire n_2994;
wire n_2998;
wire n_2984;
wire n_2995;
wire n_2969;
wire n_2971;
wire n_2965;
wire n_2676;
wire n_2673;
wire n_2751;
wire n_2754;
wire n_2675;
wire n_2710;
wire n_2681;
wire n_2992;
wire n_2993;
wire n_2991;
wire n_2684;
wire n_3044;
wire n_3043;
wire n_3042;
wire n_2687;
wire n_2693;
wire n_2692;
wire n_2698;
wire n_2702;
wire n_2705;
wire n_2701;
wire n_2706;
wire n_2700;
wire n_2704;
wire n_3039;
wire n_3038;
wire n_3036;
wire n_3037;
wire n_2703;
wire n_3035;
wire n_2988;
wire n_2987;
wire n_2986;
wire n_2709;
wire n_2708;
wire n_2713;
wire n_2712;
wire n_2715;
wire n_3031;
wire n_3033;
wire n_3045;
wire n_2714;
wire n_3034;
wire n_2737;
wire n_2719;
wire n_2734;
wire n_2733;
wire n_2721;
wire n_2725;
wire n_2727;
wire n_2730;
wire n_8858;
wire n_2736;
wire n_3341;
wire n_3340;
wire n_3338;
wire n_2735;
wire n_3339;
wire n_2743;
wire n_2747;
wire n_2742;
wire n_2745;
wire n_2749;
wire n_2748;
wire n_2746;
wire n_3053;
wire n_3052;
wire n_3051;
wire n_3342;
wire n_3336;
wire n_3334;
wire n_2750;
wire n_3335;
wire n_2752;
wire n_2753;
wire n_2978;
wire n_2975;
wire n_2963;
wire n_2757;
wire n_2759;
wire n_3014;
wire n_2758;
wire n_3019;
wire n_3021;
wire n_3028;
wire n_3024;
wire n_3022;
wire n_2760;
wire n_3020;
wire n_2953;
wire n_3012;
wire n_3009;
wire n_2764;
wire n_2766;
wire n_2767;
wire n_2784;
wire n_2783;
wire n_2776;
wire n_2770;
wire n_3072;
wire n_3075;
wire n_2773;
wire n_2933;
wire n_2940;
wire n_2782;
wire n_2777;
wire n_2781;
wire n_2778;
wire n_2779;
wire n_2780;
wire n_2943;
wire n_2948;
wire n_2952;
wire n_3068;
wire n_3067;
wire n_2950;
wire n_2919;
wire n_2786;
wire n_2921;
wire n_2918;
wire n_2785;
wire n_2789;
wire n_2788;
wire n_3223;
wire n_3224;
wire n_3286;
wire n_2790;
wire n_2793;
wire n_2911;
wire n_2802;
wire n_2800;
wire n_2801;
wire n_2799;
wire n_3025;
wire n_3027;
wire n_3030;
wire n_3056;
wire n_3055;
wire n_2804;
wire n_2812;
wire n_2810;
wire n_2806;
wire n_2807;
wire n_2809;
wire n_3249;
wire n_3246;
wire n_3256;
wire n_2808;
wire n_2811;
wire n_3326;
wire n_3318;
wire n_3329;
wire n_2816;
wire n_2908;
wire n_2910;
wire n_2907;
wire n_2815;
wire n_2819;
wire n_2827;
wire n_2826;
wire n_8955;
wire n_2832;
wire n_2835;
wire n_2834;
wire n_3315;
wire n_3314;
wire n_3313;
wire n_2836;
wire n_2839;
wire n_3310;
wire n_3309;
wire n_3308;
wire n_2842;
wire n_2843;
wire n_2847;
wire n_2849;
wire n_3268;
wire n_2850;
wire n_3269;
wire n_3267;
wire n_2865;
wire n_2855;
wire n_2853;
wire n_2854;
wire n_8909;
wire n_2864;
wire n_2870;
wire n_2869;
wire n_8946;
wire n_2903;
wire n_2877;
wire n_2905;
wire n_2902;
wire n_2876;
wire n_2900;
wire n_2886;
wire n_2899;
wire n_3344;
wire n_3332;
wire n_3331;
wire n_2882;
wire n_2883;
wire n_2898;
wire n_2885;
wire n_2895;
wire n_2894;
wire n_2893;
wire n_3195;
wire n_3194;
wire n_3193;
wire n_2896;
wire n_2897;
wire n_3264;
wire n_3263;
wire n_3262;
wire n_2901;
wire n_2904;
wire n_3299;
wire n_3305;
wire n_3304;
wire n_2906;
wire n_2909;
wire n_3294;
wire n_3297;
wire n_3289;
wire n_2913;
wire n_2916;
wire n_3227;
wire n_3232;
wire n_2914;
wire n_3237;
wire n_3247;
wire n_2915;
wire n_3276;
wire n_3274;
wire n_3235;
wire n_2917;
wire n_3233;
wire n_2920;
wire n_3218;
wire n_3225;
wire n_3220;
wire n_2922;
wire n_2925;
wire n_2938;
wire n_2934;
wire n_2939;
wire n_2927;
wire n_3358;
wire n_3366;
wire n_3142;
wire n_3137;
wire n_2935;
wire n_2936;
wire n_2937;
wire n_3145;
wire n_3149;
wire n_3150;
wire n_3217;
wire n_3151;
wire n_2942;
wire n_3070;
wire n_3071;
wire n_2941;
wire n_3069;
wire n_2944;
wire n_2947;
wire n_2945;
wire n_2946;
wire n_3159;
wire n_3158;
wire n_3153;
wire n_2949;
wire n_3066;
wire n_2951;
wire n_2954;
wire n_2958;
wire n_2956;
wire n_2957;
wire n_3238;
wire n_3243;
wire n_3240;
wire n_3239;
wire n_2962;
wire n_3006;
wire n_3008;
wire n_2961;
wire n_3005;
wire n_2964;
wire n_2967;
wire n_2966;
wire n_3190;
wire n_3189;
wire n_3187;
wire n_2968;
wire n_3188;
wire n_2970;
wire n_2974;
wire n_2972;
wire n_2973;
wire n_3203;
wire n_3202;
wire n_3201;
wire n_2981;
wire n_2976;
wire n_2980;
wire n_2979;
wire n_2983;
wire n_3182;
wire n_3196;
wire n_3185;
wire n_3178;
wire n_3181;
wire n_2982;
wire n_2985;
wire n_2990;
wire n_2989;
wire n_2997;
wire n_3003;
wire n_2996;
wire n_3000;
wire n_3001;
wire n_3004;
wire n_3002;
wire n_2999;
wire n_3439;
wire n_3438;
wire n_3436;
wire n_3422;
wire n_3421;
wire n_3420;
wire n_3007;
wire n_3172;
wire n_3179;
wire n_3176;
wire n_3174;
wire n_3173;
wire n_3011;
wire n_3010;
wire n_3013;
wire n_3062;
wire n_3065;
wire n_3016;
wire n_3015;
wire n_3018;
wire n_3410;
wire n_3407;
wire n_3017;
wire n_3403;
wire n_3058;
wire n_3023;
wire n_3029;
wire n_3054;
wire n_3026;
wire n_3417;
wire n_3416;
wire n_3415;
wire n_3032;
wire n_3048;
wire n_3047;
wire n_3050;
wire n_3041;
wire n_3040;
wire n_3046;
wire n_3717;
wire n_3716;
wire n_3714;
wire n_3049;
wire n_3715;
wire n_3451;
wire n_3450;
wire n_3449;
wire n_3057;
wire n_3060;
wire n_3059;
wire n_3455;
wire n_3459;
wire n_3458;
wire n_3061;
wire n_3063;
wire n_3064;
wire n_3170;
wire n_3162;
wire n_3165;
wire n_3169;
wire n_3383;
wire n_3395;
wire n_3384;
wire n_3398;
wire n_3396;
wire n_3390;
wire n_3376;
wire n_3372;
wire n_3387;
wire n_3370;
wire n_3388;
wire n_3381;
wire n_3073;
wire n_3074;
wire n_3141;
wire n_3076;
wire n_3138;
wire n_3140;
wire n_3078;
wire n_3086;
wire n_3094;
wire n_3080;
wire n_3083;
wire n_3085;
wire n_3084;
wire n_3373;
wire n_3367;
wire n_3362;
wire n_3578;
wire n_3087;
wire n_3093;
wire n_3089;
wire n_3097;
wire n_3090;
wire n_3092;
wire n_3091;
wire n_3108;
wire n_3497;
wire n_3107;
wire n_3096;
wire n_3095;
wire n_3099;
wire n_3102;
wire n_3100;
wire n_3101;
wire n_4031;
wire n_4027;
wire n_3104;
wire n_3105;
wire n_3494;
wire n_3519;
wire n_3110;
wire n_3109;
wire n_4101;
wire n_4107;
wire n_4106;
wire n_3111;
wire n_3113;
wire n_3114;
wire n_3116;
wire n_3581;
wire n_3117;
wire n_3579;
wire n_3890;
wire n_3118;
wire n_3121;
wire n_3120;
wire n_3119;
wire n_3123;
wire n_3899;
wire n_3895;
wire n_3893;
wire n_3125;
wire n_3130;
wire n_3134;
wire n_3126;
wire n_3127;
wire n_4326;
wire n_4325;
wire n_4323;
wire n_3129;
wire n_3133;
wire n_3132;
wire n_3131;
wire n_3813;
wire n_3811;
wire n_3884;
wire n_3357;
wire n_3136;
wire n_3139;
wire n_3375;
wire n_3475;
wire n_3474;
wire n_3369;
wire n_3144;
wire n_3352;
wire n_3143;
wire n_3351;
wire n_3146;
wire n_3148;
wire n_3147;
wire n_3589;
wire n_3586;
wire n_3666;
wire n_3665;
wire n_3585;
wire n_3152;
wire n_3216;
wire n_3157;
wire n_3154;
wire n_3156;
wire n_3155;
wire n_3769;
wire n_3766;
wire n_3771;
wire n_3770;
wire n_3765;
wire n_3212;
wire n_3161;
wire n_3160;
wire n_3211;
wire n_3163;
wire n_3164;
wire n_3545;
wire n_3539;
wire n_3544;
wire n_3166;
wire n_3171;
wire n_3167;
wire n_3168;
wire n_3208;
wire n_3596;
wire n_3594;
wire n_3609;
wire n_3209;
wire n_3552;
wire n_3551;
wire n_3550;
wire n_3543;
wire n_3175;
wire n_3542;
wire n_3177;
wire n_3206;
wire n_3205;
wire n_3180;
wire n_3204;
wire n_3184;
wire n_3183;
wire n_3199;
wire n_3197;
wire n_3200;
wire n_3186;
wire n_3192;
wire n_3191;
wire n_3198;
wire n_3625;
wire n_3624;
wire n_3623;
wire n_3607;
wire n_3600;
wire n_3598;
wire n_3599;
wire n_3207;
wire n_3597;
wire n_3210;
wire n_3595;
wire n_3213;
wire n_3215;
wire n_3214;
wire n_3538;
wire n_3556;
wire n_3555;
wire n_3537;
wire n_3219;
wire n_3669;
wire n_3700;
wire n_3699;
wire n_3222;
wire n_3221;
wire n_3226;
wire n_3278;
wire n_3284;
wire n_3283;
wire n_3277;
wire n_3285;
wire n_3228;
wire n_3230;
wire n_3229;
wire n_3729;
wire n_3231;
wire n_3703;
wire n_3722;
wire n_3242;
wire n_3241;
wire n_3234;
wire n_3275;
wire n_3236;
wire n_3705;
wire n_3708;
wire n_3721;
wire n_3244;
wire n_3272;
wire n_3271;
wire n_3245;
wire n_3254;
wire n_3253;
wire n_3270;
wire n_3248;
wire n_3255;
wire n_3252;
wire n_3250;
wire n_3251;
wire n_3790;
wire n_3789;
wire n_3788;
wire n_3257;
wire n_3261;
wire n_3259;
wire n_3258;
wire n_3605;
wire n_3604;
wire n_3602;
wire n_3603;
wire n_3260;
wire n_3601;
wire n_3266;
wire n_3265;
wire n_3791;
wire n_3786;
wire n_3785;
wire n_3273;
wire n_3787;
wire n_3775;
wire n_3777;
wire n_3780;
wire n_3280;
wire n_3279;
wire n_3282;
wire n_3677;
wire n_3678;
wire n_3281;
wire n_3671;
wire n_3287;
wire n_3348;
wire n_3350;
wire n_3288;
wire n_3292;
wire n_3290;
wire n_3291;
wire n_3442;
wire n_3430;
wire n_3429;
wire n_3433;
wire n_3431;
wire n_3293;
wire n_3296;
wire n_3295;
wire n_3298;
wire n_3317;
wire n_3303;
wire n_3301;
wire n_3300;
wire n_3727;
wire n_3726;
wire n_3725;
wire n_3302;
wire n_3307;
wire n_3306;
wire n_3316;
wire n_3312;
wire n_3311;
wire n_3320;
wire n_3319;
wire n_3322;
wire n_3432;
wire n_3321;
wire n_3325;
wire n_3323;
wire n_3324;
wire n_3434;
wire n_3441;
wire n_3328;
wire n_3327;
wire n_3330;
wire n_3345;
wire n_3347;
wire n_3333;
wire n_3337;
wire n_3343;
wire n_3346;
wire n_3719;
wire n_3712;
wire n_3710;
wire n_3402;
wire n_3426;
wire n_3349;
wire n_3428;
wire n_3453;
wire n_3423;
wire n_3401;
wire n_3427;
wire n_3353;
wire n_3356;
wire n_3354;
wire n_3355;
wire n_3750;
wire n_3753;
wire n_3584;
wire n_3360;
wire n_3359;
wire n_3361;
wire n_3365;
wire n_3363;
wire n_3364;
wire n_3580;
wire n_3583;
wire n_3577;
wire n_3576;
wire n_3489;
wire n_3368;
wire n_3371;
wire n_3379;
wire n_3377;
wire n_3374;
wire n_3488;
wire n_3473;
wire n_3378;
wire n_3380;
wire n_3761;
wire n_3762;
wire n_3755;
wire n_3386;
wire n_3382;
wire n_3400;
wire n_3385;
wire n_3468;
wire n_3466;
wire n_3469;
wire n_3472;
wire n_3389;
wire n_3391;
wire n_3394;
wire n_3392;
wire n_3393;
wire n_3628;
wire n_3626;
wire n_3592;
wire n_3397;
wire n_3467;
wire n_3399;
wire n_3405;
wire n_3404;
wire n_3620;
wire n_3619;
wire n_3617;
wire n_3618;
wire n_3406;
wire n_3616;
wire n_3409;
wire n_3408;
wire n_3411;
wire n_3413;
wire n_3414;
wire n_3412;
wire n_3697;
wire n_3696;
wire n_3694;
wire n_3419;
wire n_3418;
wire n_3424;
wire n_3425;
wire n_3443;
wire n_3448;
wire n_3435;
wire n_3437;
wire n_3440;
wire n_3446;
wire n_3444;
wire n_3445;
wire n_3932;
wire n_3931;
wire n_3933;
wire n_3447;
wire n_3452;
wire n_3454;
wire n_3456;
wire n_3457;
wire n_3464;
wire n_3461;
wire n_3462;
wire n_3465;
wire n_3460;
wire n_3463;
wire n_3966;
wire n_3965;
wire n_3963;
wire n_3945;
wire n_3942;
wire n_3944;
wire n_3638;
wire n_3641;
wire n_3653;
wire n_3470;
wire n_3471;
wire n_3534;
wire n_3533;
wire n_3529;
wire n_3484;
wire n_3477;
wire n_3487;
wire n_3483;
wire n_3476;
wire n_3479;
wire n_3478;
wire n_3481;
wire n_3508;
wire n_3506;
wire n_3480;
wire n_3482;
wire n_3503;
wire n_3501;
wire n_3485;
wire n_3486;
wire n_3526;
wire n_3525;
wire n_3520;
wire n_3490;
wire n_3493;
wire n_3491;
wire n_3492;
wire n_3495;
wire n_3518;
wire n_3499;
wire n_3496;
wire n_4040;
wire n_4045;
wire n_4044;
wire n_3498;
wire n_3517;
wire n_3516;
wire n_3500;
wire n_3502;
wire n_3504;
wire n_4139;
wire n_4134;
wire n_4118;
wire n_3505;
wire n_4113;
wire n_4114;
wire n_3507;
wire n_3636;
wire n_3511;
wire n_3642;
wire n_3590;
wire n_3510;
wire n_3509;
wire n_3515;
wire n_3660;
wire n_3643;
wire n_3591;
wire n_3513;
wire n_3512;
wire n_4181;
wire n_4180;
wire n_4174;
wire n_3514;
wire n_4176;
wire n_4175;
wire n_4041;
wire n_3524;
wire n_3521;
wire n_3523;
wire n_3522;
wire n_3817;
wire n_3823;
wire n_3824;
wire n_3816;
wire n_3571;
wire n_3528;
wire n_3527;
wire n_3570;
wire n_3530;
wire n_3532;
wire n_3531;
wire n_4070;
wire n_4057;
wire n_4056;
wire n_3536;
wire n_3569;
wire n_3567;
wire n_3535;
wire n_3566;
wire n_3541;
wire n_3540;
wire n_3546;
wire n_3548;
wire n_3549;
wire n_3547;
wire n_4131;
wire n_4130;
wire n_4129;
wire n_3553;
wire n_3564;
wire n_3559;
wire n_3558;
wire n_3563;
wire n_3562;
wire n_3557;
wire n_4126;
wire n_4125;
wire n_4124;
wire n_3560;
wire n_3561;
wire n_4127;
wire n_4082;
wire n_4081;
wire n_4079;
wire n_4078;
wire n_4080;
wire n_3565;
wire n_4084;
wire n_4087;
wire n_3568;
wire n_4112;
wire n_3573;
wire n_3572;
wire n_4058;
wire n_4053;
wire n_4048;
wire n_3574;
wire n_3575;
wire n_3807;
wire n_3582;
wire n_3664;
wire n_3588;
wire n_3587;
wire n_3593;
wire n_3615;
wire n_3612;
wire n_3611;
wire n_3606;
wire n_3608;
wire n_3614;
wire n_3610;
wire n_4161;
wire n_4160;
wire n_4159;
wire n_3613;
wire n_3622;
wire n_3621;
wire n_3627;
wire n_3631;
wire n_3634;
wire n_3630;
wire n_3635;
wire n_3629;
wire n_3633;
wire n_4156;
wire n_4154;
wire n_4155;
wire n_3632;
wire n_4151;
wire n_4150;
wire n_4149;
wire n_3637;
wire n_3662;
wire n_3661;
wire n_3640;
wire n_3639;
wire n_3646;
wire n_3645;
wire n_3651;
wire n_3648;
wire n_3644;
wire n_3652;
wire n_4355;
wire n_4354;
wire n_4352;
wire n_4353;
wire n_3647;
wire n_4351;
wire n_3649;
wire n_3650;
wire n_3655;
wire n_4363;
wire n_4364;
wire n_4362;
wire n_3659;
wire n_3690;
wire n_3654;
wire n_3656;
wire n_3657;
wire n_3658;
wire n_3689;
wire n_3692;
wire n_4136;
wire n_4147;
wire n_4142;
wire n_4141;
wire n_4146;
wire n_3663;
wire n_4148;
wire n_4153;
wire n_3746;
wire n_3668;
wire n_3748;
wire n_3667;
wire n_3745;
wire n_3670;
wire n_3673;
wire n_3672;
wire n_3960;
wire n_3675;
wire n_3959;
wire n_3674;
wire n_3676;
wire n_3687;
wire n_3680;
wire n_3686;
wire n_3681;
wire n_3685;
wire n_3679;
wire n_3939;
wire n_3683;
wire n_3938;
wire n_3682;
wire n_3684;
wire n_3688;
wire n_3691;
wire n_3693;
wire n_3695;
wire n_3698;
wire n_3741;
wire n_3702;
wire n_3743;
wire n_3740;
wire n_3701;
wire n_3704;
wire n_3732;
wire n_3738;
wire n_3736;
wire n_3731;
wire n_3706;
wire n_3707;
wire n_3723;
wire n_3728;
wire n_3711;
wire n_3709;
wire n_3713;
wire n_3720;
wire n_3724;
wire n_3730;
wire n_3735;
wire n_3843;
wire n_3842;
wire n_3841;
wire n_3733;
wire n_3734;
wire n_3934;
wire n_3737;
wire n_3929;
wire n_3930;
wire n_3739;
wire n_3928;
wire n_3742;
wire n_3950;
wire n_3956;
wire n_3955;
wire n_3744;
wire n_3747;
wire n_3913;
wire n_3749;
wire n_3919;
wire n_3910;
wire n_3917;
wire n_3916;
wire n_3752;
wire n_3751;
wire n_3754;
wire n_3803;
wire n_3806;
wire n_3760;
wire n_3757;
wire n_3756;
wire n_3759;
wire n_3867;
wire n_3861;
wire n_3758;
wire n_3862;
wire n_3764;
wire n_3797;
wire n_3801;
wire n_3763;
wire n_3796;
wire n_3767;
wire n_3768;
wire n_3926;
wire n_3924;
wire n_3922;
wire n_3773;
wire n_3794;
wire n_3793;
wire n_3772;
wire n_3792;
wire n_3774;
wire n_3776;
wire n_4086;
wire n_4085;
wire n_3779;
wire n_3778;
wire n_3781;
wire n_3783;
wire n_3784;
wire n_3782;
wire n_3854;
wire n_3853;
wire n_3852;
wire n_3835;
wire n_3839;
wire n_3845;
wire n_3838;
wire n_3795;
wire n_3844;
wire n_3827;
wire n_3799;
wire n_3798;
wire n_3830;
wire n_3800;
wire n_3831;
wire n_3832;
wire n_3802;
wire n_3905;
wire n_3804;
wire n_3898;
wire n_3909;
wire n_3805;
wire n_3973;
wire n_3974;
wire n_3911;
wire n_3908;
wire n_3906;
wire n_3808;
wire n_3810;
wire n_3814;
wire n_3809;
wire n_3883;
wire n_3878;
wire n_3812;
wire n_3815;
wire n_3821;
wire n_3818;
wire n_3820;
wire n_4785;
wire n_3819;
wire n_4782;
wire n_4784;
wire n_3822;
wire n_3826;
wire n_3860;
wire n_3825;
wire n_3859;
wire n_3828;
wire n_3829;
wire n_4915;
wire n_4913;
wire n_4914;
wire n_3834;
wire n_3856;
wire n_3858;
wire n_3833;
wire n_3837;
wire n_3836;
wire n_3846;
wire n_3851;
wire n_3840;
wire n_3848;
wire n_3847;
wire n_4920;
wire n_4919;
wire n_4918;
wire n_3849;
wire n_3850;
wire n_3855;
wire n_3857;
wire n_4909;
wire n_4908;
wire n_4907;
wire n_3874;
wire n_3870;
wire n_3873;
wire n_3869;
wire n_3864;
wire n_3863;
wire n_4779;
wire n_4773;
wire n_4772;
wire n_3865;
wire n_3866;
wire n_3872;
wire n_3868;
wire n_4901;
wire n_4898;
wire n_4900;
wire n_3871;
wire n_4899;
wire n_4792;
wire n_4791;
wire n_3876;
wire n_3875;
wire n_3877;
wire n_4794;
wire n_4797;
wire n_3880;
wire n_3879;
wire n_4838;
wire n_4837;
wire n_4822;
wire n_3881;
wire n_3882;
wire n_3886;
wire n_3885;
wire n_4761;
wire n_3888;
wire n_4780;
wire n_3887;
wire n_3889;
wire n_4803;
wire n_4801;
wire n_4781;
wire n_3891;
wire n_3894;
wire n_3892;
wire n_3975;
wire n_3897;
wire n_3896;
wire n_3900;
wire n_3903;
wire n_3904;
wire n_3901;
wire n_3902;
wire n_4336;
wire n_4335;
wire n_4329;
wire n_3907;
wire n_4347;
wire n_4367;
wire n_4368;
wire n_3971;
wire n_3949;
wire n_3920;
wire n_3970;
wire n_3912;
wire n_3918;
wire n_3915;
wire n_3914;
wire n_4359;
wire n_4358;
wire n_4350;
wire n_4349;
wire n_4357;
wire n_4360;
wire n_3921;
wire n_3923;
wire n_4796;
wire n_4795;
wire n_3925;
wire n_3937;
wire n_3927;
wire n_3936;
wire n_3935;
wire n_3940;
wire n_3948;
wire n_3941;
wire n_3943;
wire n_3946;
wire n_3947;
wire n_3954;
wire n_3952;
wire n_3951;
wire n_4778;
wire n_4777;
wire n_4775;
wire n_4776;
wire n_3953;
wire n_4774;
wire n_3958;
wire n_3957;
wire n_3969;
wire n_3961;
wire n_3968;
wire n_3962;
wire n_3964;
wire n_3967;
wire n_3972;
wire n_4767;
wire n_4770;
wire n_4763;
wire n_3976;
wire n_3979;
wire n_3977;
wire n_3978;
wire n_4169;
wire n_4171;
wire n_4110;
wire n_3990;
wire n_3982;
wire n_3983;
wire n_3989;
wire n_3985;
wire n_4224;
wire n_4226;
wire n_4228;
wire n_3988;
wire n_3987;
wire n_4230;
wire n_4259;
wire n_4231;
wire n_4235;
wire n_3991;
wire n_3997;
wire n_3994;
wire n_4410;
wire n_3995;
wire n_4284;
wire n_4412;
wire n_4612;
wire n_4613;
wire n_4413;
wire n_4411;
wire n_4213;
wire n_3999;
wire n_4002;
wire n_4005;
wire n_4303;
wire n_4003;
wire n_4004;
wire n_4309;
wire n_4312;
wire n_4403;
wire n_4408;
wire n_4310;
wire n_4304;
wire n_4009;
wire n_4014;
wire n_4012;
wire n_4008;
wire n_4013;
wire n_4643;
wire n_4010;
wire n_4011;
wire n_4663;
wire n_5010;
wire n_4666;
wire n_4867;
wire n_4664;
wire n_4644;
wire n_4017;
wire n_4020;
wire n_4018;
wire n_4019;
wire n_4866;
wire n_4667;
wire n_4023;
wire n_4208;
wire n_4099;
wire n_4204;
wire n_4205;
wire n_4028;
wire n_4030;
wire n_4029;
wire n_4734;
wire n_4758;
wire n_4756;
wire n_4733;
wire n_4033;
wire n_4032;
wire n_4036;
wire n_4035;
wire n_4039;
wire n_4038;
wire n_4890;
wire n_4889;
wire n_4037;
wire n_4871;
wire n_4042;
wire n_4043;
wire n_4921;
wire n_4893;
wire n_4894;
wire n_4904;
wire n_4092;
wire n_4047;
wire n_4046;
wire n_4091;
wire n_4050;
wire n_4049;
wire n_4896;
wire n_4895;
wire n_4051;
wire n_4052;
wire n_4055;
wire n_4054;
wire n_4059;
wire n_4065;
wire n_4077;
wire n_4072;
wire n_4069;
wire n_4064;
wire n_4060;
wire n_4061;
wire n_4454;
wire n_4453;
wire n_4446;
wire n_4062;
wire n_4063;
wire n_4455;
wire n_4066;
wire n_4068;
wire n_4067;
wire n_4451;
wire n_4450;
wire n_4448;
wire n_4076;
wire n_4071;
wire n_4073;
wire n_4075;
wire n_4074;
wire n_4459;
wire n_4458;
wire n_4457;
wire n_4083;
wire n_4090;
wire n_4089;
wire n_4088;
wire n_4095;
wire n_4093;
wire n_4094;
wire n_4441;
wire n_4438;
wire n_4436;
wire n_5781;
wire n_4435;
wire n_4437;
wire n_4096;
wire n_4203;
wire n_4098;
wire n_4100;
wire n_4102;
wire n_4105;
wire n_4103;
wire n_4104;
wire n_4461;
wire n_4462;
wire n_4434;
wire n_4196;
wire n_4109;
wire n_4108;
wire n_4195;
wire n_4133;
wire n_4111;
wire n_4117;
wire n_4116;
wire n_4115;
wire n_4119;
wire n_4123;
wire n_4121;
wire n_4120;
wire n_4490;
wire n_4489;
wire n_4487;
wire n_4122;
wire n_4128;
wire n_4132;
wire n_4137;
wire n_4135;
wire n_4144;
wire n_4145;
wire n_4138;
wire n_4166;
wire n_4164;
wire n_4163;
wire n_4140;
wire n_4143;
wire n_4708;
wire n_4710;
wire n_4707;
wire n_4152;
wire n_4158;
wire n_4157;
wire n_4162;
wire n_4165;
wire n_4484;
wire n_4167;
wire n_4483;
wire n_4168;
wire n_4170;
wire n_4173;
wire n_4190;
wire n_4193;
wire n_4172;
wire n_4504;
wire n_4503;
wire n_4502;
wire n_4178;
wire n_4179;
wire n_4177;
wire n_4184;
wire n_4188;
wire n_4187;
wire n_4183;
wire n_4182;
wire n_4186;
wire n_4690;
wire n_4689;
wire n_4687;
wire n_4185;
wire n_4688;
wire n_4711;
wire n_4705;
wire n_4703;
wire n_4704;
wire n_4189;
wire n_4702;
wire n_4192;
wire n_4481;
wire n_4191;
wire n_4478;
wire n_4480;
wire n_4194;
wire n_4197;
wire n_4200;
wire n_4198;
wire n_4199;
wire n_4201;
wire n_4493;
wire n_4477;
wire n_4202;
wire n_4508;
wire n_4507;
wire n_4494;
wire n_4870;
wire n_4939;
wire n_4207;
wire n_4206;
wire n_4948;
wire n_4938;
wire n_4936;
wire n_4942;
wire n_4210;
wire n_4212;
wire n_4211;
wire n_4422;
wire n_4429;
wire n_4428;
wire n_4424;
wire n_4423;
wire n_4286;
wire n_4215;
wire n_4294;
wire n_4293;
wire n_4287;
wire n_4218;
wire n_4219;
wire n_4253;
wire n_4256;
wire n_4283;
wire n_4221;
wire n_4223;
wire n_4225;
wire n_4241;
wire n_4232;
wire n_4245;
wire n_4227;
wire n_5730;
wire n_5728;
wire n_5737;
wire n_5732;
wire n_5727;
wire n_4255;
wire n_4257;
wire n_4234;
wire n_4233;
wire n_4236;
wire n_4246;
wire n_4243;
wire n_4275;
wire n_4237;
wire n_4240;
wire n_4238;
wire n_4239;
wire n_5995;
wire n_5740;
wire n_5994;
wire n_5733;
wire n_4242;
wire n_4244;
wire n_4281;
wire n_4271;
wire n_4268;
wire n_4251;
wire n_4247;
wire n_4250;
wire n_4248;
wire n_4249;
wire n_6382;
wire n_6381;
wire n_6094;
wire n_4254;
wire n_4265;
wire n_4261;
wire n_5015;
wire n_4258;
wire n_4262;
wire n_4264;
wire n_4260;
wire n_4615;
wire n_5019;
wire n_5741;
wire n_4263;
wire n_5746;
wire n_5748;
wire n_5747;
wire n_5743;
wire n_5742;
wire n_4266;
wire n_4270;
wire n_4267;
wire n_4269;
wire n_4606;
wire n_4416;
wire n_4603;
wire n_4273;
wire n_4272;
wire n_4280;
wire n_4276;
wire n_4274;
wire n_6096;
wire n_6124;
wire n_6123;
wire n_4278;
wire n_4279;
wire n_4277;
wire n_5032;
wire n_5035;
wire n_5028;
wire n_6097;
wire n_4282;
wire n_4285;
wire n_4288;
wire n_4292;
wire n_4289;
wire n_4290;
wire n_4291;
wire n_4617;
wire n_4633;
wire n_4636;
wire n_4642;
wire n_4634;
wire n_4296;
wire n_4302;
wire n_4301;
wire n_4295;
wire n_4298;
wire n_4297;
wire n_4571;
wire n_4419;
wire n_4574;
wire n_4299;
wire n_4300;
wire n_4305;
wire n_4308;
wire n_4306;
wire n_4307;
wire n_4520;
wire n_4522;
wire n_4421;
wire n_4311;
wire n_4402;
wire n_4314;
wire n_4318;
wire n_4317;
wire n_4433;
wire n_4387;
wire n_4322;
wire n_4321;
wire n_4386;
wire n_4324;
wire n_4547;
wire n_4554;
wire n_4553;
wire n_4328;
wire n_4378;
wire n_4327;
wire n_4377;
wire n_4330;
wire n_4332;
wire n_4331;
wire n_4334;
wire n_4500;
wire n_4333;
wire n_4495;
wire n_4499;
wire n_4346;
wire n_4339;
wire n_4338;
wire n_4345;
wire n_4337;
wire n_4692;
wire n_4341;
wire n_4685;
wire n_4340;
wire n_4344;
wire n_4343;
wire n_4342;
wire n_4698;
wire n_4695;
wire n_4697;
wire n_4348;
wire n_4356;
wire n_4361;
wire n_4365;
wire n_4371;
wire n_4375;
wire n_4374;
wire n_4370;
wire n_4369;
wire n_4373;
wire n_4696;
wire n_4372;
wire n_4694;
wire n_4819;
wire n_4818;
wire n_4816;
wire n_4376;
wire n_4817;
wire n_4379;
wire n_4382;
wire n_4380;
wire n_4381;
wire n_4713;
wire n_4383;
wire n_4684;
wire n_4384;
wire n_4716;
wire n_4715;
wire n_4385;
wire n_4802;
wire n_4805;
wire n_4814;
wire n_4388;
wire n_4391;
wire n_4389;
wire n_4390;
wire n_4539;
wire n_4537;
wire n_4533;
wire n_4393;
wire n_4401;
wire n_4396;
wire n_4398;
wire n_4399;
wire n_4395;
wire n_4400;
wire n_4397;
wire n_4589;
wire n_4588;
wire n_4586;
wire n_4530;
wire n_4529;
wire n_4525;
wire n_4577;
wire n_4404;
wire n_4405;
wire n_4581;
wire n_4585;
wire n_4598;
wire n_4406;
wire n_4407;
wire n_5948;
wire n_5924;
wire n_5958;
wire n_5954;
wire n_4583;
wire n_4409;
wire n_4414;
wire n_4611;
wire n_4417;
wire n_4415;
wire n_4418;
wire n_4602;
wire n_4420;
wire n_4427;
wire n_5058;
wire n_5056;
wire n_5052;
wire n_4425;
wire n_4426;
wire n_4515;
wire n_4431;
wire n_4430;
wire n_4514;
wire n_5782;
wire n_5783;
wire n_5780;
wire n_4440;
wire n_4439;
wire n_4444;
wire n_4442;
wire n_4445;
wire n_4443;
wire n_5789;
wire n_5788;
wire n_5787;
wire n_4447;
wire n_4449;
wire n_4452;
wire n_4456;
wire n_4460;
wire n_4465;
wire n_4470;
wire n_4464;
wire n_4469;
wire n_4463;
wire n_4468;
wire n_5085;
wire n_5077;
wire n_5078;
wire n_4467;
wire n_4466;
wire n_5086;
wire n_5784;
wire n_5777;
wire n_5778;
wire n_4471;
wire n_4472;
wire n_4476;
wire n_4513;
wire n_4511;
wire n_4510;
wire n_4475;
wire n_4506;
wire n_4479;
wire n_5811;
wire n_5812;
wire n_5810;
wire n_4482;
wire n_4485;
wire n_4492;
wire n_4486;
wire n_4488;
wire n_4491;
wire n_4498;
wire n_4496;
wire n_4497;
wire n_5938;
wire n_5937;
wire n_5936;
wire n_4501;
wire n_4505;
wire n_5807;
wire n_5806;
wire n_5805;
wire n_4509;
wire n_5801;
wire n_4512;
wire n_5768;
wire n_5771;
wire n_5764;
wire n_4517;
wire n_4516;
wire n_5762;
wire n_5791;
wire n_5790;
wire n_4518;
wire n_4519;
wire n_4521;
wire n_4524;
wire n_4568;
wire n_4567;
wire n_4523;
wire n_4526;
wire n_4528;
wire n_4527;
wire n_5828;
wire n_5826;
wire n_5829;
wire n_5823;
wire n_5825;
wire n_4532;
wire n_4566;
wire n_4564;
wire n_4531;
wire n_4563;
wire n_4534;
wire n_4536;
wire n_4535;
wire n_5798;
wire n_5803;
wire n_5794;
wire n_4538;
wire n_4544;
wire n_4541;
wire n_4545;
wire n_4540;
wire n_4542;
wire n_4543;
wire n_5838;
wire n_5836;
wire n_5832;
wire n_4552;
wire n_4546;
wire n_4548;
wire n_4550;
wire n_4549;
wire n_5944;
wire n_4551;
wire n_5943;
wire n_5945;
wire n_5942;
wire n_4561;
wire n_4557;
wire n_4556;
wire n_4560;
wire n_4559;
wire n_4555;
wire n_5933;
wire n_5932;
wire n_5930;
wire n_5931;
wire n_5929;
wire n_4558;
wire n_5935;
wire n_5893;
wire n_5892;
wire n_5890;
wire n_5891;
wire n_4562;
wire n_5889;
wire n_4565;
wire n_5939;
wire n_5927;
wire n_5925;
wire n_5926;
wire n_5760;
wire n_5818;
wire n_5821;
wire n_4569;
wire n_4570;
wire n_4573;
wire n_4572;
wire n_4575;
wire n_4599;
wire n_4601;
wire n_4576;
wire n_4579;
wire n_4578;
wire n_5865;
wire n_5871;
wire n_5870;
wire n_4580;
wire n_4582;
wire n_4597;
wire n_4596;
wire n_4584;
wire n_4587;
wire n_4672;
wire n_4679;
wire n_4721;
wire n_4852;
wire n_4591;
wire n_4595;
wire n_4593;
wire n_4592;
wire n_4590;
wire n_4862;
wire n_4855;
wire n_4594;
wire n_5878;
wire n_5881;
wire n_5874;
wire n_5923;
wire n_5752;
wire n_5755;
wire n_4600;
wire n_5854;
wire n_5759;
wire n_5757;
wire n_5756;
wire n_5753;
wire n_4604;
wire n_4605;
wire n_4607;
wire n_4625;
wire n_4608;
wire n_4609;
wire n_4628;
wire n_4619;
wire n_6127;
wire n_6151;
wire n_6144;
wire n_4610;
wire n_5014;
wire n_4614;
wire n_4616;
wire n_4618;
wire n_4621;
wire n_4620;
wire n_4622;
wire n_4624;
wire n_4623;
wire n_5914;
wire n_5863;
wire n_5917;
wire n_5864;
wire n_5916;
wire n_5915;
wire n_4626;
wire n_4627;
wire n_4629;
wire n_4652;
wire n_4630;
wire n_4632;
wire n_4654;
wire n_4649;
wire n_4631;
wire n_6194;
wire n_6147;
wire n_6146;
wire n_4641;
wire n_4635;
wire n_4638;
wire n_4637;
wire n_5042;
wire n_5047;
wire n_5046;
wire n_4639;
wire n_4640;
wire n_4645;
wire n_4648;
wire n_4647;
wire n_4646;
wire n_4959;
wire n_4651;
wire n_4650;
wire n_4955;
wire n_4961;
wire n_4660;
wire n_4653;
wire n_4659;
wire n_4656;
wire n_4657;
wire n_4658;
wire n_4655;
wire n_6430;
wire n_6431;
wire n_6426;
wire n_6158;
wire n_6154;
wire n_6155;
wire n_4661;
wire n_4662;
wire n_4665;
wire n_5009;
wire n_4668;
wire n_4675;
wire n_4671;
wire n_4674;
wire n_4673;
wire n_4680;
wire n_4683;
wire n_4720;
wire n_4678;
wire n_4676;
wire n_4743;
wire n_4677;
wire n_4749;
wire n_4736;
wire n_4681;
wire n_4682;
wire n_4754;
wire n_4750;
wire n_4739;
wire n_4738;
wire n_4719;
wire n_4714;
wire n_4701;
wire n_4693;
wire n_4686;
wire n_4691;
wire n_4700;
wire n_4699;
wire n_4706;
wire n_4709;
wire n_4712;
wire n_5906;
wire n_5905;
wire n_5904;
wire n_4717;
wire n_4718;
wire n_4808;
wire n_4722;
wire n_4724;
wire n_5928;
wire n_4723;
wire n_4725;
wire n_4726;
wire n_4727;
wire n_5940;
wire n_4729;
wire n_4732;
wire n_4848;
wire n_4731;
wire n_4737;
wire n_4735;
wire n_4742;
wire n_5900;
wire n_5899;
wire n_5898;
wire n_4740;
wire n_4741;
wire n_4744;
wire n_4827;
wire n_4748;
wire n_4745;
wire n_4752;
wire n_4746;
wire n_4747;
wire n_5984;
wire n_5982;
wire n_5983;
wire n_4826;
wire n_4836;
wire n_4751;
wire n_4753;
wire n_4755;
wire n_4835;
wire n_4760;
wire n_4757;
wire n_4820;
wire n_4759;
wire n_4800;
wire n_4762;
wire n_4765;
wire n_4764;
wire n_4812;
wire n_4811;
wire n_4810;
wire n_4766;
wire n_4768;
wire n_4769;
wire n_4771;
wire n_4783;
wire n_4831;
wire n_4832;
wire n_4830;
wire n_4786;
wire n_4790;
wire n_4788;
wire n_4787;
wire n_4987;
wire n_4986;
wire n_4984;
wire n_4789;
wire n_4985;
wire n_4793;
wire n_4799;
wire n_4798;
wire n_4813;
wire n_4804;
wire n_4806;
wire n_4809;
wire n_4807;
wire n_4815;
wire n_4821;
wire n_4824;
wire n_4823;
wire n_4825;
wire n_4829;
wire n_4828;
wire n_4834;
wire n_4833;
wire n_4841;
wire n_4846;
wire n_4845;
wire n_4840;
wire n_4844;
wire n_4839;
wire n_4996;
wire n_4994;
wire n_4995;
wire n_4842;
wire n_4843;
wire n_4981;
wire n_4980;
wire n_4977;
wire n_4847;
wire n_4979;
wire n_4849;
wire n_4851;
wire n_4850;
wire n_4861;
wire n_4853;
wire n_4854;
wire n_4856;
wire n_4879;
wire n_4857;
wire n_4858;
wire n_4880;
wire n_4873;
wire n_5979;
wire n_5978;
wire n_5977;
wire n_4860;
wire n_4859;
wire n_5980;
wire n_4863;
wire n_5888;
wire n_5886;
wire n_4865;
wire n_4864;
wire n_5887;
wire n_5895;
wire n_4869;
wire n_4953;
wire n_4952;
wire n_4951;
wire n_4868;
wire n_4937;
wire n_4935;
wire n_4888;
wire n_4874;
wire n_4872;
wire n_4876;
wire n_4875;
wire n_4878;
wire n_6180;
wire n_6179;
wire n_6178;
wire n_4877;
wire n_4882;
wire n_4887;
wire n_4881;
wire n_4884;
wire n_4883;
wire n_6451;
wire n_6450;
wire n_6449;
wire n_4885;
wire n_4886;
wire n_4892;
wire n_4933;
wire n_4932;
wire n_4891;
wire n_4931;
wire n_4929;
wire n_4928;
wire n_4924;
wire n_4923;
wire n_4912;
wire n_4906;
wire n_4897;
wire n_4903;
wire n_4902;
wire n_4911;
wire n_4905;
wire n_4910;
wire n_4917;
wire n_4916;
wire n_4927;
wire n_4922;
wire n_5090;
wire n_5088;
wire n_5089;
wire n_4925;
wire n_4926;
wire n_5083;
wire n_5080;
wire n_5082;
wire n_4930;
wire n_5081;
wire n_4991;
wire n_4974;
wire n_4975;
wire n_4934;
wire n_4970;
wire n_4940;
wire n_4946;
wire n_4947;
wire n_4941;
wire n_4943;
wire n_5071;
wire n_5066;
wire n_4945;
wire n_4944;
wire n_5072;
wire n_5076;
wire n_4950;
wire n_4972;
wire n_4949;
wire n_4964;
wire n_4968;
wire n_4971;
wire n_4954;
wire n_4956;
wire n_4958;
wire n_4957;
wire n_5965;
wire n_5963;
wire n_5970;
wire n_5966;
wire n_5006;
wire n_5005;
wire n_4963;
wire n_4960;
wire n_4962;
wire n_5004;
wire n_4965;
wire n_4967;
wire n_4966;
wire n_6446;
wire n_6445;
wire n_6444;
wire n_4969;
wire n_5000;
wire n_4973;
wire n_4993;
wire n_4976;
wire n_4978;
wire n_4982;
wire n_4990;
wire n_4983;
wire n_4989;
wire n_4988;
wire n_4992;
wire n_4999;
wire n_4997;
wire n_4998;
wire n_5002;
wire n_5001;
wire n_6182;
wire n_6176;
wire n_6175;
wire n_5003;
wire n_6169;
wire n_6170;
wire n_6165;
wire n_6161;
wire n_5007;
wire n_5008;
wire n_5011;
wire n_5013;
wire n_5012;
wire n_5051;
wire n_5093;
wire n_5092;
wire n_5050;
wire n_5016;
wire n_5027;
wire n_5022;
wire n_5021;
wire n_5018;
wire n_5017;
wire n_5020;
wire n_5026;
wire n_5025;
wire n_5860;
wire n_5859;
wire n_5751;
wire n_5023;
wire n_5024;
wire n_5029;
wire n_5031;
wire n_5030;
wire n_6393;
wire n_6392;
wire n_6456;
wire n_5034;
wire n_5033;
wire n_5036;
wire n_5041;
wire n_5037;
wire n_5039;
wire n_5038;
wire n_6548;
wire n_6551;
wire n_6552;
wire n_5040;
wire n_5043;
wire n_5045;
wire n_5044;
wire n_6398;
wire n_6403;
wire n_6402;
wire n_6401;
wire n_6399;
wire n_5104;
wire n_5049;
wire n_5048;
wire n_5103;
wire n_5054;
wire n_5053;
wire n_6441;
wire n_6440;
wire n_6439;
wire n_5055;
wire n_5057;
wire n_5065;
wire n_5062;
wire n_5059;
wire n_5064;
wire n_5061;
wire n_6410;
wire n_5060;
wire n_6407;
wire n_6409;
wire n_5063;
wire n_5070;
wire n_5068;
wire n_5067;
wire n_6414;
wire n_6413;
wire n_6412;
wire n_5069;
wire n_5074;
wire n_5073;
wire n_6475;
wire n_6474;
wire n_6472;
wire n_5075;
wire n_6473;
wire n_5087;
wire n_5079;
wire n_5084;
wire n_5091;
wire n_5099;
wire n_5095;
wire n_5101;
wire n_5096;
wire n_5098;
wire n_5094;
wire n_6486;
wire n_6462;
wire n_6466;
wire n_5097;
wire n_6465;
wire n_5100;
wire n_6406;
wire n_6419;
wire n_6417;
wire n_5102;
wire n_5106;
wire n_5105;
wire n_6493;
wire n_6459;
wire n_6460;
wire n_5107;
wire n_5109;
wire n_5111;
wire n_5113;
wire n_5560;
wire n_5115;
wire n_5510;
wire n_5557;
wire n_5117;
wire n_5120;
wire n_5118;
wire n_5119;
wire n_5129;
wire n_5123;
wire n_5124;
wire n_5127;
wire n_5125;
wire n_5126;
wire n_5156;
wire n_5154;
wire n_5128;
wire n_5151;
wire n_5153;
wire n_5134;
wire n_5611;
wire n_5518;
wire n_5132;
wire n_5133;
wire n_5131;
wire n_5564;
wire n_5609;
wire n_5515;
wire n_5517;
wire n_5141;
wire n_5136;
wire n_5146;
wire n_5147;
wire n_5150;
wire n_5148;
wire n_5142;
wire n_5143;
wire n_5145;
wire n_5144;
wire n_5183;
wire n_5179;
wire n_5191;
wire n_5193;
wire n_5178;
wire n_5167;
wire n_5164;
wire n_5149;
wire n_5527;
wire n_5181;
wire n_5152;
wire n_5184;
wire n_5182;
wire n_5180;
wire n_5155;
wire n_5161;
wire n_5163;
wire n_5158;
wire n_5157;
wire n_5160;
wire n_5437;
wire n_5436;
wire n_5435;
wire n_5159;
wire n_5162;
wire n_5196;
wire n_5203;
wire n_5201;
wire n_5197;
wire n_5165;
wire n_5166;
wire n_5433;
wire n_5370;
wire n_5429;
wire n_5432;
wire n_5170;
wire n_5169;
wire n_5174;
wire n_5177;
wire n_5267;
wire n_5212;
wire n_5215;
wire n_5176;
wire n_5547;
wire n_5526;
wire n_5549;
wire n_5190;
wire n_5572;
wire n_5185;
wire n_5187;
wire n_5186;
wire n_5189;
wire n_5407;
wire n_5399;
wire n_5188;
wire n_5400;
wire n_5595;
wire n_5571;
wire n_5192;
wire n_5195;
wire n_5208;
wire n_5211;
wire n_5194;
wire n_5198;
wire n_5200;
wire n_5199;
wire n_5292;
wire n_5295;
wire n_5294;
wire n_5291;
wire n_5205;
wire n_5202;
wire n_5552;
wire n_5206;
wire n_5204;
wire n_5550;
wire n_5555;
wire n_5207;
wire n_5489;
wire n_5492;
wire n_5488;
wire n_5209;
wire n_5210;
wire n_5288;
wire n_5287;
wire n_5276;
wire n_5213;
wire n_5214;
wire n_5219;
wire n_5396;
wire n_5224;
wire n_5221;
wire n_5218;
wire n_5220;
wire n_5372;
wire n_5394;
wire n_5222;
wire n_5244;
wire n_5382;
wire n_5227;
wire n_5238;
wire n_5228;
wire n_5230;
wire n_5232;
wire n_5378;
wire n_5234;
wire n_5233;
wire n_5377;
wire n_5379;
wire n_5236;
wire n_5386;
wire n_5387;
wire n_5237;
wire n_5385;
wire n_5239;
wire n_5240;
wire n_5381;
wire n_5245;
wire n_5375;
wire n_5247;
wire n_5251;
wire n_5250;
wire n_5308;
wire n_5305;
wire n_5303;
wire n_5252;
wire n_5254;
wire n_5256;
wire n_5313;
wire n_5258;
wire n_5257;
wire n_5312;
wire n_5314;
wire n_5260;
wire n_5264;
wire n_5266;
wire n_5279;
wire n_5278;
wire n_5285;
wire n_5268;
wire n_5270;
wire n_5269;
wire n_5369;
wire n_5272;
wire n_5320;
wire n_5275;
wire n_5318;
wire n_5274;
wire n_5319;
wire n_5277;
wire n_5280;
wire n_5282;
wire n_5281;
wire n_5354;
wire n_5357;
wire n_5353;
wire n_5283;
wire n_5403;
wire n_5404;
wire n_5284;
wire n_5402;
wire n_5286;
wire n_5362;
wire n_5360;
wire n_5364;
wire n_5290;
wire n_5304;
wire n_5302;
wire n_5289;
wire n_5301;
wire n_5293;
wire n_5462;
wire n_5470;
wire n_5468;
wire n_5299;
wire n_5600;
wire n_5582;
wire n_5297;
wire n_5298;
wire n_5296;
wire n_5581;
wire n_5579;
wire n_5598;
wire n_5300;
wire n_5608;
wire n_5306;
wire n_5307;
wire n_5316;
wire n_5310;
wire n_5315;
wire n_5309;
wire n_5311;
wire n_5317;
wire n_5420;
wire n_5418;
wire n_5425;
wire n_5322;
wire n_5325;
wire n_5331;
wire n_5326;
wire n_5330;
wire n_5332;
wire n_5481;
wire n_5334;
wire n_5485;
wire n_5479;
wire n_5337;
wire n_5336;
wire n_5339;
wire n_5341;
wire n_5342;
wire n_5340;
wire n_5460;
wire n_5458;
wire n_5456;
wire n_5343;
wire n_5346;
wire n_5351;
wire n_5347;
wire n_5352;
wire n_5355;
wire n_5356;
wire n_5465;
wire n_5464;
wire n_5466;
wire n_5359;
wire n_5361;
wire n_5365;
wire n_5363;
wire n_5497;
wire n_5367;
wire n_5366;
wire n_5496;
wire n_5498;
wire n_5373;
wire n_5371;
wire n_5393;
wire n_5374;
wire n_5392;
wire n_5380;
wire n_5376;
wire n_5383;
wire n_5389;
wire n_5384;
wire n_5388;
wire n_5390;
wire n_5391;
wire n_5412;
wire n_5411;
wire n_5413;
wire n_5395;
wire n_5398;
wire n_5445;
wire n_5428;
wire n_5450;
wire n_5397;
wire n_5416;
wire n_5409;
wire n_5415;
wire n_5401;
wire n_5405;
wire n_5406;
wire n_5605;
wire n_5604;
wire n_5606;
wire n_5414;
wire n_5408;
wire n_5410;
wire n_5417;
wire n_5424;
wire n_5419;
wire n_5421;
wire n_5586;
wire n_5423;
wire n_5422;
wire n_5585;
wire n_5587;
wire n_5593;
wire n_5427;
wire n_5426;
wire n_5592;
wire n_5594;
wire n_5446;
wire n_5434;
wire n_5430;
wire n_5431;
wire n_5454;
wire n_5457;
wire n_5441;
wire n_5443;
wire n_5537;
wire n_5439;
wire n_5622;
wire n_5617;
wire n_5646;
wire n_5440;
wire n_5438;
wire n_5545;
wire n_5536;
wire n_5442;
wire n_5451;
wire n_5444;
wire n_5448;
wire n_5447;
wire n_5641;
wire n_5449;
wire n_5644;
wire n_5639;
wire n_5650;
wire n_5452;
wire n_5453;
wire n_5648;
wire n_5654;
wire n_5455;
wire n_5487;
wire n_5459;
wire n_5477;
wire n_5476;
wire n_5461;
wire n_5469;
wire n_5475;
wire n_5467;
wire n_5463;
wire n_5472;
wire n_5471;
wire n_5541;
wire n_5474;
wire n_5473;
wire n_5540;
wire n_5542;
wire n_5486;
wire n_5478;
wire n_5480;
wire n_5482;
wire n_5503;
wire n_5484;
wire n_5483;
wire n_5502;
wire n_5504;
wire n_5500;
wire n_5494;
wire n_5490;
wire n_5628;
wire n_5491;
wire n_5635;
wire n_5625;
wire n_5499;
wire n_5493;
wire n_5495;
wire n_5501;
wire n_5508;
wire n_5507;
wire n_5511;
wire n_5514;
wire n_5513;
wire n_5512;
wire n_5516;
wire n_7303;
wire n_7233;
wire n_7301;
wire n_5522;
wire n_5525;
wire n_7083;
wire n_5520;
wire n_5521;
wire n_5519;
wire n_7080;
wire n_7053;
wire n_5523;
wire n_5524;
wire n_5546;
wire n_5531;
wire n_5529;
wire n_7371;
wire n_5528;
wire n_5530;
wire n_7370;
wire n_7411;
wire n_5532;
wire n_5535;
wire n_5533;
wire n_5534;
wire n_5538;
wire n_5543;
wire n_5539;
wire n_7149;
wire n_7150;
wire n_5544;
wire n_7148;
wire n_7398;
wire n_7393;
wire n_7406;
wire n_5548;
wire n_7091;
wire n_5556;
wire n_5551;
wire n_7171;
wire n_7179;
wire n_7165;
wire n_5553;
wire n_7189;
wire n_5554;
wire n_7188;
wire n_7198;
wire n_7089;
wire n_7087;
wire n_5558;
wire n_5559;
wire n_7048;
wire n_7005;
wire n_7046;
wire n_5562;
wire n_5561;
wire n_7003;
wire n_7047;
wire n_7006;
wire n_7022;
wire n_5563;
wire n_5566;
wire n_5565;
wire n_5567;
wire n_5568;
wire n_5570;
wire n_5569;
wire n_5596;
wire n_5574;
wire n_7118;
wire n_5580;
wire n_5576;
wire n_5573;
wire n_5575;
wire n_7115;
wire n_7153;
wire n_5578;
wire n_5577;
wire n_5590;
wire n_5583;
wire n_5588;
wire n_5584;
wire n_5589;
wire n_7098;
wire n_7100;
wire n_7097;
wire n_5591;
wire n_5597;
wire n_5599;
wire n_5602;
wire n_5607;
wire n_7106;
wire n_5601;
wire n_5603;
wire n_7104;
wire n_7109;
wire n_5610;
wire n_5613;
wire n_7162;
wire n_5616;
wire n_5614;
wire n_5612;
wire n_7157;
wire n_7161;
wire n_5618;
wire n_5615;
wire n_5621;
wire n_5620;
wire n_5619;
wire n_5623;
wire n_5637;
wire n_5624;
wire n_5627;
wire n_5626;
wire n_5629;
wire n_5632;
wire n_7409;
wire n_5631;
wire n_5630;
wire n_7408;
wire n_7410;
wire n_7176;
wire n_5634;
wire n_5633;
wire n_7175;
wire n_7177;
wire n_5636;
wire n_5638;
wire n_5640;
wire n_5642;
wire n_7194;
wire n_7195;
wire n_5643;
wire n_7193;
wire n_5645;
wire n_5647;
wire n_5649;
wire n_5651;
wire n_7182;
wire n_5653;
wire n_5652;
wire n_7181;
wire n_7183;
wire n_6998;
wire n_7199;
wire n_5657;
wire n_5659;
wire n_5662;
wire n_5661;
wire n_5698;
wire n_5696;
wire n_5712;
wire n_5708;
wire n_5663;
wire n_5664;
wire n_5667;
wire n_5687;
wire n_5686;
wire n_5674;
wire n_5670;
wire n_5673;
wire n_5671;
wire n_5672;
wire n_7571;
wire n_7574;
wire n_7479;
wire n_5677;
wire n_5676;
wire n_5714;
wire n_5722;
wire n_5713;
wire n_5681;
wire n_5679;
wire n_5680;
wire n_5710;
wire n_5682;
wire n_5685;
wire n_5683;
wire n_5684;
wire n_8068;
wire n_8066;
wire n_7920;
wire n_7472;
wire n_7471;
wire n_7469;
wire n_6088;
wire n_5691;
wire n_6011;
wire n_5693;
wire n_5694;
wire n_5707;
wire n_5700;
wire n_5697;
wire n_6042;
wire n_5701;
wire n_5699;
wire n_6016;
wire n_6044;
wire n_5702;
wire n_5705;
wire n_5703;
wire n_5704;
wire n_7485;
wire n_7484;
wire n_5706;
wire n_7481;
wire n_7483;
wire n_5709;
wire n_5711;
wire n_6852;
wire n_6770;
wire n_6849;
wire n_5718;
wire n_5721;
wire n_6058;
wire n_5716;
wire n_5717;
wire n_5715;
wire n_6060;
wire n_6050;
wire n_5719;
wire n_7581;
wire n_5720;
wire n_7576;
wire n_7717;
wire n_7585;
wire n_7643;
wire n_7583;
wire n_7582;
wire n_5723;
wire n_5725;
wire n_6008;
wire n_5731;
wire n_5729;
wire n_6093;
wire n_6602;
wire n_6601;
wire n_6092;
wire n_5739;
wire n_5736;
wire n_5735;
wire n_5734;
wire n_5996;
wire n_6000;
wire n_6002;
wire n_6003;
wire n_5738;
wire n_6395;
wire n_6390;
wire n_6385;
wire n_5744;
wire n_5745;
wire n_5750;
wire n_5992;
wire n_5991;
wire n_5749;
wire n_5990;
wire n_5754;
wire n_6559;
wire n_6586;
wire n_6585;
wire n_5758;
wire n_5853;
wire n_5761;
wire n_5763;
wire n_5766;
wire n_5765;
wire n_6483;
wire n_6482;
wire n_6480;
wire n_6481;
wire n_5767;
wire n_6479;
wire n_5770;
wire n_5769;
wire n_5772;
wire n_5776;
wire n_5774;
wire n_5773;
wire n_6583;
wire n_6582;
wire n_6581;
wire n_5775;
wire n_5786;
wire n_5779;
wire n_5785;
wire n_5793;
wire n_5815;
wire n_5814;
wire n_5792;
wire n_5813;
wire n_5796;
wire n_5795;
wire n_6576;
wire n_6575;
wire n_6573;
wire n_5797;
wire n_6574;
wire n_5799;
wire n_5802;
wire n_5800;
wire n_5804;
wire n_5809;
wire n_5808;
wire n_6477;
wire n_6468;
wire n_6470;
wire n_5816;
wire n_5817;
wire n_5820;
wire n_5819;
wire n_5822;
wire n_5851;
wire n_5847;
wire n_5824;
wire n_5831;
wire n_5843;
wire n_5844;
wire n_5827;
wire n_6578;
wire n_6570;
wire n_6571;
wire n_5830;
wire n_5835;
wire n_5833;
wire n_5834;
wire n_6655;
wire n_6654;
wire n_6653;
wire n_5837;
wire n_5840;
wire n_5839;
wire n_5842;
wire n_6293;
wire n_6292;
wire n_6290;
wire n_6291;
wire n_5841;
wire n_6289;
wire n_6650;
wire n_6649;
wire n_6648;
wire n_5846;
wire n_5845;
wire n_6651;
wire n_5849;
wire n_6563;
wire n_5848;
wire n_6560;
wire n_5850;
wire n_6566;
wire n_6565;
wire n_6569;
wire n_5852;
wire n_6562;
wire n_5856;
wire n_5855;
wire n_6636;
wire n_6658;
wire n_6661;
wire n_5857;
wire n_5858;
wire n_5862;
wire n_5988;
wire n_5987;
wire n_5986;
wire n_5861;
wire n_5866;
wire n_5868;
wire n_5867;
wire n_6644;
wire n_6646;
wire n_6640;
wire n_6638;
wire n_6637;
wire n_6643;
wire n_5869;
wire n_5909;
wire n_5873;
wire n_5872;
wire n_5908;
wire n_5876;
wire n_5875;
wire n_6676;
wire n_6675;
wire n_6674;
wire n_5877;
wire n_5880;
wire n_5879;
wire n_5882;
wire n_5884;
wire n_5883;
wire n_6303;
wire n_6300;
wire n_6302;
wire n_5885;
wire n_6301;
wire n_5903;
wire n_5897;
wire n_5894;
wire n_5902;
wire n_5896;
wire n_5901;
wire n_5907;
wire n_5910;
wire n_5912;
wire n_5911;
wire n_6665;
wire n_6663;
wire n_6664;
wire n_5913;
wire n_5918;
wire n_5922;
wire n_5920;
wire n_5919;
wire n_6258;
wire n_6257;
wire n_6256;
wire n_5921;
wire n_5950;
wire n_5947;
wire n_5934;
wire n_5941;
wire n_5946;
wire n_5949;
wire n_5952;
wire n_5951;
wire n_6315;
wire n_6313;
wire n_6314;
wire n_5953;
wire n_5955;
wire n_5957;
wire n_5956;
wire n_5960;
wire n_5959;
wire n_5964;
wire n_5972;
wire n_5962;
wire n_6310;
wire n_6308;
wire n_6309;
wire n_6282;
wire n_6281;
wire n_5961;
wire n_6312;
wire n_5976;
wire n_5967;
wire n_5969;
wire n_5968;
wire n_6295;
wire n_6288;
wire n_6287;
wire n_5971;
wire n_5973;
wire n_5975;
wire n_5974;
wire n_6220;
wire n_6219;
wire n_6217;
wire n_5981;
wire n_5985;
wire n_6626;
wire n_6633;
wire n_6631;
wire n_5989;
wire n_6616;
wire n_6623;
wire n_6612;
wire n_5993;
wire n_5997;
wire n_5999;
wire n_5998;
wire n_6117;
wire n_6028;
wire n_6030;
wire n_6029;
wire n_6027;
wire n_6001;
wire n_6605;
wire n_6613;
wire n_6610;
wire n_6606;
wire n_6004;
wire n_6006;
wire n_6005;
wire n_6021;
wire n_6018;
wire n_6024;
wire n_6022;
wire n_6007;
wire n_6012;
wire n_6015;
wire n_6013;
wire n_6014;
wire n_6043;
wire n_6017;
wire n_6019;
wire n_6020;
wire n_6861;
wire n_6859;
wire n_6854;
wire n_6023;
wire n_6026;
wire n_6038;
wire n_6041;
wire n_6025;
wire n_6120;
wire n_6102;
wire n_6032;
wire n_6331;
wire n_6037;
wire n_6034;
wire n_6031;
wire n_6033;
wire n_6334;
wire n_6325;
wire n_6035;
wire n_6036;
wire n_6076;
wire n_6074;
wire n_6072;
wire n_6039;
wire n_6040;
wire n_6063;
wire n_6066;
wire n_6062;
wire n_6045;
wire n_6049;
wire n_6052;
wire n_6047;
wire n_6046;
wire n_7488;
wire n_7558;
wire n_7555;
wire n_6048;
wire n_7497;
wire n_7489;
wire n_6051;
wire n_6059;
wire n_6053;
wire n_6054;
wire n_6057;
wire n_6055;
wire n_6056;
wire n_8079;
wire n_8078;
wire n_8073;
wire n_6084;
wire n_6061;
wire n_6702;
wire n_6704;
wire n_6696;
wire n_6065;
wire n_6064;
wire n_6068;
wire n_6067;
wire n_6071;
wire n_8217;
wire n_8216;
wire n_8211;
wire n_6069;
wire n_6070;
wire n_6073;
wire n_6106;
wire n_6108;
wire n_6104;
wire n_6075;
wire n_6340;
wire n_6083;
wire n_6358;
wire n_6077;
wire n_6082;
wire n_6080;
wire n_6078;
wire n_6079;
wire n_8260;
wire n_8257;
wire n_8250;
wire n_6081;
wire n_6338;
wire n_6085;
wire n_6086;
wire n_6087;
wire n_8209;
wire n_8197;
wire n_8235;
wire n_8196;
wire n_8198;
wire n_8234;
wire n_6091;
wire n_6766;
wire n_6090;
wire n_6095;
wire n_6098;
wire n_6101;
wire n_6100;
wire n_6099;
wire n_6105;
wire n_6103;
wire n_6243;
wire n_6238;
wire n_6236;
wire n_6107;
wire n_6115;
wire n_6111;
wire n_6110;
wire n_6116;
wire n_6109;
wire n_6114;
wire n_8154;
wire n_8153;
wire n_8146;
wire n_6112;
wire n_6113;
wire n_8120;
wire n_8118;
wire n_8111;
wire n_6119;
wire n_6118;
wire n_6121;
wire n_6136;
wire n_6122;
wire n_6249;
wire n_6139;
wire n_6130;
wire n_6252;
wire n_6234;
wire n_6126;
wire n_6320;
wire n_6319;
wire n_6125;
wire n_6150;
wire n_6128;
wire n_6131;
wire n_6129;
wire n_6133;
wire n_6132;
wire n_6135;
wire n_6364;
wire n_6363;
wire n_6361;
wire n_6360;
wire n_6134;
wire n_6362;
wire n_6137;
wire n_6138;
wire n_6140;
wire n_6206;
wire n_6142;
wire n_6141;
wire n_6207;
wire n_6199;
wire n_6347;
wire n_6345;
wire n_6343;
wire n_6342;
wire n_6344;
wire n_6143;
wire n_6346;
wire n_6353;
wire n_6145;
wire n_6149;
wire n_6232;
wire n_6153;
wire n_6192;
wire n_6148;
wire n_6197;
wire n_6195;
wire n_6233;
wire n_6231;
wire n_6152;
wire n_6193;
wire n_6191;
wire n_6160;
wire n_6186;
wire n_6185;
wire n_6156;
wire n_6157;
wire n_6284;
wire n_6279;
wire n_6276;
wire n_6278;
wire n_6159;
wire n_6184;
wire n_6163;
wire n_6162;
wire n_6228;
wire n_6227;
wire n_6225;
wire n_6226;
wire n_6164;
wire n_6224;
wire n_6167;
wire n_6166;
wire n_6171;
wire n_6173;
wire n_6168;
wire n_6174;
wire n_6172;
wire n_6541;
wire n_6540;
wire n_6539;
wire n_6177;
wire n_6181;
wire n_6183;
wire n_6222;
wire n_6188;
wire n_6215;
wire n_6187;
wire n_6190;
wire n_6189;
wire n_6196;
wire n_6200;
wire n_6198;
wire n_6274;
wire n_6283;
wire n_6269;
wire n_6201;
wire n_6205;
wire n_6204;
wire n_6202;
wire n_6203;
wire n_7522;
wire n_7521;
wire n_7520;
wire n_6209;
wire n_6214;
wire n_6213;
wire n_6208;
wire n_6211;
wire n_6210;
wire n_7528;
wire n_7527;
wire n_7525;
wire n_6212;
wire n_6223;
wire n_6230;
wire n_6216;
wire n_6218;
wire n_6221;
wire n_6229;
wire n_6235;
wire n_6239;
wire n_6237;
wire n_6241;
wire n_6240;
wire n_6244;
wire n_8151;
wire n_8150;
wire n_8148;
wire n_8149;
wire n_6242;
wire n_8147;
wire n_6247;
wire n_6246;
wire n_6245;
wire n_8159;
wire n_8158;
wire n_8157;
wire n_6248;
wire n_6254;
wire n_6250;
wire n_6251;
wire n_6270;
wire n_6280;
wire n_6275;
wire n_6268;
wire n_6253;
wire n_6255;
wire n_6261;
wire n_6266;
wire n_6265;
wire n_6260;
wire n_6259;
wire n_6264;
wire n_6377;
wire n_6375;
wire n_6376;
wire n_6262;
wire n_6263;
wire n_6350;
wire n_6352;
wire n_6267;
wire n_6351;
wire n_6271;
wire n_6273;
wire n_6272;
wire n_6369;
wire n_6367;
wire n_6368;
wire n_6297;
wire n_6277;
wire n_6285;
wire n_6307;
wire n_6298;
wire n_6306;
wire n_6286;
wire n_6294;
wire n_6296;
wire n_6299;
wire n_6305;
wire n_6304;
wire n_6311;
wire n_6318;
wire n_6316;
wire n_6317;
wire n_6321;
wire n_6324;
wire n_6323;
wire n_6322;
wire n_6326;
wire n_6328;
wire n_6327;
wire n_6330;
wire n_7508;
wire n_6329;
wire n_7501;
wire n_7506;
wire n_7505;
wire n_6333;
wire n_6332;
wire n_6336;
wire n_6335;
wire n_6380;
wire n_6511;
wire n_6359;
wire n_6337;
wire n_6339;
wire n_6348;
wire n_6356;
wire n_6341;
wire n_6357;
wire n_6349;
wire n_6355;
wire n_6354;
wire n_6374;
wire n_6366;
wire n_6373;
wire n_6365;
wire n_6371;
wire n_6672;
wire n_6370;
wire n_6372;
wire n_6671;
wire n_6668;
wire n_6379;
wire n_6378;
wire n_6514;
wire n_6506;
wire n_6384;
wire n_6597;
wire n_6383;
wire n_6596;
wire n_6386;
wire n_6389;
wire n_6387;
wire n_6799;
wire n_6388;
wire n_6840;
wire n_6839;
wire n_6800;
wire n_6795;
wire n_6391;
wire n_6394;
wire n_6397;
wire n_6454;
wire n_6453;
wire n_6547;
wire n_6396;
wire n_6455;
wire n_6400;
wire n_6521;
wire n_6528;
wire n_6516;
wire n_6425;
wire n_6405;
wire n_6424;
wire n_6404;
wire n_6416;
wire n_6408;
wire n_6814;
wire n_6815;
wire n_6813;
wire n_6411;
wire n_6415;
wire n_6418;
wire n_6421;
wire n_6420;
wire n_6423;
wire n_6834;
wire n_6833;
wire n_6832;
wire n_6422;
wire n_6428;
wire n_6427;
wire n_6536;
wire n_6535;
wire n_6534;
wire n_6429;
wire n_6527;
wire n_6437;
wire n_6434;
wire n_6433;
wire n_6436;
wire n_6432;
wire n_6810;
wire n_6809;
wire n_6807;
wire n_6808;
wire n_6435;
wire n_6806;
wire n_6438;
wire n_6443;
wire n_6442;
wire n_6448;
wire n_6447;
wire n_6452;
wire n_6457;
wire n_6504;
wire n_6503;
wire n_6458;
wire n_6500;
wire n_6495;
wire n_6499;
wire n_6497;
wire n_6461;
wire n_6464;
wire n_6463;
wire n_6489;
wire n_6487;
wire n_6490;
wire n_6492;
wire n_6467;
wire n_6469;
wire n_6471;
wire n_6476;
wire n_6478;
wire n_6485;
wire n_6484;
wire n_6488;
wire n_6739;
wire n_6738;
wire n_6736;
wire n_6491;
wire n_6722;
wire n_6721;
wire n_6720;
wire n_6498;
wire n_6494;
wire n_6496;
wire n_6824;
wire n_6829;
wire n_6828;
wire n_6823;
wire n_6816;
wire n_6805;
wire n_6804;
wire n_6501;
wire n_6502;
wire n_6510;
wire n_6505;
wire n_6508;
wire n_6507;
wire n_7515;
wire n_7517;
wire n_7514;
wire n_6509;
wire n_6512;
wire n_6513;
wire n_6546;
wire n_6544;
wire n_6517;
wire n_6525;
wire n_6522;
wire n_6543;
wire n_6515;
wire n_6520;
wire n_6518;
wire n_6519;
wire n_7619;
wire n_7618;
wire n_7617;
wire n_6523;
wire n_6524;
wire n_6530;
wire n_7610;
wire n_7611;
wire n_7608;
wire n_6526;
wire n_6529;
wire n_6533;
wire n_6531;
wire n_7609;
wire n_6532;
wire n_7607;
wire n_6538;
wire n_6537;
wire n_6542;
wire n_6545;
wire n_7614;
wire n_7613;
wire n_7606;
wire n_6550;
wire n_6549;
wire n_6900;
wire n_6904;
wire n_6907;
wire n_6558;
wire n_6554;
wire n_6556;
wire n_6553;
wire n_6557;
wire n_6555;
wire n_6801;
wire n_6820;
wire n_6819;
wire n_6802;
wire n_6561;
wire n_6751;
wire n_6752;
wire n_6750;
wire n_6564;
wire n_6746;
wire n_6745;
wire n_6744;
wire n_6567;
wire n_6568;
wire n_6580;
wire n_6572;
wire n_6579;
wire n_6589;
wire n_6593;
wire n_6592;
wire n_6588;
wire n_6587;
wire n_6591;
wire n_6717;
wire n_6714;
wire n_6716;
wire n_6590;
wire n_6715;
wire n_6741;
wire n_6733;
wire n_6734;
wire n_6594;
wire n_6595;
wire n_6598;
wire n_6600;
wire n_6599;
wire n_6782;
wire n_6787;
wire n_6790;
wire n_6781;
wire n_6604;
wire n_6764;
wire n_6763;
wire n_6762;
wire n_6603;
wire n_6607;
wire n_6609;
wire n_6608;
wire n_6873;
wire n_6865;
wire n_6916;
wire n_6914;
wire n_6864;
wire n_6611;
wire n_6694;
wire n_6620;
wire n_6621;
wire n_6693;
wire n_6614;
wire n_6622;
wire n_6615;
wire n_6617;
wire n_6619;
wire n_6618;
wire n_6727;
wire n_6711;
wire n_6756;
wire n_6753;
wire n_6710;
wire n_6624;
wire n_6689;
wire n_6625;
wire n_6627;
wire n_6630;
wire n_6628;
wire n_6629;
wire n_6725;
wire n_6712;
wire n_6635;
wire n_6632;
wire n_6684;
wire n_6683;
wire n_6634;
wire n_6639;
wire n_6641;
wire n_6895;
wire n_6642;
wire n_6896;
wire n_6894;
wire n_6645;
wire n_6657;
wire n_6647;
wire n_6656;
wire n_6652;
wire n_6659;
wire n_6660;
wire n_6662;
wire n_6679;
wire n_6666;
wire n_6673;
wire n_6669;
wire n_6667;
wire n_6670;
wire n_6681;
wire n_6680;
wire n_6891;
wire n_6889;
wire n_6890;
wire n_6881;
wire n_6880;
wire n_6682;
wire n_6893;
wire n_6688;
wire n_6883;
wire n_6686;
wire n_6685;
wire n_6687;
wire n_6882;
wire n_6876;
wire n_6875;
wire n_6879;
wire n_6878;
wire n_6690;
wire n_6692;
wire n_6691;
wire n_6870;
wire n_6866;
wire n_6698;
wire n_6695;
wire n_6697;
wire n_6700;
wire n_6699;
wire n_6703;
wire n_8103;
wire n_8106;
wire n_8084;
wire n_6701;
wire n_8085;
wire n_6709;
wire n_6705;
wire n_6706;
wire n_6708;
wire n_6707;
wire n_8138;
wire n_8141;
wire n_8133;
wire n_6713;
wire n_6719;
wire n_6718;
wire n_6724;
wire n_6723;
wire n_6732;
wire n_6726;
wire n_6729;
wire n_6728;
wire n_6731;
wire n_8116;
wire n_8115;
wire n_8113;
wire n_8114;
wire n_6730;
wire n_8112;
wire n_6749;
wire n_6743;
wire n_6737;
wire n_6735;
wire n_6748;
wire n_6742;
wire n_6747;
wire n_6755;
wire n_6754;
wire n_6757;
wire n_6759;
wire n_6761;
wire n_6760;
wire n_6758;
wire n_7664;
wire n_7667;
wire n_7660;
wire n_8096;
wire n_8095;
wire n_8087;
wire n_8086;
wire n_8094;
wire n_8097;
wire n_6772;
wire n_6778;
wire n_6777;
wire n_6765;
wire n_6767;
wire n_6769;
wire n_6768;
wire n_6771;
wire n_6773;
wire n_6775;
wire n_7490;
wire n_7498;
wire n_6774;
wire n_7494;
wire n_6776;
wire n_6780;
wire n_6844;
wire n_6779;
wire n_6843;
wire n_6783;
wire n_6784;
wire n_7531;
wire n_7530;
wire n_7507;
wire n_7500;
wire n_6785;
wire n_6786;
wire n_6789;
wire n_6788;
wire n_6792;
wire n_6791;
wire n_6794;
wire n_7602;
wire n_7601;
wire n_7597;
wire n_6793;
wire n_7599;
wire n_7598;
wire n_6838;
wire n_6797;
wire n_6796;
wire n_7543;
wire n_7542;
wire n_7538;
wire n_6798;
wire n_7540;
wire n_7539;
wire n_6818;
wire n_6803;
wire n_6812;
wire n_6811;
wire n_6822;
wire n_6821;
wire n_6837;
wire n_6826;
wire n_6825;
wire n_7678;
wire n_7677;
wire n_7676;
wire n_6827;
wire n_6831;
wire n_6830;
wire n_6835;
wire n_7621;
wire n_7624;
wire n_7605;
wire n_6841;
wire n_6842;
wire n_6845;
wire n_6848;
wire n_6846;
wire n_6847;
wire n_7595;
wire n_7588;
wire n_7593;
wire n_7594;
wire n_6850;
wire n_6851;
wire n_6853;
wire n_6929;
wire n_6855;
wire n_6857;
wire n_6856;
wire n_7656;
wire n_7646;
wire n_7695;
wire n_7693;
wire n_6858;
wire n_6863;
wire n_6860;
wire n_6925;
wire n_6928;
wire n_6862;
wire n_6868;
wire n_6867;
wire n_7684;
wire n_7683;
wire n_7670;
wire n_6869;
wire n_7669;
wire n_6872;
wire n_6871;
wire n_6874;
wire n_6899;
wire n_8101;
wire n_8100;
wire n_8099;
wire n_6877;
wire n_6884;
wire n_6888;
wire n_6886;
wire n_6885;
wire n_8126;
wire n_8125;
wire n_8123;
wire n_6887;
wire n_8124;
wire n_6892;
wire n_6898;
wire n_6897;
wire n_6901;
wire n_6903;
wire n_6902;
wire n_7689;
wire n_7688;
wire n_7687;
wire n_6906;
wire n_6905;
wire n_6909;
wire n_6908;
wire n_6912;
wire n_6911;
wire n_8092;
wire n_8091;
wire n_8089;
wire n_6910;
wire n_8090;
wire n_7679;
wire n_7672;
wire n_7674;
wire n_6913;
wire n_7673;
wire n_6922;
wire n_6915;
wire n_6924;
wire n_6917;
wire n_6919;
wire n_6921;
wire n_6918;
wire n_7699;
wire n_7698;
wire n_6920;
wire n_6923;
wire n_7648;
wire n_7654;
wire n_7647;
wire n_6926;
wire n_6927;
wire n_8130;
wire n_8129;
wire n_8082;
wire n_6930;
wire n_6933;
wire n_6931;
wire n_6932;
wire n_7638;
wire n_7586;
wire n_6937;
wire n_7914;
wire n_7736;
wire n_7734;
wire n_6940;
wire n_6946;
wire n_6944;
wire n_6945;
wire n_6951;
wire n_6947;
wire n_6950;
wire n_6948;
wire n_6949;
wire n_6986;
wire n_6981;
wire n_6978;
wire n_6953;
wire n_6956;
wire n_7759;
wire n_6957;
wire n_6960;
wire n_6955;
wire n_7741;
wire n_7761;
wire n_6958;
wire n_6959;
wire n_7208;
wire n_7207;
wire n_7205;
wire n_6966;
wire n_6962;
wire n_6976;
wire n_6972;
wire n_6967;
wire n_6968;
wire n_6971;
wire n_6969;
wire n_6970;
wire n_7216;
wire n_7219;
wire n_7203;
wire n_6977;
wire n_6973;
wire n_6974;
wire n_6994;
wire n_6996;
wire n_6979;
wire n_8656;
wire n_8658;
wire n_6980;
wire n_8323;
wire n_8404;
wire n_6982;
wire n_6984;
wire n_6993;
wire n_6983;
wire n_6990;
wire n_6988;
wire n_6985;
wire n_7011;
wire n_7013;
wire n_7015;
wire n_6987;
wire n_6992;
wire n_6991;
wire n_6989;
wire n_7025;
wire n_7031;
wire n_7029;
wire n_7010;
wire n_6995;
wire n_7007;
wire n_7021;
wire n_7008;
wire n_6999;
wire n_7201;
wire n_7001;
wire n_7002;
wire n_7004;
wire n_7009;
wire n_8865;
wire n_7012;
wire n_8841;
wire n_8867;
wire n_7014;
wire n_7839;
wire n_7019;
wire n_7017;
wire n_7020;
wire n_7016;
wire n_7018;
wire n_7841;
wire n_7827;
wire n_7824;
wire n_7315;
wire n_7308;
wire n_7314;
wire n_7042;
wire n_7024;
wire n_7023;
wire n_7041;
wire n_7026;
wire n_7028;
wire n_7027;
wire n_7067;
wire n_7066;
wire n_7064;
wire n_7030;
wire n_7039;
wire n_7034;
wire n_7033;
wire n_7037;
wire n_7032;
wire n_7038;
wire n_7279;
wire n_7276;
wire n_7278;
wire n_7035;
wire n_7036;
wire n_7040;
wire n_7357;
wire n_7358;
wire n_7349;
wire n_7043;
wire n_7045;
wire n_7044;
wire n_7058;
wire n_7056;
wire n_7061;
wire n_7059;
wire n_7055;
wire n_7155;
wire n_7052;
wire n_7049;
wire n_7051;
wire n_7050;
wire n_7054;
wire n_7374;
wire n_7378;
wire n_7057;
wire n_7379;
wire n_7377;
wire n_7375;
wire n_7063;
wire n_7060;
wire n_7078;
wire n_7076;
wire n_7062;
wire n_7065;
wire n_7908;
wire n_7902;
wire n_7911;
wire n_7074;
wire n_7069;
wire n_7070;
wire n_7073;
wire n_7068;
wire n_7338;
wire n_7336;
wire n_7337;
wire n_7071;
wire n_7072;
wire n_7777;
wire n_7075;
wire n_7780;
wire n_7775;
wire n_7077;
wire n_7127;
wire n_7126;
wire n_7120;
wire n_7079;
wire n_7125;
wire n_7082;
wire n_7081;
wire n_7084;
wire n_7112;
wire n_7114;
wire n_7085;
wire n_7088;
wire n_7086;
wire n_7102;
wire n_7101;
wire n_7090;
wire n_7093;
wire n_7095;
wire n_7092;
wire n_7266;
wire n_7094;
wire n_7269;
wire n_7264;
wire n_7096;
wire n_7099;
wire n_7134;
wire n_7131;
wire n_7135;
wire n_7103;
wire n_7108;
wire n_7105;
wire n_7107;
wire n_7143;
wire n_7144;
wire n_7140;
wire n_7123;
wire n_7111;
wire n_7110;
wire n_7122;
wire n_7124;
wire n_7113;
wire n_7328;
wire n_7154;
wire n_7117;
wire n_7116;
wire n_7119;
wire n_7146;
wire n_7121;
wire n_7139;
wire n_7130;
wire n_7138;
wire n_7129;
wire n_7137;
wire n_7128;
wire n_7136;
wire n_7132;
wire n_7133;
wire n_7145;
wire n_7141;
wire n_7142;
wire n_7147;
wire n_7151;
wire n_7152;
wire n_7333;
wire n_7332;
wire n_7334;
wire n_7326;
wire n_7343;
wire n_7156;
wire n_7159;
wire n_7158;
wire n_7160;
wire n_7273;
wire n_7271;
wire n_7262;
wire n_7164;
wire n_7168;
wire n_7187;
wire n_7185;
wire n_7163;
wire n_7184;
wire n_7167;
wire n_7166;
wire n_7169;
wire n_7170;
wire n_7173;
wire n_7178;
wire n_7431;
wire n_7172;
wire n_7174;
wire n_7428;
wire n_7445;
wire n_7180;
wire n_7186;
wire n_7197;
wire n_7191;
wire n_7190;
wire n_7192;
wire n_7196;
wire n_7457;
wire n_7458;
wire n_7454;
wire n_7202;
wire n_7228;
wire n_7204;
wire n_7206;
wire n_7846;
wire n_7819;
wire n_7848;
wire n_7212;
wire n_7810;
wire n_7210;
wire n_7209;
wire n_7211;
wire n_7813;
wire n_7767;
wire n_7213;
wire n_7215;
wire n_7214;
wire n_7894;
wire n_7238;
wire n_7241;
wire n_7239;
wire n_7237;
wire n_7218;
wire n_7217;
wire n_7220;
wire n_7224;
wire n_7227;
wire n_7221;
wire n_7223;
wire n_7222;
wire n_7306;
wire n_7321;
wire n_7320;
wire n_7307;
wire n_7225;
wire n_7226;
wire n_7251;
wire n_7248;
wire n_7235;
wire n_7229;
wire n_7232;
wire n_7231;
wire n_7230;
wire n_7234;
wire n_7236;
wire n_7896;
wire n_7880;
wire n_7247;
wire n_7784;
wire n_7240;
wire n_7243;
wire n_7242;
wire n_7246;
wire n_7289;
wire n_7292;
wire n_7291;
wire n_7244;
wire n_7245;
wire n_7783;
wire n_7771;
wire n_7249;
wire n_7260;
wire n_7253;
wire n_7250;
wire n_7252;
wire n_7259;
wire n_7258;
wire n_7254;
wire n_7257;
wire n_7255;
wire n_7256;
wire n_7423;
wire n_7422;
wire n_7413;
wire n_7261;
wire n_7263;
wire n_7265;
wire n_7267;
wire n_7268;
wire n_7284;
wire n_7283;
wire n_7285;
wire n_7270;
wire n_7272;
wire n_7275;
wire n_7287;
wire n_7274;
wire n_7277;
wire n_7281;
wire n_7286;
wire n_7803;
wire n_7280;
wire n_7282;
wire n_7800;
wire n_7809;
wire n_7288;
wire n_7290;
wire n_7462;
wire n_7464;
wire n_7461;
wire n_7295;
wire n_7299;
wire n_7298;
wire n_7294;
wire n_7293;
wire n_7297;
wire n_7450;
wire n_7449;
wire n_7447;
wire n_7448;
wire n_7296;
wire n_7446;
wire n_7443;
wire n_7442;
wire n_7440;
wire n_7441;
wire n_7300;
wire n_7439;
wire n_7302;
wire n_7305;
wire n_7367;
wire n_7369;
wire n_7304;
wire n_7313;
wire n_7310;
wire n_7309;
wire n_7417;
wire n_7419;
wire n_7414;
wire n_7311;
wire n_7312;
wire n_7319;
wire n_7317;
wire n_8848;
wire n_7833;
wire n_7318;
wire n_7316;
wire n_8863;
wire n_8850;
wire n_7836;
wire n_7828;
wire n_7348;
wire n_7323;
wire n_7324;
wire n_7347;
wire n_7322;
wire n_7344;
wire n_7325;
wire n_7330;
wire n_7327;
wire n_7335;
wire n_7329;
wire n_7331;
wire n_7342;
wire n_8879;
wire n_7905;
wire n_7340;
wire n_8891;
wire n_8894;
wire n_8888;
wire n_7341;
wire n_7339;
wire n_7904;
wire n_7907;
wire n_8878;
wire n_8881;
wire n_7365;
wire n_7346;
wire n_7345;
wire n_7364;
wire n_7366;
wire n_7353;
wire n_7350;
wire n_7351;
wire n_7383;
wire n_7352;
wire n_7355;
wire n_7384;
wire n_7354;
wire n_7356;
wire n_7385;
wire n_7362;
wire n_8883;
wire n_7360;
wire n_7361;
wire n_7359;
wire n_8870;
wire n_8885;
wire n_7363;
wire n_8857;
wire n_8861;
wire n_8854;
wire n_7368;
wire n_7412;
wire n_7373;
wire n_7392;
wire n_7396;
wire n_7372;
wire n_7391;
wire n_7376;
wire n_7404;
wire n_7405;
wire n_7402;
wire n_7380;
wire n_7389;
wire n_7381;
wire n_7382;
wire n_7388;
wire n_7831;
wire n_7387;
wire n_7386;
wire n_7830;
wire n_7832;
wire n_7390;
wire n_7395;
wire n_7394;
wire n_7397;
wire n_7400;
wire n_7399;
wire n_7403;
wire n_7401;
wire n_7407;
wire n_7416;
wire n_7791;
wire n_7415;
wire n_7794;
wire n_7789;
wire n_7418;
wire n_7421;
wire n_7436;
wire n_7420;
wire n_7435;
wire n_7437;
wire n_7434;
wire n_7453;
wire n_7426;
wire n_7452;
wire n_7425;
wire n_7451;
wire n_7424;
wire n_7427;
wire n_7444;
wire n_7430;
wire n_7429;
wire n_7432;
wire n_7438;
wire n_7433;
wire n_7459;
wire n_7455;
wire n_7456;
wire n_7460;
wire n_7463;
wire n_7732;
wire n_7466;
wire n_7468;
wire n_7919;
wire n_8185;
wire n_8182;
wire n_7473;
wire n_7474;
wire n_7726;
wire n_7478;
wire n_7477;
wire n_7725;
wire n_7480;
wire n_7482;
wire n_8072;
wire n_8168;
wire n_8170;
wire n_8071;
wire n_7487;
wire n_7567;
wire n_7486;
wire n_7566;
wire n_7491;
wire n_7493;
wire n_7492;
wire n_8265;
wire n_8268;
wire n_8249;
wire n_7499;
wire n_7495;
wire n_7496;
wire n_7552;
wire n_7554;
wire n_7504;
wire n_7502;
wire n_7503;
wire n_8290;
wire n_8289;
wire n_8287;
wire n_7509;
wire n_7513;
wire n_7511;
wire n_7510;
wire n_8255;
wire n_8254;
wire n_8252;
wire n_7512;
wire n_7516;
wire n_7519;
wire n_7523;
wire n_7518;
wire n_7524;
wire n_7526;
wire n_7529;
wire n_7533;
wire n_7537;
wire n_7535;
wire n_7532;
wire n_7536;
wire n_7534;
wire n_8225;
wire n_8230;
wire n_8233;
wire n_8226;
wire n_7994;
wire n_7993;
wire n_7991;
wire n_7541;
wire n_7992;
wire n_7546;
wire n_7550;
wire n_7549;
wire n_7545;
wire n_7544;
wire n_7548;
wire n_8004;
wire n_8003;
wire n_8001;
wire n_8002;
wire n_7547;
wire n_8000;
wire n_8011;
wire n_8010;
wire n_8008;
wire n_8009;
wire n_7551;
wire n_8007;
wire n_7553;
wire n_8281;
wire n_8295;
wire n_8294;
wire n_8282;
wire n_7557;
wire n_7556;
wire n_7559;
wire n_7561;
wire n_7563;
wire n_7562;
wire n_7560;
wire n_8014;
wire n_7987;
wire n_8025;
wire n_8024;
wire n_7986;
wire n_8273;
wire n_8247;
wire n_8272;
wire n_7564;
wire n_7565;
wire n_7568;
wire n_7570;
wire n_8208;
wire n_8201;
wire n_7569;
wire n_8245;
wire n_8243;
wire n_8195;
wire n_7573;
wire n_7572;
wire n_7575;
wire n_7722;
wire n_7721;
wire n_7577;
wire n_7580;
wire n_7578;
wire n_7579;
wire n_7983;
wire n_7981;
wire n_7960;
wire n_7584;
wire n_7716;
wire n_7587;
wire n_7589;
wire n_7591;
wire n_7590;
wire n_7998;
wire n_7988;
wire n_8013;
wire n_7592;
wire n_7596;
wire n_7633;
wire n_7995;
wire n_7989;
wire n_7600;
wire n_7604;
wire n_7630;
wire n_7629;
wire n_7603;
wire n_7628;
wire n_7612;
wire n_7616;
wire n_7615;
wire n_7620;
wire n_7622;
wire n_7623;
wire n_7625;
wire n_7627;
wire n_7626;
wire n_8038;
wire n_8036;
wire n_8037;
wire n_8291;
wire n_8285;
wire n_8284;
wire n_7631;
wire n_7632;
wire n_7635;
wire n_7634;
wire n_8042;
wire n_8046;
wire n_8033;
wire n_8028;
wire n_7636;
wire n_7637;
wire n_7639;
wire n_7645;
wire n_7640;
wire n_7714;
wire n_7641;
wire n_7642;
wire n_8438;
wire n_8437;
wire n_8411;
wire n_7644;
wire n_7712;
wire n_7650;
wire n_7649;
wire n_8030;
wire n_8029;
wire n_7651;
wire n_7652;
wire n_7653;
wire n_7655;
wire n_7658;
wire n_7668;
wire n_7657;
wire n_7659;
wire n_7662;
wire n_7661;
wire n_8449;
wire n_8448;
wire n_8446;
wire n_8447;
wire n_7663;
wire n_8445;
wire n_7665;
wire n_7666;
wire n_7682;
wire n_7671;
wire n_7675;
wire n_7681;
wire n_7680;
wire n_7686;
wire n_7685;
wire n_7692;
wire n_7690;
wire n_7694;
wire n_7697;
wire n_7710;
wire n_7709;
wire n_7696;
wire n_7707;
wire n_7702;
wire n_7706;
wire n_7701;
wire n_7705;
wire n_7700;
wire n_8563;
wire n_8561;
wire n_8562;
wire n_7703;
wire n_7704;
wire n_8452;
wire n_8451;
wire n_8444;
wire n_7708;
wire n_8443;
wire n_8441;
wire n_8458;
wire n_8455;
wire n_7711;
wire n_8442;
wire n_7713;
wire n_7715;
wire n_7718;
wire n_7720;
wire n_7719;
wire n_8410;
wire n_8470;
wire n_8469;
wire n_8409;
wire n_8188;
wire n_8192;
wire n_8202;
wire n_7723;
wire n_7724;
wire n_7728;
wire n_7727;
wire n_7751;
wire n_7743;
wire n_7749;
wire n_7729;
wire n_7730;
wire n_7731;
wire n_7750;
wire n_7922;
wire n_7753;
wire n_7735;
wire n_7739;
wire n_7738;
wire n_8317;
wire n_7918;
wire n_7917;
wire n_7758;
wire n_7740;
wire n_7742;
wire n_7744;
wire n_7746;
wire n_7745;
wire n_8660;
wire n_8662;
wire n_8665;
wire n_7747;
wire n_8661;
wire n_7748;
wire n_8911;
wire n_7754;
wire n_7757;
wire n_7752;
wire n_7958;
wire n_7926;
wire n_7755;
wire n_7756;
wire n_7864;
wire n_7863;
wire n_7850;
wire n_7760;
wire n_7763;
wire n_7818;
wire n_7766;
wire n_7816;
wire n_7762;
wire n_7817;
wire n_7765;
wire n_7764;
wire n_7768;
wire n_7770;
wire n_7769;
wire n_7773;
wire n_7772;
wire n_7781;
wire n_7774;
wire n_7776;
wire n_7778;
wire n_7889;
wire n_7779;
wire n_7891;
wire n_7888;
wire n_8335;
wire n_8336;
wire n_7782;
wire n_8334;
wire n_7798;
wire n_7797;
wire n_7787;
wire n_7786;
wire n_7796;
wire n_7785;
wire n_7795;
wire n_7788;
wire n_7790;
wire n_7792;
wire n_7793;
wire n_8396;
wire n_8395;
wire n_8397;
wire n_7799;
wire n_7808;
wire n_7802;
wire n_7801;
wire n_7804;
wire n_7805;
wire n_8346;
wire n_8348;
wire n_8343;
wire n_8387;
wire n_7807;
wire n_7806;
wire n_8386;
wire n_8388;
wire n_7812;
wire n_7811;
wire n_7814;
wire n_8772;
wire n_7815;
wire n_8326;
wire n_8769;
wire n_8738;
wire n_8328;
wire n_8353;
wire n_7820;
wire n_7823;
wire n_7822;
wire n_7821;
wire n_7826;
wire n_7825;
wire n_7829;
wire n_7835;
wire n_7834;
wire n_7837;
wire n_8961;
wire n_7838;
wire n_8939;
wire n_8965;
wire n_8962;
wire n_8936;
wire n_8933;
wire n_7840;
wire n_8338;
wire n_7844;
wire n_7842;
wire n_7857;
wire n_7843;
wire n_7860;
wire n_7855;
wire n_8332;
wire n_7845;
wire n_8339;
wire n_8367;
wire n_8372;
wire n_8365;
wire n_7847;
wire n_7879;
wire n_7876;
wire n_7849;
wire n_7875;
wire n_7851;
wire n_7854;
wire n_7853;
wire n_7852;
wire n_7856;
wire n_8899;
wire n_8900;
wire n_8898;
wire n_7858;
wire n_7859;
wire n_7861;
wire n_8696;
wire n_7862;
wire n_7949;
wire n_8692;
wire n_8698;
wire n_7947;
wire n_7953;
wire n_7866;
wire n_7931;
wire n_7874;
wire n_7873;
wire n_7865;
wire n_7871;
wire n_7867;
wire n_7869;
wire n_7883;
wire n_7868;
wire n_7881;
wire n_7870;
wire n_7886;
wire n_7885;
wire n_7893;
wire n_7937;
wire n_7872;
wire n_7882;
wire n_7930;
wire n_7954;
wire n_7878;
wire n_7877;
wire n_7884;
wire n_7892;
wire n_7887;
wire n_7890;
wire n_7936;
wire n_7942;
wire n_7895;
wire n_7900;
wire n_7899;
wire n_7897;
wire n_8391;
wire n_7898;
wire n_8389;
wire n_8385;
wire n_8383;
wire n_7909;
wire n_7901;
wire n_7910;
wire n_7903;
wire n_7906;
wire n_7915;
wire n_7916;
wire n_8065;
wire n_7924;
wire n_7921;
wire n_7923;
wire n_8064;
wire n_8061;
wire n_7959;
wire n_7925;
wire n_7957;
wire n_7956;
wire n_7928;
wire n_7927;
wire n_7929;
wire n_7945;
wire n_7934;
wire n_7944;
wire n_7933;
wire n_7943;
wire n_7932;
wire n_7935;
wire n_7941;
wire n_7939;
wire n_7976;
wire n_7938;
wire n_7940;
wire n_7975;
wire n_7972;
wire n_7946;
wire n_7952;
wire n_7948;
wire n_8722;
wire n_8721;
wire n_8725;
wire n_7950;
wire n_7951;
wire n_8724;
wire n_7965;
wire n_7979;
wire n_7955;
wire n_7964;
wire n_8060;
wire n_7962;
wire n_7961;
wire n_7963;
wire n_7978;
wire n_7968;
wire n_7973;
wire n_7971;
wire n_7967;
wire n_7966;
wire n_7970;
wire n_8377;
wire n_8376;
wire n_8374;
wire n_8375;
wire n_7969;
wire n_8373;
wire n_7974;
wire n_7977;
wire n_7980;
wire n_8416;
wire n_8415;
wire n_8431;
wire n_7982;
wire n_7985;
wire n_8058;
wire n_8055;
wire n_7984;
wire n_7990;
wire n_7996;
wire n_7997;
wire n_7999;
wire n_8006;
wire n_8005;
wire n_8012;
wire n_8022;
wire n_8017;
wire n_8021;
wire n_8016;
wire n_8020;
wire n_8015;
wire n_8428;
wire n_8427;
wire n_8426;
wire n_8018;
wire n_8019;
wire n_8436;
wire n_8435;
wire n_8433;
wire n_8023;
wire n_8434;
wire n_8027;
wire n_8052;
wire n_8051;
wire n_8026;
wire n_8050;
wire n_8031;
wire n_8032;
wire n_8034;
wire n_8041;
wire n_8035;
wire n_8039;
wire n_8040;
wire n_8043;
wire n_8048;
wire n_8044;
wire n_8045;
wire n_8421;
wire n_8419;
wire n_8420;
wire n_8047;
wire n_8049;
wire n_8706;
wire n_8704;
wire n_8703;
wire n_8053;
wire n_8054;
wire n_8057;
wire n_8674;
wire n_8056;
wire n_8669;
wire n_8673;
wire n_8059;
wire n_8062;
wire n_8063;
wire n_8358;
wire n_8357;
wire n_8356;
wire n_8067;
wire n_8070;
wire n_8178;
wire n_8181;
wire n_8069;
wire n_8074;
wire n_8077;
wire n_8075;
wire n_8076;
wire n_8568;
wire n_8566;
wire n_8553;
wire n_8164;
wire n_8081;
wire n_8080;
wire n_8163;
wire n_8083;
wire n_8088;
wire n_8093;
wire n_8098;
wire n_8102;
wire n_8105;
wire n_8104;
wire n_8109;
wire n_8107;
wire n_8110;
wire n_8108;
wire n_8541;
wire n_8540;
wire n_8538;
wire n_8117;
wire n_8119;
wire n_8121;
wire n_8128;
wire n_8122;
wire n_8127;
wire n_8132;
wire n_8162;
wire n_8161;
wire n_8131;
wire n_8160;
wire n_8135;
wire n_8134;
wire n_8548;
wire n_8547;
wire n_8546;
wire n_8136;
wire n_8137;
wire n_8140;
wire n_8139;
wire n_8142;
wire n_8144;
wire n_8145;
wire n_8143;
wire n_8605;
wire n_8604;
wire n_8602;
wire n_8152;
wire n_8156;
wire n_8155;
wire n_8558;
wire n_8557;
wire n_8555;
wire n_8554;
wire n_8556;
wire n_8559;
wire n_8165;
wire n_8166;
wire n_8527;
wire n_8530;
wire n_8518;
wire n_8519;
wire n_8167;
wire n_8529;
wire n_8531;
wire n_8543;
wire n_8535;
wire n_8169;
wire n_8177;
wire n_8174;
wire n_8172;
wire n_8175;
wire n_8171;
wire n_8176;
wire n_8173;
wire n_8595;
wire n_8625;
wire n_8628;
wire n_8594;
wire n_8517;
wire n_8550;
wire n_8549;
wire n_8406;
wire n_8180;
wire n_8179;
wire n_8512;
wire n_8513;
wire n_8516;
wire n_8514;
wire n_8407;
wire n_8183;
wire n_8184;
wire n_8314;
wire n_8186;
wire n_8312;
wire n_8313;
wire n_8187;
wire n_8189;
wire n_8191;
wire n_8190;
wire n_8584;
wire n_8587;
wire n_8586;
wire n_8583;
wire n_8194;
wire n_8193;
wire n_8203;
wire n_8199;
wire n_8200;
wire n_8236;
wire n_8238;
wire n_8239;
wire n_8242;
wire n_8246;
wire n_8310;
wire n_8307;
wire n_8207;
wire n_8204;
wire n_8206;
wire n_8205;
wire n_8687;
wire n_8686;
wire n_8668;
wire n_8210;
wire n_8212;
wire n_8213;
wire n_8542;
wire n_8536;
wire n_8214;
wire n_8215;
wire n_8544;
wire n_8224;
wire n_8219;
wire n_8220;
wire n_8223;
wire n_8218;
wire n_8608;
wire n_8607;
wire n_8600;
wire n_8221;
wire n_8222;
wire n_8609;
wire n_8227;
wire n_8229;
wire n_8228;
wire n_8613;
wire n_8612;
wire n_8611;
wire n_8231;
wire n_8237;
wire n_8597;
wire n_8616;
wire n_8615;
wire n_8598;
wire n_8240;
wire n_8241;
wire n_8648;
wire n_8646;
wire n_8631;
wire n_8244;
wire n_8306;
wire n_8305;
wire n_8248;
wire n_8256;
wire n_8253;
wire n_8251;
wire n_8258;
wire n_8259;
wire n_8261;
wire n_8263;
wire n_8262;
wire n_8639;
wire n_8640;
wire n_8637;
wire n_8264;
wire n_8638;
wire n_8266;
wire n_8267;
wire n_8269;
wire n_8271;
wire n_8270;
wire n_8643;
wire n_8635;
wire n_8633;
wire n_8280;
wire n_8276;
wire n_8275;
wire n_8279;
wire n_8274;
wire n_8678;
wire n_8677;
wire n_8676;
wire n_8277;
wire n_8278;
wire n_8283;
wire n_8288;
wire n_8286;
wire n_8292;
wire n_8302;
wire n_8298;
wire n_8301;
wire n_8297;
wire n_8300;
wire n_8296;
wire n_8712;
wire n_8711;
wire n_8709;
wire n_8299;
wire n_8710;
wire n_8683;
wire n_8682;
wire n_8681;
wire n_8303;
wire n_8304;
wire n_8308;
wire n_8309;
wire n_8716;
wire n_8715;
wire n_8311;
wire n_8702;
wire n_8316;
wire n_8315;
wire n_8324;
wire n_8327;
wire n_8402;
wire n_8403;
wire n_8319;
wire n_8318;
wire n_8321;
wire n_8655;
wire n_8320;
wire n_8322;
wire n_8325;
wire n_8354;
wire n_8352;
wire n_8329;
wire n_8331;
wire n_8330;
wire n_8340;
wire n_8333;
wire n_8337;
wire n_8351;
wire n_8368;
wire n_8342;
wire n_8341;
wire n_8350;
wire n_8349;
wire n_8344;
wire n_8345;
wire n_8355;
wire n_8378;
wire n_8500;
wire n_8489;
wire n_8499;
wire n_8363;
wire n_8477;
wire n_8362;
wire n_8360;
wire n_8361;
wire n_8359;
wire n_8475;
wire n_8483;
wire n_8371;
wire n_8364;
wire n_8366;
wire n_8369;
wire n_8496;
wire n_8370;
wire n_8495;
wire n_8497;
wire n_8380;
wire n_8379;
wire n_8382;
wire n_8381;
wire n_8384;
wire n_8399;
wire n_8390;
wire n_8393;
wire n_8394;
wire n_8398;
wire n_8392;
wire n_8750;
wire n_8400;
wire n_8401;
wire n_8742;
wire n_8749;
wire n_8405;
wire n_8582;
wire n_8408;
wire n_8413;
wire n_8412;
wire n_8414;
wire n_8430;
wire n_8425;
wire n_8418;
wire n_8424;
wire n_8417;
wire n_8422;
wire n_8432;
wire n_8440;
wire n_8466;
wire n_8465;
wire n_8439;
wire n_8464;
wire n_8450;
wire n_8453;
wire n_8454;
wire n_8457;
wire n_8456;
wire n_8459;
wire n_8460;
wire n_8461;
wire n_8509;
wire n_8508;
wire n_8507;
wire n_8463;
wire n_8462;
wire n_8510;
wire n_8504;
wire n_8502;
wire n_8503;
wire n_8467;
wire n_8468;
wire n_8488;
wire n_8486;
wire n_8473;
wire n_8472;
wire n_8485;
wire n_8471;
wire n_8484;
wire n_8474;
wire n_8476;
wire n_8480;
wire n_8479;
wire n_8482;
wire n_8524;
wire n_8478;
wire n_8747;
wire n_8746;
wire n_8744;
wire n_8745;
wire n_8481;
wire n_8743;
wire n_8523;
wire n_8526;
wire n_8487;
wire n_8492;
wire n_8490;
wire n_8498;
wire n_8491;
wire n_8493;
wire n_8494;
wire n_8501;
wire n_8506;
wire n_8505;
wire n_8580;
wire n_8579;
wire n_8515;
wire n_8522;
wire n_8520;
wire n_8521;
wire n_8528;
wire n_8533;
wire n_8532;
wire n_8827;
wire n_8826;
wire n_8824;
wire n_8534;
wire n_8825;
wire n_8539;
wire n_8537;
wire n_8545;
wire n_8575;
wire n_8552;
wire n_8551;
wire n_8574;
wire n_8560;
wire n_8564;
wire n_8565;
wire n_8567;
wire n_8570;
wire n_8569;
wire n_8766;
wire n_8765;
wire n_8764;
wire n_8571;
wire n_8572;
wire n_8577;
wire n_8576;
wire n_8761;
wire n_8759;
wire n_8760;
wire n_8578;
wire n_8806;
wire n_8830;
wire n_8805;
wire n_8581;
wire n_8813;
wire n_8771;
wire n_8585;
wire n_8775;
wire n_8777;
wire n_8780;
wire n_8590;
wire n_8593;
wire n_8589;
wire n_8588;
wire n_8592;
wire n_8753;
wire n_8740;
wire n_8757;
wire n_8591;
wire n_8741;
wire n_8596;
wire n_8599;
wire n_8601;
wire n_8603;
wire n_8606;
wire n_8610;
wire n_8614;
wire n_8623;
wire n_8619;
wire n_8622;
wire n_8618;
wire n_8621;
wire n_8617;
wire n_8792;
wire n_8791;
wire n_8789;
wire n_8790;
wire n_8620;
wire n_8788;
wire n_8819;
wire n_8818;
wire n_8816;
wire n_8817;
wire n_8624;
wire n_8815;
wire n_8626;
wire n_8627;
wire n_8654;
wire n_8629;
wire n_8652;
wire n_8653;
wire n_8630;
wire n_8634;
wire n_8632;
wire n_8636;
wire n_8641;
wire n_8642;
wire n_8647;
wire n_8650;
wire n_8649;
wire n_8802;
wire n_8801;
wire n_8799;
wire n_8651;
wire n_8800;
wire n_8808;
wire n_8812;
wire n_8657;
wire n_8843;
wire n_8840;
wire n_8659;
wire n_8839;
wire n_8930;
wire n_8929;
wire n_8664;
wire n_8663;
wire n_8666;
wire n_8735;
wire n_8737;
wire n_8667;
wire n_8670;
wire n_8672;
wire n_8671;
wire n_8785;
wire n_8796;
wire n_8787;
wire n_8675;
wire n_8680;
wire n_8679;
wire n_8685;
wire n_8684;
wire n_8689;
wire n_8701;
wire n_8691;
wire n_8688;
wire n_8700;
wire n_8690;
wire n_8693;
wire n_8694;
wire n_8695;
wire n_8905;
wire n_8903;
wire n_8904;
wire n_8697;
wire n_8699;
wire n_8731;
wire n_8730;
wire n_8734;
wire n_8705;
wire n_8707;
wire n_8714;
wire n_8708;
wire n_8713;
wire n_8728;
wire n_8719;
wire n_8727;
wire n_8718;
wire n_8726;
wire n_8717;
wire n_8720;
wire n_8723;
wire n_8729;
wire n_8733;
wire n_8732;
wire n_8736;
wire n_8739;
wire n_8756;
wire n_8748;
wire n_8754;
wire n_8755;
wire n_8758;
wire n_8763;
wire n_8762;
wire n_8768;
wire n_8770;
wire n_8774;
wire n_8773;
wire n_8803;
wire n_8776;
wire n_8943;
wire n_8945;
wire n_8942;
wire n_8779;
wire n_8778;
wire n_8783;
wire n_8781;
wire n_8784;
wire n_8782;
wire n_8954;
wire n_8953;
wire n_8951;
wire n_8786;
wire n_8797;
wire n_8793;
wire n_8798;
wire n_8804;
wire n_8833;
wire n_8837;
wire n_8836;
wire n_8832;
wire n_8807;
wire n_8811;
wire n_8810;
wire n_8809;
wire n_8814;
wire n_8822;
wire n_8820;
wire n_8823;
wire n_8828;
wire n_8831;
wire n_8835;
wire n_8925;
wire n_8924;
wire n_8922;
wire n_8923;
wire n_8834;
wire n_8921;
wire n_8970;
wire n_8969;
wire n_8968;
wire n_8838;
wire n_8842;
wire n_8844;
wire n_8845;
wire n_8847;
wire n_8846;
wire n_8919;
wire n_8864;
wire n_8853;
wire n_8852;
wire n_8851;
wire n_8862;
wire n_8855;
wire n_8856;
wire n_8916;
wire n_8913;
wire n_8866;
wire n_8871;
wire n_8869;
wire n_8910;
wire n_8868;
wire n_8872;
wire n_8882;
wire n_8875;
wire n_8873;
wire n_8874;
wire n_8876;
wire n_8877;
wire n_8884;
wire n_8897;
wire n_8887;
wire n_8886;
wire n_8896;
wire n_8895;
wire n_8889;
wire n_8890;
wire n_8902;
wire n_8901;
wire n_8914;
wire n_8912;
wire n_8915;
wire n_8917;
wire n_8918;
wire n_8920;
wire n_8928;
wire n_8934;
wire n_8963;
wire n_8960;
wire n_8932;
wire n_8931;
wire n_8959;
wire n_8935;
wire n_8938;
wire n_8937;
wire n_8940;
wire n_8949;
wire n_8941;
wire n_8944;
wire n_8952;
wire n_8950;
wire n_8966;
wire n_8964;
wire n_8967;
wire n_8977;
wire n_9022;
wire n_8978;
wire n_9007;
wire n_8980;
wire n_8982;
wire n_8987;
wire n_8985;
wire n_8988;
wire n_8991;
wire n_8997;
wire n_8998;
wire n_9001;
wire n_9010;
wire n_9014;
wire n_9011;
wire n_9033;
wire n_9012;
wire n_9013;
wire n_9032;
wire n_9034;
wire n_9015;
wire n_9018;
wire n_9023;
wire n_9024;
wire n_9031;
wire n_9035;
wire n_9030;
wire n_9028;
wire n_9029;
wire n_9036;
wire sgo__sro_n128;
wire sgo__sro_n129;
wire sgo__sro_n130;
wire sgo__sro_n81;
wire sgo__sro_n82;
wire sgo__sro_n83;
wire sgo__sro_n156;
wire sgo__sro_n157;
wire sgo__sro_n158;
wire CLOCK_opt_ipo_n324;
wire CLOCK_opt_ipo_n326;
wire CLOCK_opt_ipo_n333;
wire CLOCK_opt_ipo_n337;
wire CLOCK_opt_ipo_n345;
wire CLOCK_opt_ipo_n351;
wire CLOCK_opt_ipo_n418;
wire CLOCK_opt_ipo_n423;
wire CLOCK_opt_ipo_n425;
wire CLOCK_opt_ipo_n433;
wire CLOCK_opt_ipo_n528;


INV_X2 i_9102 (.ZN (n_9038), .A (B_imm[31]));
INV_X4 i_9101 (.ZN (n_9037), .A (A_imm[31]));
AOI22_X1 i_9100 (.ZN (n_9036), .A1 (A_imm[30]), .A2 (B_imm[31]), .B1 (B_imm[30]), .B2 (opt_ipoPP_0));
INV_X1 i_9099 (.ZN (n_9035), .A (n_9036));
AOI22_X1 i_9098 (.ZN (n_9034), .A1 (A_imm[29]), .A2 (B_imm[31]), .B1 (B_imm[29]), .B2 (opt_ipoPP_0));
NAND2_X1 i_9097 (.ZN (n_9033), .A1 (A_imm[30]), .A2 (B_imm[30]));
NAND4_X1 i_9096 (.ZN (n_9032), .A1 (A_imm[29]), .A2 (B_imm[31]), .A3 (B_imm[29]), .A4 (opt_ipoPP_0));
AOI21_X1 i_9095 (.ZN (n_9031), .A (n_9034), .B1 (n_9033), .B2 (n_9032));
NAND4_X1 i_9094 (.ZN (n_9030), .A1 (A_imm[30]), .A2 (B_imm[31]), .A3 (B_imm[30]), .A4 (opt_ipoPP_0));
INV_X1 i_9093 (.ZN (n_9029), .A (n_9030));
OAI21_X1 i_9092 (.ZN (n_9028), .A (n_9035), .B1 (n_9031), .B2 (n_9029));
OR3_X1 i_9091 (.ZN (n_9027), .A1 (n_9028), .A2 (n_9038), .A3 (n_9037));
OAI21_X1 i_9090 (.ZN (n_9026), .A (n_9028), .B1 (n_9038), .B2 (n_9037));
INV_X1 i_9089 (.ZN (n_9025), .A (n_9026));
NAND2_X1 i_9088 (.ZN (n_9024), .A1 (n_9035), .A2 (n_9030));
XNOR2_X1 i_9087 (.ZN (n_9023), .A (n_9024), .B (n_9031));
INV_X1 i_9086 (.ZN (n_9022), .A (n_9023));
INV_X2 i_9085 (.ZN (n_9021), .A (B_imm[28]));
INV_X2 i_9084 (.ZN (n_9020), .A (A_imm[28]));
OAI22_X1 i_9083 (.ZN (n_9019), .A1 (n_9038), .A2 (n_9020), .B1 (n_9021), .B2 (n_9037));
NAND2_X1 i_9082 (.ZN (n_9018), .A1 (A_imm[29]), .A2 (B_imm[30]));
INV_X1 i_9081 (.ZN (n_9017), .A (n_9018));
NAND4_X1 i_9080 (.ZN (n_9016), .A1 (B_imm[31]), .A2 (B_imm[28]), .A3 (opt_ipoPP_0), .A4 (A_imm[28]));
INV_X1 i_9079 (.ZN (n_9015), .A (n_9016));
OAI21_X1 i_9078 (.ZN (n_9014), .A (n_9019), .B1 (n_9017), .B2 (n_9015));
INV_X1 i_9077 (.ZN (n_9013), .A (n_9034));
NAND2_X1 i_9076 (.ZN (n_9012), .A1 (n_9013), .A2 (n_9032));
XOR2_X1 i_9075 (.Z (n_9011), .A (n_9033), .B (n_9012));
INV_X1 i_9074 (.ZN (n_9010), .A (n_9011));
OR2_X1 i_9073 (.ZN (n_9009), .A1 (n_9010), .A2 (n_9014));
NAND2_X1 i_9072 (.ZN (n_9008), .A1 (n_9010), .A2 (n_9014));
INV_X1 i_9071 (.ZN (n_9007), .A (n_9008));
INV_X4 i_9070 (.ZN (n_9006), .A (B_imm[29]));
INV_X2 i_9069 (.ZN (n_9005), .A (A_imm[30]));
INV_X2 i_9068 (.ZN (n_9004), .A (B_imm[30]));
INV_X8 i_9067 (.ZN (n_9003), .A (B_imm[27]));
OAI22_X1 i_9066 (.ZN (n_9002), .A1 (n_9004), .A2 (n_9020), .B1 (CLOCK_opt_ipo_n433), .B2 (n_9037));
NAND2_X1 i_9065 (.ZN (n_9001), .A1 (B_imm[31]), .A2 (A_imm[27]));
INV_X1 i_9064 (.ZN (n_9000), .A (n_9001));
NAND4_X1 i_9063 (.ZN (n_8999), .A1 (B_imm[30]), .A2 (B_imm[27]), .A3 (opt_ipoPP_0), .A4 (A_imm[28]));
INV_X1 i_9062 (.ZN (n_8998), .A (n_8999));
OAI21_X1 i_9061 (.ZN (n_8997), .A (n_9002), .B1 (n_8998), .B2 (n_9000));
OAI21_X1 i_9060 (.ZN (n_8996), .A (n_8997), .B1 (n_9005), .B2 (n_9006));
OR3_X1 i_9059 (.ZN (n_8995), .A1 (n_8997), .A2 (n_9005), .A3 (n_9006));
INV_X4 i_9058 (.ZN (n_8994), .A (A_imm[29]));
INV_X4 i_9057 (.ZN (n_8993), .A (B_imm[26]));
OAI22_X1 i_9056 (.ZN (n_8992), .A1 (n_9020), .A2 (n_9006), .B1 (n_8993), .B2 (n_9037));
NAND2_X1 i_9055 (.ZN (n_8991), .A1 (B_imm[30]), .A2 (A_imm[27]));
INV_X1 i_9054 (.ZN (n_8990), .A (n_8991));
NAND4_X1 i_9053 (.ZN (n_8989), .A1 (A_imm[28]), .A2 (B_imm[29]), .A3 (B_imm[26]), .A4 (opt_ipoPP_0));
INV_X1 i_9052 (.ZN (n_8988), .A (n_8989));
OAI21_X1 i_9051 (.ZN (n_8987), .A (n_8992), .B1 (n_8990), .B2 (n_8988));
OAI21_X1 i_9050 (.ZN (n_8986), .A (n_8987), .B1 (n_9006), .B2 (n_8994));
NAND2_X1 i_9049 (.ZN (n_8985), .A1 (A_imm[30]), .A2 (B_imm[28]));
INV_X1 i_9048 (.ZN (n_8984), .A (n_8985));
OR3_X1 i_9047 (.ZN (n_8983), .A1 (n_8987), .A2 (n_9006), .A3 (n_8994));
INV_X1 i_9046 (.ZN (n_8982), .A (n_8983));
OAI21_X1 i_9045 (.ZN (n_8981), .A (n_8986), .B1 (n_8982), .B2 (n_8984));
NAND2_X1 i_9044 (.ZN (n_8980), .A1 (n_8981), .A2 (n_8995));
NAND2_X1 i_9043 (.ZN (n_8979), .A1 (n_8980), .A2 (n_8996));
OAI21_X1 i_9042 (.ZN (n_8978), .A (n_9009), .B1 (n_9007), .B2 (n_8979));
INV_X1 i_9041 (.ZN (n_8977), .A (n_8978));
NOR2_X1 i_9040 (.ZN (n_8976), .A1 (n_8977), .A2 (n_9022));
NAND2_X1 i_9039 (.ZN (n_8975), .A1 (n_8977), .A2 (n_9022));
INV_X2 i_9038 (.ZN (n_8974), .A (B_imm[25]));
INV_X2 i_9037 (.ZN (n_8973), .A (B_imm[13]));
INV_X4 i_9036 (.ZN (n_8972), .A (A_imm[26]));
INV_X4 i_9035 (.ZN (n_8971), .A (A_imm[14]));
OAI22_X1 i_9034 (.ZN (n_8970), .A1 (n_8974), .A2 (n_8971), .B1 (n_8973), .B2 (n_8972));
NAND2_X1 i_9033 (.ZN (n_8969), .A1 (B_imm[20]), .A2 (A_imm[19]));
NAND4_X1 i_9032 (.ZN (n_8968), .A1 (B_imm[25]), .A2 (B_imm[13]), .A3 (A_imm[26]), .A4 (A_imm[14]));
NAND2_X1 i_9031 (.ZN (n_8967), .A1 (n_8968), .A2 (n_8969));
AOI22_X1 i_9030 (.ZN (n_8966), .A1 (n_8967), .A2 (n_8970), .B1 (B_imm[30]), .B2 (A_imm[10]));
NAND4_X1 i_9029 (.ZN (n_8965), .A1 (n_8967), .A2 (n_8970), .A3 (B_imm[30]), .A4 (A_imm[10]));
INV_X1 i_9028 (.ZN (n_8964), .A (n_8965));
OAI211_X1 i_9027 (.ZN (n_8963), .A (B_imm[31]), .B (A_imm[9]), .C1 (n_8964), .C2 (n_8966));
NAND2_X1 i_9026 (.ZN (n_8962), .A1 (B_imm[31]), .A2 (A_imm[9]));
INV_X1 i_9025 (.ZN (n_8961), .A (n_8966));
NAND3_X1 i_9024 (.ZN (n_8960), .A1 (n_8961), .A2 (n_8962), .A3 (n_8965));
NAND2_X1 i_9023 (.ZN (n_8959), .A1 (n_8963), .A2 (n_8960));
INV_X4 i_9022 (.ZN (n_8958), .A (B_imm[22]));
INV_X2 i_9021 (.ZN (n_8957), .A (B_imm[21]));
INV_X4 i_9020 (.ZN (n_8956), .A (A_imm[18]));
INV_X2 i_9019 (.ZN (n_8955), .A (A_imm[17]));
OAI22_X1 i_9018 (.ZN (n_8954), .A1 (n_8958), .A2 (n_8955), .B1 (n_8957), .B2 (n_8956));
NAND2_X1 i_9017 (.ZN (n_8953), .A1 (B_imm[15]), .A2 (A_imm[24]));
INV_X1 i_9016 (.ZN (n_8952), .A (n_8953));
NAND4_X1 i_9015 (.ZN (n_8951), .A1 (B_imm[22]), .A2 (B_imm[21]), .A3 (A_imm[18]), .A4 (A_imm[17]));
INV_X1 i_9014 (.ZN (n_8950), .A (n_8951));
OAI21_X1 i_9013 (.ZN (n_8949), .A (n_8954), .B1 (n_8952), .B2 (n_8950));
INV_X4 i_9012 (.ZN (n_8948), .A (B_imm[24]));
INV_X4 i_9011 (.ZN (n_8947), .A (B_imm[8]));
INV_X4 i_9010 (.ZN (n_8946), .A (A_imm[15]));
OAI22_X1 i_9009 (.ZN (n_8945), .A1 (n_8948), .A2 (n_8946), .B1 (n_9037), .B2 (n_8947));
NAND2_X1 i_9008 (.ZN (n_8944), .A1 (B_imm[23]), .A2 (A_imm[16]));
INV_X1 i_9007 (.ZN (n_8943), .A (n_8944));
NAND4_X1 i_9006 (.ZN (n_8942), .A1 (B_imm[24]), .A2 (A_imm[31]), .A3 (B_imm[8]), .A4 (A_imm[15]));
INV_X1 i_9005 (.ZN (n_8941), .A (n_8942));
OAI21_X1 i_9004 (.ZN (n_8940), .A (n_8945), .B1 (n_8943), .B2 (n_8941));
NAND2_X1 i_9003 (.ZN (n_8939), .A1 (n_8949), .A2 (n_8940));
INV_X1 i_9002 (.ZN (n_8938), .A (n_8949));
INV_X1 i_9001 (.ZN (n_8937), .A (n_8940));
NAND2_X1 i_9000 (.ZN (n_8936), .A1 (n_8938), .A2 (n_8937));
NAND2_X1 i_8999 (.ZN (n_8935), .A1 (n_8936), .A2 (n_8939));
NAND3_X1 i_8998 (.ZN (n_8934), .A1 (n_8935), .A2 (B_imm[13]), .A3 (A_imm[27]));
NAND2_X1 i_8997 (.ZN (n_8933), .A1 (A_imm[27]), .A2 (B_imm[13]));
NAND3_X1 i_8996 (.ZN (n_8932), .A1 (n_8936), .A2 (n_8933), .A3 (n_8939));
NAND2_X1 i_8995 (.ZN (n_8931), .A1 (n_8934), .A2 (n_8932));
NAND2_X1 i_8994 (.ZN (n_8930), .A1 (n_8931), .A2 (n_8959));
NAND4_X1 i_8993 (.ZN (n_8929), .A1 (n_8934), .A2 (n_8963), .A3 (n_8960), .A4 (n_8932));
NAND2_X1 i_8992 (.ZN (n_8928), .A1 (B_imm[14]), .A2 (A_imm[26]));
INV_X4 i_8991 (.ZN (n_8927), .A (A_imm[13]));
INV_X8 i_8990 (.ZN (n_8926), .A (A_imm[11]));
OAI22_X1 i_8989 (.ZN (n_8925), .A1 (n_9021), .A2 (n_8926), .B1 (n_8993), .B2 (n_8927));
NAND2_X1 i_8988 (.ZN (n_8924), .A1 (B_imm[19]), .A2 (A_imm[20]));
INV_X1 i_8987 (.ZN (n_8923), .A (n_8924));
NAND4_X1 i_8986 (.ZN (n_8922), .A1 (B_imm[28]), .A2 (B_imm[26]), .A3 (A_imm[13]), .A4 (A_imm[11]));
INV_X1 i_8985 (.ZN (n_8921), .A (n_8922));
OAI21_X1 i_8984 (.ZN (n_8920), .A (n_8925), .B1 (n_8923), .B2 (n_8921));
NAND2_X1 i_8983 (.ZN (n_8919), .A1 (n_8920), .A2 (n_8928));
INV_X1 i_8982 (.ZN (n_8918), .A (n_8928));
INV_X1 i_8981 (.ZN (n_8917), .A (n_8920));
NAND2_X1 i_8980 (.ZN (n_8916), .A1 (n_8917), .A2 (n_8918));
NAND2_X1 i_8979 (.ZN (n_8915), .A1 (n_8916), .A2 (n_8919));
NAND3_X1 i_8978 (.ZN (n_8914), .A1 (n_8915), .A2 (B_imm[11]), .A3 (A_imm[29]));
NAND2_X1 i_8977 (.ZN (n_8913), .A1 (A_imm[29]), .A2 (B_imm[11]));
NAND3_X1 i_8976 (.ZN (n_8912), .A1 (n_8916), .A2 (n_8913), .A3 (n_8919));
NAND2_X1 i_8975 (.ZN (n_8911), .A1 (n_8914), .A2 (n_8912));
NAND2_X1 i_8974 (.ZN (n_8910), .A1 (n_8929), .A2 (n_8911));
INV_X8 i_8973 (.ZN (n_8909), .A (B_imm[17]));
INV_X4 i_8972 (.ZN (n_8908), .A (B_imm[16]));
INV_X8 i_8971 (.ZN (n_8907), .A (A_imm[23]));
INV_X4 i_8970 (.ZN (n_8906), .A (A_imm[22]));
OAI22_X1 i_8969 (.ZN (n_8905), .A1 (n_8907), .A2 (n_8908), .B1 (n_8909), .B2 (n_8906));
NAND2_X1 i_8968 (.ZN (n_8904), .A1 (B_imm[18]), .A2 (A_imm[21]));
NAND4_X1 i_8967 (.ZN (n_8903), .A1 (A_imm[23]), .A2 (B_imm[17]), .A3 (B_imm[16]), .A4 (A_imm[22]));
NAND2_X1 i_8966 (.ZN (n_8902), .A1 (n_8903), .A2 (n_8904));
NAND2_X1 i_8965 (.ZN (n_8901), .A1 (n_8902), .A2 (n_8905));
OAI21_X1 i_8964 (.ZN (n_8900), .A (n_8901), .B1 (n_9006), .B2 (n_8926));
NAND2_X1 i_8963 (.ZN (n_8899), .A1 (A_imm[28]), .A2 (B_imm[12]));
NAND4_X1 i_8962 (.ZN (n_8898), .A1 (n_8902), .A2 (n_8905), .A3 (B_imm[29]), .A4 (A_imm[11]));
NAND2_X1 i_8961 (.ZN (n_8897), .A1 (n_8898), .A2 (n_8899));
NAND2_X1 i_8960 (.ZN (n_8896), .A1 (n_8897), .A2 (n_8900));
NAND2_X1 i_8959 (.ZN (n_8895), .A1 (B_imm[15]), .A2 (A_imm[26]));
INV_X1 i_8958 (.ZN (n_8894), .A (n_8895));
INV_X4 i_8957 (.ZN (n_8893), .A (A_imm[20]));
INV_X2 i_8956 (.ZN (n_8892), .A (A_imm[19]));
OAI22_X1 i_8955 (.ZN (n_8891), .A1 (n_8958), .A2 (n_8892), .B1 (n_8957), .B2 (n_8893));
INV_X1 i_8954 (.ZN (n_8890), .A (n_8891));
NAND4_X1 i_8953 (.ZN (n_8889), .A1 (B_imm[22]), .A2 (B_imm[21]), .A3 (A_imm[20]), .A4 (A_imm[19]));
INV_X1 i_8952 (.ZN (n_8888), .A (n_8889));
OAI21_X1 i_8951 (.ZN (n_8887), .A (n_8894), .B1 (n_8890), .B2 (n_8888));
NAND3_X1 i_8950 (.ZN (n_8886), .A1 (n_8891), .A2 (n_8895), .A3 (n_8889));
NAND3_X1 i_8949 (.ZN (n_8885), .A1 (n_8896), .A2 (n_8887), .A3 (n_8886));
NAND2_X1 i_8948 (.ZN (n_8884), .A1 (n_8887), .A2 (n_8886));
NAND3_X1 i_8947 (.ZN (n_8883), .A1 (n_8884), .A2 (n_8900), .A3 (n_8897));
NAND2_X1 i_8946 (.ZN (n_8882), .A1 (n_8883), .A2 (n_8885));
NAND2_X1 i_8945 (.ZN (n_8881), .A1 (B_imm[23]), .A2 (A_imm[18]));
INV_X8 i_8944 (.ZN (n_8880), .A (B_imm[10]));
OAI22_X1 i_8943 (.ZN (n_8879), .A1 (n_8948), .A2 (n_8955), .B1 (n_9037), .B2 (n_8880));
NAND4_X1 i_8942 (.ZN (n_8878), .A1 (B_imm[24]), .A2 (A_imm[31]), .A3 (B_imm[10]), .A4 (A_imm[17]));
NAND2_X1 i_8941 (.ZN (n_8877), .A1 (n_8879), .A2 (n_8878));
INV_X1 i_8940 (.ZN (n_8876), .A (n_8877));
NOR2_X1 i_8939 (.ZN (n_8875), .A1 (n_8876), .A2 (n_8881));
NAND2_X1 i_8938 (.ZN (n_8874), .A1 (n_8876), .A2 (n_8881));
INV_X1 i_8937 (.ZN (n_8873), .A (n_8874));
NOR2_X1 i_8936 (.ZN (n_8872), .A1 (n_8875), .A2 (n_8873));
NAND2_X1 i_8935 (.ZN (n_8871), .A1 (n_8882), .A2 (n_8872));
INV_X1 i_8934 (.ZN (n_8870), .A (n_8872));
NAND3_X1 i_8933 (.ZN (n_8869), .A1 (n_8883), .A2 (n_8870), .A3 (n_8885));
NAND2_X1 i_8932 (.ZN (n_8868), .A1 (n_8871), .A2 (n_8869));
NAND3_X1 i_8931 (.ZN (n_8867), .A1 (n_8910), .A2 (n_8868), .A3 (n_8930));
NAND2_X1 i_8930 (.ZN (n_8866), .A1 (n_8910), .A2 (n_8930));
NAND3_X1 i_8929 (.ZN (n_8865), .A1 (n_8866), .A2 (n_8871), .A3 (n_8869));
NAND2_X1 i_8928 (.ZN (n_8864), .A1 (n_8916), .A2 (n_8913));
NAND2_X1 i_8927 (.ZN (n_8863), .A1 (n_8864), .A2 (n_8919));
NAND2_X1 i_8926 (.ZN (n_8862), .A1 (B_imm[28]), .A2 (A_imm[13]));
INV_X1 i_8925 (.ZN (n_8861), .A (n_8862));
INV_X4 i_8924 (.ZN (n_8860), .A (B_imm[20]));
INV_X4 i_8923 (.ZN (n_8859), .A (A_imm[21]));
INV_X4 i_8922 (.ZN (n_8858), .A (A_imm[16]));
OAI22_X1 i_8921 (.ZN (n_8857), .A1 (n_8860), .A2 (n_8859), .B1 (n_8974), .B2 (n_8858));
INV_X1 i_8920 (.ZN (n_8856), .A (n_8857));
NAND4_X1 i_8919 (.ZN (n_8855), .A1 (B_imm[20]), .A2 (B_imm[25]), .A3 (A_imm[21]), .A4 (A_imm[16]));
INV_X1 i_8918 (.ZN (n_8854), .A (n_8855));
OAI21_X1 i_8917 (.ZN (n_8853), .A (n_8861), .B1 (n_8856), .B2 (n_8854));
NAND3_X1 i_8916 (.ZN (n_8852), .A1 (n_8857), .A2 (n_8862), .A3 (n_8855));
NAND2_X1 i_8915 (.ZN (n_8851), .A1 (n_8853), .A2 (n_8852));
NAND3_X1 i_8914 (.ZN (n_8850), .A1 (n_8851), .A2 (B_imm[11]), .A3 (A_imm[30]));
INV_X8 i_8913 (.ZN (n_8849), .A (B_imm[11]));
OAI211_X1 i_8912 (.ZN (n_8848), .A (n_8853), .B (n_8852), .C1 (n_9005), .C2 (n_8849));
NAND3_X1 i_8911 (.ZN (n_8847), .A1 (n_8863), .A2 (n_8850), .A3 (n_8848));
NAND2_X1 i_8910 (.ZN (n_8846), .A1 (n_8848), .A2 (n_8850));
NAND3_X1 i_8909 (.ZN (n_8845), .A1 (n_8846), .A2 (n_8919), .A3 (n_8864));
NAND2_X1 i_8908 (.ZN (n_8844), .A1 (n_8845), .A2 (n_8847));
NAND3_X1 i_8907 (.ZN (n_8843), .A1 (n_8865), .A2 (n_8867), .A3 (n_8844));
NAND2_X1 i_8906 (.ZN (n_8842), .A1 (n_8865), .A2 (n_8867));
INV_X1 i_8905 (.ZN (n_8841), .A (n_8844));
NAND2_X1 i_8904 (.ZN (n_8840), .A1 (n_8842), .A2 (n_8841));
NAND2_X1 i_8903 (.ZN (n_8839), .A1 (n_8840), .A2 (n_8843));
NAND2_X1 i_8902 (.ZN (n_8838), .A1 (n_8970), .A2 (n_8968));
NAND3_X1 i_8901 (.ZN (n_8837), .A1 (n_8838), .A2 (B_imm[20]), .A3 (A_imm[19]));
NAND3_X1 i_8900 (.ZN (n_8836), .A1 (n_8970), .A2 (n_8969), .A3 (n_8968));
NAND2_X1 i_8899 (.ZN (n_8835), .A1 (n_8837), .A2 (n_8836));
INV_X1 i_8898 (.ZN (n_8834), .A (n_8925));
OAI21_X1 i_8897 (.ZN (n_8833), .A (n_8923), .B1 (n_8834), .B2 (n_8921));
NAND3_X1 i_8896 (.ZN (n_8832), .A1 (n_8925), .A2 (n_8924), .A3 (n_8922));
NAND2_X1 i_8895 (.ZN (n_8831), .A1 (n_8833), .A2 (n_8832));
NAND2_X1 i_8894 (.ZN (n_8830), .A1 (n_8831), .A2 (n_8835));
INV_X4 i_8893 (.ZN (n_8829), .A (B_imm[15]));
NAND2_X1 i_8892 (.ZN (n_8828), .A1 (B_imm[22]), .A2 (A_imm[15]));
OAI21_X1 i_8891 (.ZN (n_8827), .A (n_8828), .B1 (n_8829), .B2 (n_8906));
NAND2_X1 i_8890 (.ZN (n_8826), .A1 (B_imm[25]), .A2 (A_imm[12]));
INV_X1 i_8889 (.ZN (n_8825), .A (n_8826));
NAND4_X1 i_8888 (.ZN (n_8824), .A1 (B_imm[15]), .A2 (B_imm[22]), .A3 (A_imm[22]), .A4 (A_imm[15]));
INV_X1 i_8887 (.ZN (n_8823), .A (n_8824));
OAI21_X1 i_8886 (.ZN (n_8822), .A (n_8827), .B1 (n_8823), .B2 (n_8825));
INV_X2 i_8885 (.ZN (n_8821), .A (B_imm[23]));
NAND2_X1 i_8884 (.ZN (n_8820), .A1 (A_imm[31]), .A2 (B_imm[6]));
OAI21_X1 i_8883 (.ZN (n_8819), .A (n_8820), .B1 (n_8821), .B2 (n_8971));
NAND2_X1 i_8882 (.ZN (n_8818), .A1 (B_imm[21]), .A2 (A_imm[16]));
INV_X1 i_8881 (.ZN (n_8817), .A (n_8818));
NAND4_X1 i_8880 (.ZN (n_8816), .A1 (B_imm[23]), .A2 (A_imm[31]), .A3 (B_imm[6]), .A4 (A_imm[14]));
INV_X1 i_8879 (.ZN (n_8815), .A (n_8816));
OAI21_X1 i_8878 (.ZN (n_8814), .A (n_8819), .B1 (n_8815), .B2 (n_8817));
NAND2_X1 i_8877 (.ZN (n_8813), .A1 (n_8822), .A2 (n_8814));
NAND2_X1 i_8876 (.ZN (n_8812), .A1 (A_imm[27]), .A2 (B_imm[11]));
INV_X1 i_8875 (.ZN (n_8811), .A (n_8812));
INV_X1 i_8874 (.ZN (n_8810), .A (n_8822));
INV_X1 i_8873 (.ZN (n_8809), .A (n_8814));
NAND2_X1 i_8872 (.ZN (n_8808), .A1 (n_8810), .A2 (n_8809));
INV_X1 i_8871 (.ZN (n_8807), .A (n_8808));
OAI21_X1 i_8870 (.ZN (n_8806), .A (n_8813), .B1 (n_8807), .B2 (n_8811));
NAND4_X1 i_8869 (.ZN (n_8805), .A1 (n_8833), .A2 (n_8837), .A3 (n_8836), .A4 (n_8832));
INV_X1 i_8868 (.ZN (n_8804), .A (n_8805));
OAI21_X1 i_8867 (.ZN (n_8803), .A (n_8830), .B1 (n_8804), .B2 (n_8806));
OAI22_X1 i_8866 (.ZN (n_8802), .A1 (n_8893), .A2 (n_8909), .B1 (n_8859), .B2 (n_8908));
NAND2_X1 i_8865 (.ZN (n_8801), .A1 (B_imm[18]), .A2 (A_imm[19]));
INV_X1 i_8864 (.ZN (n_8800), .A (n_8801));
NAND4_X1 i_8863 (.ZN (n_8799), .A1 (A_imm[20]), .A2 (B_imm[17]), .A3 (B_imm[16]), .A4 (A_imm[21]));
INV_X1 i_8862 (.ZN (n_8798), .A (n_8799));
OAI21_X1 i_8861 (.ZN (n_8797), .A (n_8802), .B1 (n_8800), .B2 (n_8798));
OAI21_X1 i_8860 (.ZN (n_8796), .A (n_8797), .B1 (n_8880), .B2 (n_9020));
INV_X4 i_8859 (.ZN (n_8795), .A (B_imm[12]));
INV_X4 i_8858 (.ZN (n_8794), .A (A_imm[25]));
NAND2_X1 i_8857 (.ZN (n_8793), .A1 (A_imm[26]), .A2 (B_imm[11]));
OAI21_X1 i_8856 (.ZN (n_8792), .A (n_8793), .B1 (n_8794), .B2 (n_8795));
NAND2_X1 i_8855 (.ZN (n_8791), .A1 (B_imm[24]), .A2 (A_imm[13]));
INV_X1 i_8854 (.ZN (n_8790), .A (n_8791));
NAND4_X1 i_8853 (.ZN (n_8789), .A1 (A_imm[26]), .A2 (A_imm[25]), .A3 (B_imm[11]), .A4 (B_imm[12]));
INV_X1 i_8852 (.ZN (n_8788), .A (n_8789));
OAI21_X1 i_8851 (.ZN (n_8787), .A (n_8792), .B1 (n_8788), .B2 (n_8790));
INV_X1 i_8850 (.ZN (n_8786), .A (n_8797));
NAND3_X1 i_8849 (.ZN (n_8785), .A1 (n_8786), .A2 (B_imm[10]), .A3 (A_imm[28]));
NAND2_X1 i_8848 (.ZN (n_8784), .A1 (n_8785), .A2 (n_8787));
AOI21_X1 i_8847 (.ZN (n_8783), .A (n_8953), .B1 (n_8954), .B2 (n_8951));
NAND3_X1 i_8846 (.ZN (n_8782), .A1 (n_8954), .A2 (n_8953), .A3 (n_8951));
INV_X1 i_8845 (.ZN (n_8781), .A (n_8782));
OAI211_X1 i_8844 (.ZN (n_8780), .A (n_8784), .B (n_8796), .C1 (n_8783), .C2 (n_8781));
NAND2_X1 i_8843 (.ZN (n_8779), .A1 (n_8784), .A2 (n_8796));
NOR2_X1 i_8842 (.ZN (n_8778), .A1 (n_8783), .A2 (n_8781));
NAND2_X1 i_8841 (.ZN (n_8777), .A1 (n_8779), .A2 (n_8778));
NAND2_X1 i_8840 (.ZN (n_8776), .A1 (n_8945), .A2 (n_8942));
XNOR2_X1 i_8839 (.ZN (n_8775), .A (n_8776), .B (n_8943));
NAND2_X1 i_8838 (.ZN (n_8774), .A1 (n_8777), .A2 (n_8775));
NAND2_X1 i_8837 (.ZN (n_8773), .A1 (n_8774), .A2 (n_8780));
NAND2_X1 i_8836 (.ZN (n_8772), .A1 (n_8773), .A2 (n_8803));
NAND2_X1 i_8835 (.ZN (n_8771), .A1 (n_8808), .A2 (n_8812));
NAND3_X1 i_8834 (.ZN (n_8770), .A1 (n_8805), .A2 (n_8813), .A3 (n_8771));
NAND4_X1 i_8833 (.ZN (n_8769), .A1 (n_8770), .A2 (n_8774), .A3 (n_8830), .A4 (n_8780));
NAND2_X1 i_8832 (.ZN (n_8768), .A1 (B_imm[30]), .A2 (A_imm[8]));
INV_X4 i_8831 (.ZN (n_8767), .A (A_imm[24]));
OAI22_X1 i_8830 (.ZN (n_8766), .A1 (n_8860), .A2 (n_8955), .B1 (n_8973), .B2 (n_8767));
NAND2_X1 i_8829 (.ZN (n_8765), .A1 (B_imm[28]), .A2 (A_imm[9]));
NAND4_X1 i_8828 (.ZN (n_8764), .A1 (B_imm[20]), .A2 (B_imm[13]), .A3 (A_imm[24]), .A4 (A_imm[17]));
NAND2_X1 i_8827 (.ZN (n_8763), .A1 (n_8764), .A2 (n_8765));
NAND2_X1 i_8826 (.ZN (n_8762), .A1 (n_8763), .A2 (n_8766));
NAND2_X1 i_8825 (.ZN (n_8761), .A1 (n_8762), .A2 (n_8768));
NAND2_X1 i_8824 (.ZN (n_8760), .A1 (B_imm[31]), .A2 (A_imm[7]));
NAND4_X1 i_8823 (.ZN (n_8759), .A1 (n_8763), .A2 (n_8766), .A3 (B_imm[30]), .A4 (A_imm[8]));
NAND2_X1 i_8822 (.ZN (n_8758), .A1 (n_8759), .A2 (n_8760));
NAND4_X1 i_8821 (.ZN (n_8757), .A1 (n_8758), .A2 (B_imm[9]), .A3 (A_imm[30]), .A4 (n_8761));
INV_X1 i_8820 (.ZN (n_8756), .A (n_8757));
NAND2_X1 i_8819 (.ZN (n_8755), .A1 (A_imm[30]), .A2 (B_imm[9]));
NAND2_X1 i_8818 (.ZN (n_8754), .A1 (n_8758), .A2 (n_8761));
NAND2_X1 i_8817 (.ZN (n_8753), .A1 (n_8754), .A2 (n_8755));
INV_X2 i_8816 (.ZN (n_8752), .A (A_imm[12]));
INV_X4 i_8815 (.ZN (n_8751), .A (A_imm[10]));
OAI22_X1 i_8814 (.ZN (n_8750), .A1 (n_9006), .A2 (n_8751), .B1 (n_9003), .B2 (n_8752));
NAND4_X1 i_8813 (.ZN (n_8749), .A1 (B_imm[29]), .A2 (B_imm[27]), .A3 (A_imm[12]), .A4 (A_imm[10]));
NAND2_X1 i_8812 (.ZN (n_8748), .A1 (n_8750), .A2 (n_8749));
OAI22_X1 i_8811 (.ZN (n_8747), .A1 (n_8908), .A2 (n_8906), .B1 (n_8859), .B2 (n_8909));
NAND2_X1 i_8810 (.ZN (n_8746), .A1 (B_imm[18]), .A2 (A_imm[20]));
INV_X1 i_8809 (.ZN (n_8745), .A (n_8746));
NAND4_X1 i_8808 (.ZN (n_8744), .A1 (A_imm[21]), .A2 (A_imm[22]), .A3 (B_imm[16]), .A4 (B_imm[17]));
INV_X1 i_8807 (.ZN (n_8743), .A (n_8744));
OAI21_X1 i_8806 (.ZN (n_8742), .A (n_8747), .B1 (n_8745), .B2 (n_8743));
XNOR2_X1 i_8805 (.ZN (n_8741), .A (n_8748), .B (n_8742));
INV_X1 i_8804 (.ZN (n_8740), .A (n_8741));
AOI21_X1 i_8803 (.ZN (n_8739), .A (n_8756), .B1 (n_8740), .B2 (n_8753));
INV_X1 i_8802 (.ZN (n_8738), .A (n_8739));
NAND3_X1 i_8801 (.ZN (n_8737), .A1 (n_8772), .A2 (n_8769), .A3 (n_8738));
NAND2_X1 i_8800 (.ZN (n_8736), .A1 (n_8769), .A2 (n_8772));
NAND2_X1 i_8799 (.ZN (n_8735), .A1 (n_8736), .A2 (n_8739));
NAND2_X1 i_8798 (.ZN (n_8734), .A1 (B_imm[29]), .A2 (A_imm[9]));
INV_X1 i_8797 (.ZN (n_8733), .A (n_8734));
NAND2_X1 i_8796 (.ZN (n_8732), .A1 (B_imm[19]), .A2 (A_imm[19]));
OAI21_X1 i_8795 (.ZN (n_8731), .A (n_8732), .B1 (n_9003), .B2 (n_8926));
NAND4_X1 i_8794 (.ZN (n_8730), .A1 (B_imm[27]), .A2 (B_imm[19]), .A3 (A_imm[19]), .A4 (A_imm[11]));
NAND2_X1 i_8793 (.ZN (n_8729), .A1 (n_8731), .A2 (n_8730));
NAND2_X1 i_8792 (.ZN (n_8728), .A1 (n_8729), .A2 (n_8733));
NAND3_X1 i_8791 (.ZN (n_8727), .A1 (n_8731), .A2 (n_8734), .A3 (n_8730));
NAND2_X1 i_8790 (.ZN (n_8726), .A1 (n_8728), .A2 (n_8727));
NAND2_X1 i_8789 (.ZN (n_8725), .A1 (B_imm[26]), .A2 (A_imm[12]));
INV_X1 i_8788 (.ZN (n_8724), .A (n_8725));
NAND2_X1 i_8787 (.ZN (n_8723), .A1 (B_imm[20]), .A2 (A_imm[18]));
OAI21_X1 i_8786 (.ZN (n_8722), .A (n_8723), .B1 (n_9021), .B2 (n_8751));
NAND4_X1 i_8785 (.ZN (n_8721), .A1 (B_imm[28]), .A2 (B_imm[20]), .A3 (A_imm[18]), .A4 (A_imm[10]));
NAND2_X1 i_8784 (.ZN (n_8720), .A1 (n_8722), .A2 (n_8721));
NAND2_X1 i_8783 (.ZN (n_8719), .A1 (n_8720), .A2 (n_8724));
NAND3_X1 i_8782 (.ZN (n_8718), .A1 (n_8722), .A2 (n_8725), .A3 (n_8721));
NAND2_X1 i_8781 (.ZN (n_8717), .A1 (n_8719), .A2 (n_8718));
NAND2_X1 i_8780 (.ZN (n_8716), .A1 (n_8726), .A2 (n_8717));
NAND4_X1 i_8779 (.ZN (n_8715), .A1 (n_8728), .A2 (n_8719), .A3 (n_8727), .A4 (n_8718));
NAND2_X1 i_8778 (.ZN (n_8714), .A1 (A_imm[27]), .A2 (B_imm[10]));
NAND2_X1 i_8777 (.ZN (n_8713), .A1 (B_imm[13]), .A2 (A_imm[23]));
OAI21_X1 i_8776 (.ZN (n_8712), .A (n_8713), .B1 (n_8974), .B2 (n_8926));
NAND2_X1 i_8775 (.ZN (n_8711), .A1 (B_imm[20]), .A2 (A_imm[16]));
INV_X1 i_8774 (.ZN (n_8710), .A (n_8711));
NAND4_X1 i_8773 (.ZN (n_8709), .A1 (B_imm[25]), .A2 (B_imm[13]), .A3 (A_imm[23]), .A4 (A_imm[11]));
INV_X1 i_8772 (.ZN (n_8708), .A (n_8709));
OAI21_X1 i_8771 (.ZN (n_8707), .A (n_8712), .B1 (n_8708), .B2 (n_8710));
NAND2_X1 i_8770 (.ZN (n_8706), .A1 (n_8707), .A2 (n_8714));
NAND2_X1 i_8769 (.ZN (n_8705), .A1 (n_8709), .A2 (n_8711));
NAND4_X1 i_8768 (.ZN (n_8704), .A1 (n_8705), .A2 (B_imm[10]), .A3 (A_imm[27]), .A4 (n_8712));
NAND2_X1 i_8767 (.ZN (n_8703), .A1 (B_imm[30]), .A2 (A_imm[7]));
NAND2_X1 i_8766 (.ZN (n_8702), .A1 (n_8704), .A2 (n_8703));
NAND3_X1 i_8765 (.ZN (n_8701), .A1 (n_8715), .A2 (n_8706), .A3 (n_8702));
NAND2_X1 i_8764 (.ZN (n_8700), .A1 (n_8701), .A2 (n_8716));
NAND2_X1 i_8763 (.ZN (n_8699), .A1 (n_8730), .A2 (n_8734));
NAND4_X1 i_8762 (.ZN (n_8698), .A1 (n_8699), .A2 (A_imm[29]), .A3 (B_imm[10]), .A4 (n_8731));
NAND2_X1 i_8761 (.ZN (n_8697), .A1 (n_8699), .A2 (n_8731));
OAI21_X1 i_8760 (.ZN (n_8696), .A (n_8697), .B1 (n_8880), .B2 (n_8994));
INV_X1 i_8759 (.ZN (n_8695), .A (n_8904));
NAND2_X1 i_8758 (.ZN (n_8694), .A1 (n_8905), .A2 (n_8903));
XNOR2_X1 i_8757 (.ZN (n_8693), .A (n_8694), .B (n_8695));
INV_X1 i_8756 (.ZN (n_8692), .A (n_8693));
NAND3_X1 i_8755 (.ZN (n_8691), .A1 (n_8696), .A2 (n_8692), .A3 (n_8698));
NAND2_X1 i_8754 (.ZN (n_8690), .A1 (n_8696), .A2 (n_8698));
NAND2_X1 i_8753 (.ZN (n_8689), .A1 (n_8690), .A2 (n_8693));
NAND2_X1 i_8752 (.ZN (n_8688), .A1 (n_8689), .A2 (n_8691));
NAND2_X1 i_8751 (.ZN (n_8687), .A1 (n_8688), .A2 (n_8700));
NAND4_X1 i_8750 (.ZN (n_8686), .A1 (n_8689), .A2 (n_8701), .A3 (n_8716), .A4 (n_8691));
NAND2_X1 i_8749 (.ZN (n_8685), .A1 (B_imm[31]), .A2 (A_imm[6]));
NAND2_X1 i_8748 (.ZN (n_8684), .A1 (B_imm[28]), .A2 (A_imm[8]));
OAI21_X1 i_8747 (.ZN (n_8683), .A (n_8684), .B1 (n_8993), .B2 (n_8751));
NAND2_X1 i_8746 (.ZN (n_8682), .A1 (B_imm[19]), .A2 (A_imm[17]));
NAND4_X1 i_8745 (.ZN (n_8681), .A1 (B_imm[28]), .A2 (B_imm[26]), .A3 (A_imm[10]), .A4 (A_imm[8]));
NAND2_X1 i_8744 (.ZN (n_8680), .A1 (n_8681), .A2 (n_8682));
NAND2_X1 i_8743 (.ZN (n_8679), .A1 (n_8680), .A2 (n_8683));
NAND2_X1 i_8742 (.ZN (n_8678), .A1 (n_8679), .A2 (n_8685));
NAND4_X1 i_8741 (.ZN (n_8677), .A1 (n_8680), .A2 (B_imm[31]), .A3 (A_imm[6]), .A4 (n_8683));
NAND2_X1 i_8740 (.ZN (n_8676), .A1 (B_imm[14]), .A2 (A_imm[23]));
NAND2_X1 i_8739 (.ZN (n_8675), .A1 (n_8677), .A2 (n_8676));
NAND4_X1 i_8738 (.ZN (n_8674), .A1 (n_8675), .A2 (B_imm[8]), .A3 (A_imm[30]), .A4 (n_8678));
AOI22_X1 i_8737 (.ZN (n_8673), .A1 (n_8675), .A2 (n_8678), .B1 (A_imm[30]), .B2 (B_imm[8]));
AOI21_X1 i_8736 (.ZN (n_8672), .A (n_8787), .B1 (n_8796), .B2 (n_8785));
NAND3_X1 i_8735 (.ZN (n_8671), .A1 (n_8785), .A2 (n_8796), .A3 (n_8787));
INV_X1 i_8734 (.ZN (n_8670), .A (n_8671));
NOR2_X1 i_8733 (.ZN (n_8669), .A1 (n_8670), .A2 (n_8672));
OAI21_X1 i_8732 (.ZN (n_8668), .A (n_8674), .B1 (n_8673), .B2 (n_8669));
NAND2_X1 i_8731 (.ZN (n_8667), .A1 (n_8686), .A2 (n_8668));
NAND2_X1 i_8730 (.ZN (n_8666), .A1 (n_8667), .A2 (n_8687));
NAND3_X1 i_8729 (.ZN (n_8665), .A1 (n_8735), .A2 (n_8737), .A3 (n_8666));
NAND2_X1 i_8728 (.ZN (n_8664), .A1 (n_8735), .A2 (n_8737));
INV_X1 i_8727 (.ZN (n_8663), .A (n_8666));
NAND2_X1 i_8726 (.ZN (n_8662), .A1 (n_8664), .A2 (n_8663));
NAND2_X1 i_8725 (.ZN (n_8661), .A1 (n_8930), .A2 (n_8929));
XNOR2_X1 i_8724 (.ZN (n_8660), .A (n_8661), .B (n_8911));
NAND2_X1 i_8723 (.ZN (n_8659), .A1 (n_8662), .A2 (n_8660));
NAND3_X1 i_8722 (.ZN (n_8658), .A1 (n_8839), .A2 (n_8659), .A3 (n_8665));
NAND2_X1 i_8721 (.ZN (n_8657), .A1 (n_8659), .A2 (n_8665));
NAND3_X1 i_8720 (.ZN (n_8656), .A1 (n_8657), .A2 (n_8843), .A3 (n_8840));
NAND2_X1 i_8719 (.ZN (n_8655), .A1 (n_8656), .A2 (n_8658));
AOI21_X1 i_8718 (.ZN (n_8654), .A (n_8812), .B1 (n_8813), .B2 (n_8808));
INV_X1 i_8717 (.ZN (n_8653), .A (n_8654));
NAND3_X1 i_8716 (.ZN (n_8652), .A1 (n_8808), .A2 (n_8813), .A3 (n_8812));
NAND2_X1 i_8715 (.ZN (n_8651), .A1 (n_8802), .A2 (n_8799));
NAND2_X1 i_8714 (.ZN (n_8650), .A1 (n_8651), .A2 (n_8800));
NAND3_X1 i_8713 (.ZN (n_8649), .A1 (n_8802), .A2 (n_8801), .A3 (n_8799));
OAI211_X1 i_8712 (.ZN (n_8648), .A (n_8650), .B (n_8649), .C1 (n_8994), .C2 (n_8947));
NAND2_X1 i_8711 (.ZN (n_8647), .A1 (n_8650), .A2 (n_8649));
NAND3_X1 i_8710 (.ZN (n_8646), .A1 (n_8647), .A2 (B_imm[8]), .A3 (A_imm[29]));
INV_X4 i_8709 (.ZN (n_8645), .A (A_imm[9]));
INV_X2 i_8708 (.ZN (n_8644), .A (A_imm[7]));
OAI22_X1 i_8707 (.ZN (n_8643), .A1 (n_9006), .A2 (n_8644), .B1 (n_9003), .B2 (n_8645));
NAND2_X1 i_8706 (.ZN (n_8642), .A1 (B_imm[16]), .A2 (A_imm[19]));
NAND2_X1 i_8705 (.ZN (n_8641), .A1 (A_imm[18]), .A2 (B_imm[17]));
NAND2_X1 i_8704 (.ZN (n_8640), .A1 (n_8641), .A2 (n_8642));
NAND2_X1 i_8703 (.ZN (n_8639), .A1 (B_imm[12]), .A2 (A_imm[23]));
INV_X1 i_8702 (.ZN (n_8638), .A (n_8639));
NAND4_X1 i_8701 (.ZN (n_8637), .A1 (A_imm[18]), .A2 (B_imm[16]), .A3 (B_imm[17]), .A4 (A_imm[19]));
INV_X1 i_8700 (.ZN (n_8636), .A (n_8637));
OAI21_X1 i_8699 (.ZN (n_8635), .A (n_8640), .B1 (n_8638), .B2 (n_8636));
INV_X1 i_8698 (.ZN (n_8634), .A (n_8635));
NAND4_X1 i_8697 (.ZN (n_8633), .A1 (B_imm[29]), .A2 (B_imm[27]), .A3 (A_imm[9]), .A4 (A_imm[7]));
INV_X1 i_8696 (.ZN (n_8632), .A (n_8633));
OAI21_X1 i_8695 (.ZN (n_8631), .A (n_8643), .B1 (n_8634), .B2 (n_8632));
NAND2_X1 i_8694 (.ZN (n_8630), .A1 (n_8646), .A2 (n_8631));
NAND2_X1 i_8693 (.ZN (n_8629), .A1 (n_8630), .A2 (n_8648));
NAND3_X1 i_8692 (.ZN (n_8628), .A1 (n_8653), .A2 (n_8629), .A3 (n_8652));
INV_X1 i_8691 (.ZN (n_8627), .A (n_8652));
INV_X1 i_8690 (.ZN (n_8626), .A (n_8629));
OAI21_X1 i_8689 (.ZN (n_8625), .A (n_8626), .B1 (n_8627), .B2 (n_8654));
INV_X1 i_8688 (.ZN (n_8624), .A (n_8819));
OAI21_X1 i_8687 (.ZN (n_8623), .A (n_8817), .B1 (n_8624), .B2 (n_8815));
NAND3_X1 i_8686 (.ZN (n_8622), .A1 (n_8819), .A2 (n_8818), .A3 (n_8816));
NAND2_X1 i_8685 (.ZN (n_8621), .A1 (n_8623), .A2 (n_8622));
INV_X1 i_8684 (.ZN (n_8620), .A (n_8792));
OAI21_X1 i_8683 (.ZN (n_8619), .A (n_8790), .B1 (n_8620), .B2 (n_8788));
NAND3_X1 i_8682 (.ZN (n_8618), .A1 (n_8792), .A2 (n_8791), .A3 (n_8789));
NAND2_X1 i_8681 (.ZN (n_8617), .A1 (n_8619), .A2 (n_8618));
NAND2_X1 i_8680 (.ZN (n_8616), .A1 (n_8621), .A2 (n_8617));
NAND4_X1 i_8679 (.ZN (n_8615), .A1 (n_8623), .A2 (n_8619), .A3 (n_8622), .A4 (n_8618));
NAND2_X1 i_8678 (.ZN (n_8614), .A1 (B_imm[11]), .A2 (A_imm[24]));
OAI21_X1 i_8677 (.ZN (n_8613), .A (n_8614), .B1 (n_8794), .B2 (n_8880));
NAND2_X1 i_8676 (.ZN (n_8612), .A1 (B_imm[18]), .A2 (A_imm[17]));
NAND4_X1 i_8675 (.ZN (n_8611), .A1 (A_imm[25]), .A2 (B_imm[11]), .A3 (B_imm[10]), .A4 (A_imm[24]));
NAND2_X1 i_8674 (.ZN (n_8610), .A1 (n_8611), .A2 (n_8612));
AOI22_X1 i_8673 (.ZN (n_8609), .A1 (n_8610), .A2 (n_8613), .B1 (A_imm[28]), .B2 (B_imm[8]));
INV_X1 i_8672 (.ZN (n_8608), .A (n_8609));
NAND4_X1 i_8671 (.ZN (n_8607), .A1 (n_8610), .A2 (B_imm[8]), .A3 (A_imm[28]), .A4 (n_8613));
NAND2_X1 i_8670 (.ZN (n_8606), .A1 (B_imm[9]), .A2 (A_imm[26]));
OAI21_X1 i_8669 (.ZN (n_8605), .A (n_8606), .B1 (n_8948), .B2 (n_8926));
NAND2_X1 i_8668 (.ZN (n_8604), .A1 (A_imm[31]), .A2 (B_imm[4]));
INV_X1 i_8667 (.ZN (n_8603), .A (n_8604));
NAND4_X1 i_8666 (.ZN (n_8602), .A1 (B_imm[24]), .A2 (B_imm[9]), .A3 (A_imm[26]), .A4 (A_imm[11]));
INV_X1 i_8665 (.ZN (n_8601), .A (n_8602));
OAI21_X1 i_8664 (.ZN (n_8600), .A (n_8605), .B1 (n_8601), .B2 (n_8603));
NAND2_X1 i_8663 (.ZN (n_8599), .A1 (n_8607), .A2 (n_8600));
NAND2_X1 i_8662 (.ZN (n_8598), .A1 (n_8599), .A2 (n_8608));
INV_X1 i_8661 (.ZN (n_8597), .A (n_8598));
NAND2_X1 i_8660 (.ZN (n_8596), .A1 (n_8597), .A2 (n_8615));
NAND2_X1 i_8659 (.ZN (n_8595), .A1 (n_8596), .A2 (n_8616));
INV_X1 i_8658 (.ZN (n_8594), .A (n_8595));
NAND2_X1 i_8657 (.ZN (n_8593), .A1 (n_8594), .A2 (n_8625));
NAND2_X1 i_8656 (.ZN (n_8592), .A1 (n_8593), .A2 (n_8628));
NAND2_X1 i_8655 (.ZN (n_8591), .A1 (n_8753), .A2 (n_8757));
NAND2_X1 i_8654 (.ZN (n_8590), .A1 (n_8591), .A2 (n_8741));
NAND3_X1 i_8653 (.ZN (n_8589), .A1 (n_8753), .A2 (n_8740), .A3 (n_8757));
NAND2_X1 i_8652 (.ZN (n_8588), .A1 (n_8590), .A2 (n_8589));
NAND2_X1 i_8651 (.ZN (n_8587), .A1 (n_8588), .A2 (n_8592));
NAND4_X2 i_8650 (.ZN (n_8586), .A1 (n_8590), .A2 (n_8593), .A3 (n_8628), .A4 (n_8589));
NAND2_X1 i_8649 (.ZN (n_8585), .A1 (n_8777), .A2 (n_8780));
XNOR2_X1 i_8648 (.ZN (n_8584), .A (n_8585), .B (n_8775));
INV_X1 i_8647 (.ZN (n_8583), .A (n_8584));
NAND2_X1 i_8646 (.ZN (n_8582), .A1 (n_8586), .A2 (n_8583));
NAND2_X1 i_8645 (.ZN (n_8581), .A1 (n_8830), .A2 (n_8805));
NAND3_X1 i_8644 (.ZN (n_8580), .A1 (n_8581), .A2 (n_8813), .A3 (n_8771));
NAND3_X1 i_8643 (.ZN (n_8579), .A1 (n_8806), .A2 (n_8830), .A3 (n_8805));
NAND2_X1 i_8642 (.ZN (n_8578), .A1 (n_8759), .A2 (n_8761));
NAND3_X1 i_8641 (.ZN (n_8577), .A1 (n_8578), .A2 (B_imm[31]), .A3 (A_imm[7]));
NAND3_X1 i_8640 (.ZN (n_8576), .A1 (n_8761), .A2 (n_8759), .A3 (n_8760));
NAND2_X1 i_8639 (.ZN (n_8575), .A1 (n_8577), .A2 (n_8576));
INV_X1 i_8638 (.ZN (n_8574), .A (n_8575));
INV_X2 i_8637 (.ZN (n_8573), .A (B_imm[7]));
INV_X1 i_8636 (.ZN (n_8572), .A (n_8765));
NAND2_X1 i_8635 (.ZN (n_8571), .A1 (n_8766), .A2 (n_8764));
NAND2_X1 i_8634 (.ZN (n_8570), .A1 (n_8571), .A2 (n_8572));
NAND3_X1 i_8633 (.ZN (n_8569), .A1 (n_8766), .A2 (n_8765), .A3 (n_8764));
OAI211_X1 i_8632 (.ZN (n_8568), .A (n_8570), .B (n_8569), .C1 (n_9005), .C2 (n_8573));
NAND2_X1 i_8631 (.ZN (n_8567), .A1 (n_8570), .A2 (n_8569));
NAND3_X1 i_8630 (.ZN (n_8566), .A1 (n_8567), .A2 (B_imm[7]), .A3 (A_imm[30]));
NAND2_X1 i_8629 (.ZN (n_8565), .A1 (B_imm[20]), .A2 (A_imm[15]));
NAND2_X1 i_8628 (.ZN (n_8564), .A1 (B_imm[28]), .A2 (A_imm[7]));
NAND2_X1 i_8627 (.ZN (n_8563), .A1 (n_8564), .A2 (n_8565));
NAND2_X1 i_8626 (.ZN (n_8562), .A1 (B_imm[26]), .A2 (A_imm[9]));
NAND4_X1 i_8625 (.ZN (n_8561), .A1 (B_imm[28]), .A2 (B_imm[20]), .A3 (A_imm[15]), .A4 (A_imm[7]));
NAND2_X1 i_8624 (.ZN (n_8560), .A1 (n_8561), .A2 (n_8562));
AOI22_X1 i_8623 (.ZN (n_8559), .A1 (n_8560), .A2 (n_8563), .B1 (B_imm[30]), .B2 (A_imm[6]));
INV_X1 i_8622 (.ZN (n_8558), .A (n_8559));
NAND4_X1 i_8621 (.ZN (n_8557), .A1 (n_8560), .A2 (B_imm[30]), .A3 (A_imm[6]), .A4 (n_8563));
INV_X1 i_8620 (.ZN (n_8556), .A (n_8557));
NAND2_X1 i_8619 (.ZN (n_8555), .A1 (B_imm[31]), .A2 (A_imm[5]));
INV_X1 i_8618 (.ZN (n_8554), .A (n_8555));
OAI21_X1 i_8617 (.ZN (n_8553), .A (n_8558), .B1 (n_8556), .B2 (n_8554));
NAND2_X1 i_8616 (.ZN (n_8552), .A1 (n_8566), .A2 (n_8553));
NAND2_X1 i_8615 (.ZN (n_8551), .A1 (n_8552), .A2 (n_8568));
NAND2_X1 i_8614 (.ZN (n_8550), .A1 (n_8551), .A2 (n_8574));
NAND3_X1 i_8613 (.ZN (n_8549), .A1 (n_8575), .A2 (n_8552), .A3 (n_8568));
OAI22_X1 i_8612 (.ZN (n_8548), .A1 (n_8957), .A2 (n_8971), .B1 (n_8821), .B2 (n_8752));
NAND2_X1 i_8611 (.ZN (n_8547), .A1 (B_imm[22]), .A2 (A_imm[13]));
NAND4_X1 i_8610 (.ZN (n_8546), .A1 (B_imm[21]), .A2 (B_imm[23]), .A3 (A_imm[14]), .A4 (A_imm[12]));
NAND2_X1 i_8609 (.ZN (n_8545), .A1 (n_8546), .A2 (n_8547));
AOI22_X1 i_8608 (.ZN (n_8544), .A1 (n_8548), .A2 (n_8545), .B1 (A_imm[27]), .B2 (B_imm[9]));
INV_X1 i_8607 (.ZN (n_8543), .A (n_8544));
NAND4_X1 i_8606 (.ZN (n_8542), .A1 (n_8545), .A2 (n_8548), .A3 (B_imm[9]), .A4 (A_imm[27]));
OAI22_X1 i_8605 (.ZN (n_8541), .A1 (n_8974), .A2 (n_8751), .B1 (n_8829), .B2 (n_8893));
NAND2_X1 i_8604 (.ZN (n_8540), .A1 (B_imm[13]), .A2 (A_imm[22]));
INV_X1 i_8603 (.ZN (n_8539), .A (n_8540));
NAND4_X1 i_8602 (.ZN (n_8538), .A1 (B_imm[25]), .A2 (B_imm[15]), .A3 (A_imm[20]), .A4 (A_imm[10]));
INV_X1 i_8601 (.ZN (n_8537), .A (n_8538));
OAI21_X1 i_8600 (.ZN (n_8536), .A (n_8541), .B1 (n_8539), .B2 (n_8537));
NAND2_X1 i_8599 (.ZN (n_8535), .A1 (n_8542), .A2 (n_8536));
NAND2_X1 i_8598 (.ZN (n_8534), .A1 (n_8827), .A2 (n_8824));
NAND2_X1 i_8597 (.ZN (n_8533), .A1 (n_8534), .A2 (n_8825));
NAND3_X1 i_8596 (.ZN (n_8532), .A1 (n_8827), .A2 (n_8826), .A3 (n_8824));
NAND2_X1 i_8595 (.ZN (n_8531), .A1 (n_8533), .A2 (n_8532));
NAND3_X1 i_8594 (.ZN (n_8530), .A1 (n_8535), .A2 (n_8543), .A3 (n_8531));
INV_X1 i_8593 (.ZN (n_8529), .A (n_8530));
NAND2_X1 i_8592 (.ZN (n_8528), .A1 (n_8535), .A2 (n_8543));
NAND3_X1 i_8591 (.ZN (n_8527), .A1 (n_8528), .A2 (n_8533), .A3 (n_8532));
NAND2_X1 i_8590 (.ZN (n_8526), .A1 (B_imm[27]), .A2 (A_imm[10]));
INV_X4 i_8589 (.ZN (n_8525), .A (B_imm[19]));
OAI22_X1 i_8588 (.ZN (n_8524), .A1 (n_8525), .A2 (n_8956), .B1 (n_8993), .B2 (n_8926));
NAND4_X1 i_8587 (.ZN (n_8523), .A1 (B_imm[19]), .A2 (B_imm[26]), .A3 (A_imm[18]), .A4 (A_imm[11]));
AOI21_X1 i_8586 (.ZN (n_8522), .A (n_8526), .B1 (n_8524), .B2 (n_8523));
NAND3_X1 i_8585 (.ZN (n_8521), .A1 (n_8524), .A2 (n_8526), .A3 (n_8523));
INV_X1 i_8584 (.ZN (n_8520), .A (n_8521));
NOR2_X1 i_8583 (.ZN (n_8519), .A1 (n_8522), .A2 (n_8520));
INV_X1 i_8582 (.ZN (n_8518), .A (n_8519));
AOI21_X1 i_8581 (.ZN (n_8517), .A (n_8529), .B1 (n_8527), .B2 (n_8518));
NAND2_X2 i_8580 (.ZN (n_8516), .A1 (n_8549), .A2 (n_8517));
NAND2_X1 i_8579 (.ZN (n_8515), .A1 (n_8516), .A2 (n_8550));
NAND3_X1 i_8578 (.ZN (n_8514), .A1 (n_8515), .A2 (n_8580), .A3 (n_8579));
NAND2_X1 i_8577 (.ZN (n_8513), .A1 (n_8580), .A2 (n_8579));
NAND3_X1 i_8576 (.ZN (n_8512), .A1 (n_8516), .A2 (n_8513), .A3 (n_8550));
INV_X4 i_8575 (.ZN (n_8511), .A (A_imm[8]));
AOI22_X1 i_8574 (.ZN (n_8510), .A1 (A_imm[20]), .A2 (B_imm[16]), .B1 (B_imm[17]), .B2 (A_imm[19]));
INV_X1 i_8573 (.ZN (n_8509), .A (n_8510));
NAND2_X1 i_8572 (.ZN (n_8508), .A1 (B_imm[12]), .A2 (A_imm[24]));
NAND4_X1 i_8571 (.ZN (n_8507), .A1 (A_imm[20]), .A2 (B_imm[17]), .A3 (B_imm[16]), .A4 (A_imm[19]));
NAND2_X1 i_8570 (.ZN (n_8506), .A1 (n_8507), .A2 (n_8508));
NAND2_X1 i_8569 (.ZN (n_8505), .A1 (n_8506), .A2 (n_8509));
OAI21_X1 i_8568 (.ZN (n_8504), .A (n_8505), .B1 (n_9006), .B2 (n_8511));
NAND2_X1 i_8567 (.ZN (n_8503), .A1 (A_imm[28]), .A2 (B_imm[9]));
NAND4_X1 i_8566 (.ZN (n_8502), .A1 (n_8506), .A2 (B_imm[29]), .A3 (n_8509), .A4 (A_imm[8]));
NAND2_X1 i_8565 (.ZN (n_8501), .A1 (n_8502), .A2 (n_8503));
NAND4_X1 i_8564 (.ZN (n_8500), .A1 (n_8501), .A2 (n_8504), .A3 (B_imm[9]), .A4 (A_imm[29]));
AOI22_X1 i_8563 (.ZN (n_8499), .A1 (n_8501), .A2 (n_8504), .B1 (A_imm[29]), .B2 (B_imm[9]));
INV_X1 i_8562 (.ZN (n_8498), .A (n_8499));
NAND2_X1 i_8561 (.ZN (n_8497), .A1 (A_imm[31]), .A2 (B_imm[7]));
OAI22_X1 i_8560 (.ZN (n_8496), .A1 (n_8948), .A2 (n_8971), .B1 (n_8972), .B2 (n_8795));
NAND4_X1 i_8559 (.ZN (n_8495), .A1 (B_imm[24]), .A2 (A_imm[26]), .A3 (B_imm[12]), .A4 (A_imm[14]));
NAND2_X1 i_8558 (.ZN (n_8494), .A1 (n_8496), .A2 (n_8495));
INV_X1 i_8557 (.ZN (n_8493), .A (n_8494));
NOR2_X1 i_8556 (.ZN (n_8492), .A1 (n_8493), .A2 (n_8497));
NAND2_X1 i_8555 (.ZN (n_8491), .A1 (n_8493), .A2 (n_8497));
INV_X1 i_8554 (.ZN (n_8490), .A (n_8491));
NOR2_X1 i_8553 (.ZN (n_8489), .A1 (n_8492), .A2 (n_8490));
NAND3_X1 i_8552 (.ZN (n_8488), .A1 (n_8498), .A2 (n_8489), .A3 (n_8500));
INV_X1 i_8551 (.ZN (n_8487), .A (n_8500));
OAI22_X1 i_8550 (.ZN (n_8486), .A1 (n_8487), .A2 (n_8499), .B1 (n_8492), .B2 (n_8490));
NAND2_X1 i_8549 (.ZN (n_8485), .A1 (n_8486), .A2 (n_8488));
NAND2_X1 i_8548 (.ZN (n_8484), .A1 (B_imm[14]), .A2 (A_imm[24]));
INV_X1 i_8547 (.ZN (n_8483), .A (n_8484));
NAND2_X1 i_8546 (.ZN (n_8482), .A1 (n_8523), .A2 (n_8526));
INV_X1 i_8545 (.ZN (n_8481), .A (n_8747));
OAI21_X1 i_8544 (.ZN (n_8480), .A (n_8745), .B1 (n_8481), .B2 (n_8743));
NAND3_X1 i_8543 (.ZN (n_8479), .A1 (n_8747), .A2 (n_8746), .A3 (n_8744));
NAND2_X1 i_8542 (.ZN (n_8478), .A1 (n_8480), .A2 (n_8479));
NAND3_X1 i_8541 (.ZN (n_8477), .A1 (n_8478), .A2 (n_8524), .A3 (n_8482));
NAND2_X1 i_8540 (.ZN (n_8476), .A1 (n_8482), .A2 (n_8524));
NAND3_X1 i_8539 (.ZN (n_8475), .A1 (n_8476), .A2 (n_8480), .A3 (n_8479));
NAND2_X1 i_8538 (.ZN (n_8474), .A1 (n_8475), .A2 (n_8477));
NAND2_X1 i_8537 (.ZN (n_8473), .A1 (n_8474), .A2 (n_8483));
NAND3_X1 i_8536 (.ZN (n_8472), .A1 (n_8475), .A2 (n_8484), .A3 (n_8477));
NAND2_X1 i_8535 (.ZN (n_8471), .A1 (n_8473), .A2 (n_8472));
NAND2_X1 i_8534 (.ZN (n_8470), .A1 (n_8485), .A2 (n_8471));
NAND4_X2 i_8533 (.ZN (n_8469), .A1 (n_8488), .A2 (n_8486), .A3 (n_8473), .A4 (n_8472));
INV_X1 i_8532 (.ZN (n_8468), .A (n_8503));
NAND2_X1 i_8531 (.ZN (n_8467), .A1 (n_8504), .A2 (n_8502));
NAND2_X1 i_8530 (.ZN (n_8466), .A1 (n_8467), .A2 (n_8468));
NAND3_X1 i_8529 (.ZN (n_8465), .A1 (n_8504), .A2 (n_8502), .A3 (n_8503));
NAND2_X1 i_8528 (.ZN (n_8464), .A1 (n_8466), .A2 (n_8465));
INV_X1 i_8527 (.ZN (n_8463), .A (n_8508));
INV_X1 i_8526 (.ZN (n_8462), .A (n_8507));
OAI21_X1 i_8525 (.ZN (n_8461), .A (n_8463), .B1 (n_8462), .B2 (n_8510));
NAND3_X1 i_8524 (.ZN (n_8460), .A1 (n_8509), .A2 (n_8508), .A3 (n_8507));
NAND2_X1 i_8523 (.ZN (n_8459), .A1 (n_8460), .A2 (n_8461));
NAND3_X1 i_8522 (.ZN (n_8458), .A1 (n_8459), .A2 (B_imm[14]), .A3 (A_imm[22]));
NAND2_X1 i_8521 (.ZN (n_8457), .A1 (B_imm[14]), .A2 (A_imm[22]));
INV_X1 i_8520 (.ZN (n_8456), .A (n_8459));
NAND2_X1 i_8519 (.ZN (n_8455), .A1 (n_8457), .A2 (n_8456));
NAND2_X1 i_8518 (.ZN (n_8454), .A1 (B_imm[19]), .A2 (A_imm[16]));
NAND2_X1 i_8517 (.ZN (n_8453), .A1 (B_imm[27]), .A2 (A_imm[8]));
NAND2_X1 i_8516 (.ZN (n_8452), .A1 (n_8453), .A2 (n_8454));
NAND4_X1 i_8515 (.ZN (n_8451), .A1 (B_imm[27]), .A2 (B_imm[19]), .A3 (A_imm[16]), .A4 (A_imm[8]));
INV_X1 i_8514 (.ZN (n_8450), .A (n_8451));
OAI22_X1 i_8513 (.ZN (n_8449), .A1 (n_8956), .A2 (n_8908), .B1 (n_8955), .B2 (n_8909));
NAND2_X1 i_8512 (.ZN (n_8448), .A1 (A_imm[24]), .A2 (B_imm[10]));
INV_X1 i_8511 (.ZN (n_8447), .A (n_8448));
NAND4_X1 i_8510 (.ZN (n_8446), .A1 (A_imm[18]), .A2 (B_imm[16]), .A3 (A_imm[17]), .A4 (B_imm[17]));
INV_X1 i_8509 (.ZN (n_8445), .A (n_8446));
OAI21_X1 i_8508 (.ZN (n_8444), .A (n_8449), .B1 (n_8447), .B2 (n_8445));
INV_X1 i_8507 (.ZN (n_8443), .A (n_8444));
OAI21_X1 i_8506 (.ZN (n_8442), .A (n_8452), .B1 (n_8450), .B2 (n_8443));
INV_X1 i_8505 (.ZN (n_8441), .A (n_8442));
NAND2_X1 i_8504 (.ZN (n_8440), .A1 (n_8441), .A2 (n_8455));
NAND2_X1 i_8503 (.ZN (n_8439), .A1 (n_8440), .A2 (n_8458));
NAND2_X1 i_8502 (.ZN (n_8438), .A1 (n_8439), .A2 (n_8464));
NAND4_X1 i_8501 (.ZN (n_8437), .A1 (n_8440), .A2 (n_8466), .A3 (n_8465), .A4 (n_8458));
OAI22_X1 i_8500 (.ZN (n_8436), .A1 (n_8958), .A2 (n_8971), .B1 (n_8957), .B2 (n_8946));
NAND2_X1 i_8499 (.ZN (n_8435), .A1 (B_imm[15]), .A2 (A_imm[21]));
INV_X1 i_8498 (.ZN (n_8434), .A (n_8435));
NAND4_X1 i_8497 (.ZN (n_8433), .A1 (B_imm[22]), .A2 (B_imm[21]), .A3 (A_imm[15]), .A4 (A_imm[14]));
INV_X1 i_8496 (.ZN (n_8432), .A (n_8433));
OAI21_X1 i_8495 (.ZN (n_8431), .A (n_8436), .B1 (n_8434), .B2 (n_8432));
INV_X1 i_8494 (.ZN (n_8430), .A (n_8431));
INV_X4 i_8493 (.ZN (n_8429), .A (B_imm[5]));
OAI22_X1 i_8492 (.ZN (n_8428), .A1 (n_8948), .A2 (n_8752), .B1 (n_9037), .B2 (n_8429));
NAND2_X1 i_8491 (.ZN (n_8427), .A1 (B_imm[23]), .A2 (A_imm[13]));
NAND4_X1 i_8490 (.ZN (n_8426), .A1 (B_imm[24]), .A2 (A_imm[31]), .A3 (B_imm[5]), .A4 (A_imm[12]));
NAND2_X1 i_8489 (.ZN (n_8425), .A1 (n_8426), .A2 (n_8427));
NAND2_X1 i_8488 (.ZN (n_8424), .A1 (n_8425), .A2 (n_8428));
INV_X4 i_8487 (.ZN (n_8423), .A (B_imm[18]));
NAND2_X1 i_8486 (.ZN (n_8422), .A1 (A_imm[26]), .A2 (B_imm[10]));
OAI21_X1 i_8485 (.ZN (n_8421), .A (n_8422), .B1 (n_8423), .B2 (n_8956));
NAND2_X1 i_8484 (.ZN (n_8420), .A1 (A_imm[25]), .A2 (B_imm[11]));
NAND4_X1 i_8483 (.ZN (n_8419), .A1 (B_imm[18]), .A2 (A_imm[26]), .A3 (B_imm[10]), .A4 (A_imm[18]));
NAND2_X1 i_8482 (.ZN (n_8418), .A1 (n_8419), .A2 (n_8420));
NAND2_X1 i_8481 (.ZN (n_8417), .A1 (n_8418), .A2 (n_8421));
NAND2_X1 i_8480 (.ZN (n_8416), .A1 (n_8424), .A2 (n_8417));
NAND4_X1 i_8479 (.ZN (n_8415), .A1 (n_8425), .A2 (n_8428), .A3 (n_8418), .A4 (n_8421));
NAND2_X1 i_8478 (.ZN (n_8414), .A1 (n_8415), .A2 (n_8416));
NAND2_X1 i_8477 (.ZN (n_8413), .A1 (n_8414), .A2 (n_8430));
NAND3_X1 i_8476 (.ZN (n_8412), .A1 (n_8416), .A2 (n_8415), .A3 (n_8431));
NAND2_X1 i_8475 (.ZN (n_8411), .A1 (n_8413), .A2 (n_8412));
NAND2_X1 i_8474 (.ZN (n_8410), .A1 (n_8437), .A2 (n_8411));
NAND2_X1 i_8473 (.ZN (n_8409), .A1 (n_8410), .A2 (n_8438));
NAND2_X1 i_8472 (.ZN (n_8408), .A1 (n_8469), .A2 (n_8409));
NAND2_X2 i_8471 (.ZN (n_8407), .A1 (n_8408), .A2 (n_8470));
INV_X1 i_8470 (.ZN (n_8406), .A (n_8407));
NAND2_X1 i_8469 (.ZN (n_8405), .A1 (n_8512), .A2 (n_8406));
NAND4_X2 i_8468 (.ZN (n_8404), .A1 (n_8405), .A2 (n_8514), .A3 (n_8582), .A4 (n_8587));
NAND2_X1 i_8467 (.ZN (n_8403), .A1 (n_8582), .A2 (n_8587));
NAND2_X1 i_8466 (.ZN (n_8402), .A1 (n_8405), .A2 (n_8514));
INV_X1 i_8465 (.ZN (n_8401), .A (n_8749));
INV_X1 i_8464 (.ZN (n_8400), .A (n_8742));
OAI21_X1 i_8463 (.ZN (n_8399), .A (n_8750), .B1 (n_8400), .B2 (n_8401));
INV_X1 i_8462 (.ZN (n_8398), .A (n_8399));
NAND2_X1 i_8461 (.ZN (n_8397), .A1 (B_imm[18]), .A2 (A_imm[22]));
OAI22_X1 i_8460 (.ZN (n_8396), .A1 (n_8909), .A2 (n_8907), .B1 (n_8767), .B2 (n_8908));
NAND4_X1 i_8459 (.ZN (n_8395), .A1 (A_imm[23]), .A2 (A_imm[24]), .A3 (B_imm[17]), .A4 (B_imm[16]));
AOI21_X1 i_8458 (.ZN (n_8394), .A (n_8397), .B1 (n_8396), .B2 (n_8395));
NAND3_X1 i_8457 (.ZN (n_8393), .A1 (n_8396), .A2 (n_8397), .A3 (n_8395));
INV_X1 i_8456 (.ZN (n_8392), .A (n_8393));
OAI21_X1 i_8455 (.ZN (n_8391), .A (n_8398), .B1 (n_8394), .B2 (n_8392));
INV_X1 i_8454 (.ZN (n_8390), .A (n_8394));
NAND3_X1 i_8453 (.ZN (n_8389), .A1 (n_8399), .A2 (n_8390), .A3 (n_8393));
NAND2_X1 i_8452 (.ZN (n_8388), .A1 (B_imm[15]), .A2 (A_imm[25]));
OAI22_X1 i_8451 (.ZN (n_8387), .A1 (n_8958), .A2 (n_8956), .B1 (n_8957), .B2 (n_8892));
NAND4_X1 i_8450 (.ZN (n_8386), .A1 (B_imm[22]), .A2 (B_imm[21]), .A3 (A_imm[19]), .A4 (A_imm[18]));
AOI21_X1 i_8449 (.ZN (n_8385), .A (n_8388), .B1 (n_8387), .B2 (n_8386));
NAND3_X1 i_8448 (.ZN (n_8384), .A1 (n_8387), .A2 (n_8388), .A3 (n_8386));
INV_X1 i_8447 (.ZN (n_8383), .A (n_8384));
NOR2_X1 i_8446 (.ZN (n_8382), .A1 (n_8385), .A2 (n_8383));
NAND3_X1 i_8445 (.ZN (n_8381), .A1 (n_8391), .A2 (n_8389), .A3 (n_8382));
INV_X1 i_8444 (.ZN (n_8380), .A (n_8381));
AOI21_X1 i_8443 (.ZN (n_8379), .A (n_8382), .B1 (n_8391), .B2 (n_8389));
NOR2_X1 i_8442 (.ZN (n_8378), .A1 (n_8380), .A2 (n_8379));
OAI22_X1 i_8441 (.ZN (n_8377), .A1 (n_8957), .A2 (n_8955), .B1 (n_8821), .B2 (n_8946));
NAND2_X1 i_8440 (.ZN (n_8376), .A1 (B_imm[22]), .A2 (A_imm[16]));
INV_X1 i_8439 (.ZN (n_8375), .A (n_8376));
NAND4_X1 i_8438 (.ZN (n_8374), .A1 (B_imm[21]), .A2 (B_imm[23]), .A3 (A_imm[17]), .A4 (A_imm[15]));
INV_X1 i_8437 (.ZN (n_8373), .A (n_8374));
OAI21_X1 i_8436 (.ZN (n_8372), .A (n_8377), .B1 (n_8375), .B2 (n_8373));
INV_X1 i_8435 (.ZN (n_8371), .A (n_8372));
NAND2_X1 i_8434 (.ZN (n_8370), .A1 (n_8495), .A2 (n_8497));
NAND2_X1 i_8433 (.ZN (n_8369), .A1 (n_8496), .A2 (n_8370));
OAI21_X1 i_8432 (.ZN (n_8368), .A (n_8369), .B1 (n_8849), .B2 (n_9020));
INV_X1 i_8431 (.ZN (n_8367), .A (n_8368));
INV_X1 i_8430 (.ZN (n_8366), .A (n_8369));
NAND3_X1 i_8429 (.ZN (n_8365), .A1 (n_8366), .A2 (B_imm[11]), .A3 (A_imm[28]));
INV_X1 i_8428 (.ZN (n_8364), .A (n_8365));
OAI21_X1 i_8427 (.ZN (n_8363), .A (n_8371), .B1 (n_8367), .B2 (n_8364));
NAND3_X1 i_8426 (.ZN (n_8362), .A1 (n_8365), .A2 (n_8372), .A3 (n_8368));
NAND2_X1 i_8425 (.ZN (n_8361), .A1 (n_8363), .A2 (n_8362));
NAND2_X1 i_8424 (.ZN (n_8360), .A1 (n_8475), .A2 (n_8483));
NAND2_X1 i_8423 (.ZN (n_8359), .A1 (n_8360), .A2 (n_8477));
NAND2_X1 i_8422 (.ZN (n_8358), .A1 (n_8361), .A2 (n_8359));
NAND4_X2 i_8421 (.ZN (n_8357), .A1 (n_8363), .A2 (n_8477), .A3 (n_8362), .A4 (n_8360));
OAI21_X1 i_8420 (.ZN (n_8356), .A (n_8500), .B1 (n_8489), .B2 (n_8499));
NAND2_X2 i_8419 (.ZN (n_8355), .A1 (n_8357), .A2 (n_8356));
AOI21_X1 i_8418 (.ZN (n_8354), .A (n_8378), .B1 (n_8358), .B2 (n_8355));
NAND3_X2 i_8417 (.ZN (n_8353), .A1 (n_8355), .A2 (n_8378), .A3 (n_8358));
INV_X1 i_8416 (.ZN (n_8352), .A (n_8353));
NAND2_X1 i_8415 (.ZN (n_8351), .A1 (n_8365), .A2 (n_8372));
NAND2_X1 i_8414 (.ZN (n_8350), .A1 (n_8351), .A2 (n_8368));
NAND2_X1 i_8413 (.ZN (n_8349), .A1 (B_imm[23]), .A2 (A_imm[17]));
INV_X1 i_8412 (.ZN (n_8348), .A (n_8349));
INV_X2 i_8411 (.ZN (n_8347), .A (B_imm[9]));
OAI22_X1 i_8410 (.ZN (n_8346), .A1 (n_8347), .A2 (n_9037), .B1 (n_8948), .B2 (n_8858));
INV_X1 i_8409 (.ZN (n_8345), .A (n_8346));
NAND4_X1 i_8408 (.ZN (n_8344), .A1 (B_imm[24]), .A2 (opt_ipoPP_0), .A3 (B_imm[9]), .A4 (A_imm[16]));
INV_X1 i_8407 (.ZN (n_8343), .A (n_8344));
OAI21_X1 i_8406 (.ZN (n_8342), .A (n_8348), .B1 (n_8345), .B2 (n_8343));
NAND3_X1 i_8405 (.ZN (n_8341), .A1 (n_8346), .A2 (n_8349), .A3 (n_8344));
NAND3_X1 i_8404 (.ZN (n_8340), .A1 (n_8350), .A2 (n_8342), .A3 (n_8341));
NAND2_X1 i_8403 (.ZN (n_8339), .A1 (n_8342), .A2 (n_8341));
NAND3_X1 i_8402 (.ZN (n_8338), .A1 (n_8351), .A2 (n_8368), .A3 (n_8339));
NAND2_X1 i_8401 (.ZN (n_8337), .A1 (B_imm[27]), .A2 (A_imm[13]));
INV_X1 i_8400 (.ZN (n_8336), .A (n_8337));
OAI22_X1 i_8399 (.ZN (n_8335), .A1 (n_8525), .A2 (n_8859), .B1 (n_8993), .B2 (n_8971));
NAND4_X1 i_8398 (.ZN (n_8334), .A1 (B_imm[19]), .A2 (B_imm[26]), .A3 (A_imm[21]), .A4 (A_imm[14]));
NAND2_X1 i_8397 (.ZN (n_8333), .A1 (n_8335), .A2 (n_8334));
XNOR2_X1 i_8396 (.ZN (n_8332), .A (n_8333), .B (n_8336));
AOI21_X1 i_8395 (.ZN (n_8331), .A (n_8332), .B1 (n_8340), .B2 (n_8338));
NAND3_X1 i_8394 (.ZN (n_8330), .A1 (n_8340), .A2 (n_8338), .A3 (n_8332));
INV_X1 i_8393 (.ZN (n_8329), .A (n_8330));
NOR2_X1 i_8392 (.ZN (n_8328), .A1 (n_8329), .A2 (n_8331));
OAI21_X1 i_8391 (.ZN (n_8327), .A (n_8328), .B1 (n_8354), .B2 (n_8352));
INV_X2 i_8390 (.ZN (n_8326), .A (n_8354));
INV_X1 i_8389 (.ZN (n_8325), .A (n_8328));
NAND3_X1 i_8388 (.ZN (n_8324), .A1 (n_8326), .A2 (n_8353), .A3 (n_8325));
AOI22_X1 i_8387 (.ZN (n_8323), .A1 (n_8402), .A2 (n_8403), .B1 (n_8327), .B2 (n_8324));
INV_X1 i_8386 (.ZN (n_8322), .A (n_8323));
NAND2_X1 i_8385 (.ZN (n_8321), .A1 (n_8322), .A2 (n_8404));
INV_X1 i_8384 (.ZN (n_8320), .A (n_8321));
NAND2_X1 i_8383 (.ZN (n_8319), .A1 (n_8655), .A2 (n_8320));
NAND3_X1 i_8382 (.ZN (n_8318), .A1 (n_8321), .A2 (n_8658), .A3 (n_8656));
NAND2_X1 i_8381 (.ZN (n_8317), .A1 (n_8319), .A2 (n_8318));
NAND2_X1 i_8380 (.ZN (n_8316), .A1 (n_8402), .A2 (n_8403));
NAND2_X1 i_8379 (.ZN (n_8315), .A1 (n_8324), .A2 (n_8327));
AOI21_X1 i_8378 (.ZN (n_8314), .A (n_8315), .B1 (n_8316), .B2 (n_8404));
INV_X1 i_8377 (.ZN (n_8313), .A (n_8314));
NAND3_X1 i_8376 (.ZN (n_8312), .A1 (n_8316), .A2 (n_8404), .A3 (n_8315));
NAND2_X1 i_8375 (.ZN (n_8311), .A1 (n_8702), .A2 (n_8706));
NAND3_X1 i_8374 (.ZN (n_8310), .A1 (n_8716), .A2 (n_8311), .A3 (n_8715));
INV_X1 i_8373 (.ZN (n_8309), .A (n_8311));
NAND2_X1 i_8372 (.ZN (n_8308), .A1 (n_8716), .A2 (n_8715));
NAND2_X1 i_8371 (.ZN (n_8307), .A1 (n_8308), .A2 (n_8309));
NAND2_X1 i_8370 (.ZN (n_8306), .A1 (n_8307), .A2 (n_8310));
INV_X1 i_8369 (.ZN (n_8305), .A (n_8306));
INV_X1 i_8368 (.ZN (n_8304), .A (n_8682));
NAND2_X1 i_8367 (.ZN (n_8303), .A1 (n_8683), .A2 (n_8681));
NAND2_X1 i_8366 (.ZN (n_8302), .A1 (n_8303), .A2 (n_8304));
NAND3_X1 i_8365 (.ZN (n_8301), .A1 (n_8683), .A2 (n_8682), .A3 (n_8681));
NAND2_X1 i_8364 (.ZN (n_8300), .A1 (n_8302), .A2 (n_8301));
NAND2_X1 i_8363 (.ZN (n_8299), .A1 (n_8712), .A2 (n_8709));
NAND2_X1 i_8362 (.ZN (n_8298), .A1 (n_8299), .A2 (n_8710));
NAND3_X1 i_8361 (.ZN (n_8297), .A1 (n_8712), .A2 (n_8711), .A3 (n_8709));
NAND2_X1 i_8360 (.ZN (n_8296), .A1 (n_8298), .A2 (n_8297));
NAND2_X1 i_8359 (.ZN (n_8295), .A1 (n_8300), .A2 (n_8296));
NAND4_X1 i_8358 (.ZN (n_8294), .A1 (n_8302), .A2 (n_8298), .A3 (n_8301), .A4 (n_8297));
INV_X4 i_8357 (.ZN (n_8293), .A (A_imm[5]));
NAND2_X1 i_8356 (.ZN (n_8292), .A1 (A_imm[27]), .A2 (B_imm[8]));
OAI21_X1 i_8355 (.ZN (n_8291), .A (n_8292), .B1 (n_9004), .B2 (n_8293));
OAI22_X1 i_8354 (.ZN (n_8290), .A1 (n_8860), .A2 (n_8971), .B1 (n_8973), .B2 (n_8859));
NAND2_X1 i_8353 (.ZN (n_8289), .A1 (B_imm[28]), .A2 (A_imm[6]));
INV_X1 i_8352 (.ZN (n_8288), .A (n_8289));
NAND4_X1 i_8351 (.ZN (n_8287), .A1 (B_imm[20]), .A2 (B_imm[13]), .A3 (A_imm[21]), .A4 (A_imm[14]));
INV_X1 i_8350 (.ZN (n_8286), .A (n_8287));
OAI21_X1 i_8349 (.ZN (n_8285), .A (n_8290), .B1 (n_8288), .B2 (n_8286));
NAND4_X1 i_8348 (.ZN (n_8284), .A1 (B_imm[30]), .A2 (A_imm[27]), .A3 (B_imm[8]), .A4 (A_imm[5]));
NAND2_X1 i_8347 (.ZN (n_8283), .A1 (n_8285), .A2 (n_8284));
NAND2_X1 i_8346 (.ZN (n_8282), .A1 (n_8283), .A2 (n_8291));
INV_X1 i_8345 (.ZN (n_8281), .A (n_8282));
NAND2_X1 i_8344 (.ZN (n_8280), .A1 (n_8281), .A2 (n_8294));
NAND2_X1 i_8343 (.ZN (n_8279), .A1 (n_8280), .A2 (n_8295));
INV_X1 i_8342 (.ZN (n_8278), .A (n_8676));
NAND2_X1 i_8341 (.ZN (n_8277), .A1 (n_8678), .A2 (n_8677));
NAND2_X1 i_8340 (.ZN (n_8276), .A1 (n_8277), .A2 (n_8278));
NAND3_X1 i_8339 (.ZN (n_8275), .A1 (n_8678), .A2 (n_8677), .A3 (n_8676));
NAND2_X1 i_8338 (.ZN (n_8274), .A1 (n_8276), .A2 (n_8275));
NAND2_X1 i_8337 (.ZN (n_8273), .A1 (n_8279), .A2 (n_8274));
NAND4_X1 i_8336 (.ZN (n_8272), .A1 (n_8280), .A2 (n_8276), .A3 (n_8295), .A4 (n_8275));
AOI21_X1 i_8335 (.ZN (n_8271), .A (n_8635), .B1 (n_8643), .B2 (n_8633));
NAND3_X1 i_8334 (.ZN (n_8270), .A1 (n_8643), .A2 (n_8635), .A3 (n_8633));
INV_X1 i_8333 (.ZN (n_8269), .A (n_8270));
OAI211_X1 i_8332 (.ZN (n_8268), .A (B_imm[6]), .B (A_imm[30]), .C1 (n_8269), .C2 (n_8271));
NAND2_X1 i_8331 (.ZN (n_8267), .A1 (A_imm[30]), .A2 (B_imm[6]));
NOR2_X1 i_8330 (.ZN (n_8266), .A1 (n_8269), .A2 (n_8271));
NAND2_X1 i_8329 (.ZN (n_8265), .A1 (n_8266), .A2 (n_8267));
NAND2_X1 i_8328 (.ZN (n_8264), .A1 (n_8640), .A2 (n_8637));
NAND2_X1 i_8327 (.ZN (n_8263), .A1 (n_8264), .A2 (n_8638));
NAND3_X1 i_8326 (.ZN (n_8262), .A1 (n_8639), .A2 (n_8640), .A3 (n_8637));
NAND2_X1 i_8325 (.ZN (n_8261), .A1 (n_8263), .A2 (n_8262));
NAND3_X1 i_8324 (.ZN (n_8260), .A1 (n_8261), .A2 (B_imm[31]), .A3 (A_imm[4]));
NAND2_X1 i_8323 (.ZN (n_8259), .A1 (B_imm[31]), .A2 (A_imm[4]));
INV_X1 i_8322 (.ZN (n_8258), .A (n_8261));
NAND2_X1 i_8321 (.ZN (n_8257), .A1 (n_8258), .A2 (n_8259));
INV_X1 i_8320 (.ZN (n_8256), .A (n_8257));
OAI22_X1 i_8319 (.ZN (n_8255), .A1 (n_8525), .A2 (n_8946), .B1 (n_8993), .B2 (n_8511));
NAND2_X1 i_8318 (.ZN (n_8254), .A1 (B_imm[27]), .A2 (A_imm[7]));
INV_X1 i_8317 (.ZN (n_8253), .A (n_8254));
NAND4_X1 i_8316 (.ZN (n_8252), .A1 (B_imm[19]), .A2 (B_imm[26]), .A3 (A_imm[15]), .A4 (A_imm[8]));
INV_X1 i_8315 (.ZN (n_8251), .A (n_8252));
OAI21_X1 i_8314 (.ZN (n_8250), .A (n_8255), .B1 (n_8253), .B2 (n_8251));
OAI21_X1 i_8313 (.ZN (n_8249), .A (n_8260), .B1 (n_8256), .B2 (n_8250));
NAND2_X1 i_8312 (.ZN (n_8248), .A1 (n_8265), .A2 (n_8249));
NAND2_X1 i_8311 (.ZN (n_8247), .A1 (n_8248), .A2 (n_8268));
NAND2_X1 i_8310 (.ZN (n_8246), .A1 (n_8247), .A2 (n_8272));
NAND3_X1 i_8309 (.ZN (n_8245), .A1 (n_8246), .A2 (n_8305), .A3 (n_8273));
NAND2_X1 i_8308 (.ZN (n_8244), .A1 (n_8246), .A2 (n_8273));
NAND2_X1 i_8307 (.ZN (n_8243), .A1 (n_8244), .A2 (n_8306));
NAND3_X1 i_8306 (.ZN (n_8242), .A1 (n_8648), .A2 (n_8646), .A3 (n_8631));
INV_X1 i_8305 (.ZN (n_8241), .A (n_8631));
NAND2_X1 i_8304 (.ZN (n_8240), .A1 (n_8648), .A2 (n_8646));
NAND2_X1 i_8303 (.ZN (n_8239), .A1 (n_8240), .A2 (n_8241));
NAND3_X1 i_8302 (.ZN (n_8238), .A1 (n_8616), .A2 (n_8598), .A3 (n_8615));
NAND2_X1 i_8301 (.ZN (n_8237), .A1 (n_8616), .A2 (n_8615));
NAND2_X1 i_8300 (.ZN (n_8236), .A1 (n_8237), .A2 (n_8597));
AOI22_X1 i_8299 (.ZN (n_8235), .A1 (n_8236), .A2 (n_8238), .B1 (n_8239), .B2 (n_8242));
NAND4_X1 i_8298 (.ZN (n_8234), .A1 (n_8236), .A2 (n_8239), .A3 (n_8242), .A4 (n_8238));
NAND4_X1 i_8297 (.ZN (n_8233), .A1 (A_imm[29]), .A2 (B_imm[14]), .A3 (B_imm[6]), .A4 (A_imm[21]));
INV_X2 i_8296 (.ZN (n_8232), .A (B_imm[6]));
NAND2_X1 i_8295 (.ZN (n_8231), .A1 (B_imm[14]), .A2 (A_imm[21]));
OAI21_X1 i_8294 (.ZN (n_8230), .A (n_8231), .B1 (n_8994), .B2 (n_8232));
AOI21_X1 i_8293 (.ZN (n_8229), .A (n_8612), .B1 (n_8613), .B2 (n_8611));
NAND3_X1 i_8292 (.ZN (n_8228), .A1 (n_8613), .A2 (n_8612), .A3 (n_8611));
INV_X1 i_8291 (.ZN (n_8227), .A (n_8228));
NOR2_X1 i_8290 (.ZN (n_8226), .A1 (n_8227), .A2 (n_8229));
INV_X1 i_8289 (.ZN (n_8225), .A (n_8226));
NAND2_X1 i_8288 (.ZN (n_8224), .A1 (n_8230), .A2 (n_8225));
NAND2_X1 i_8287 (.ZN (n_8223), .A1 (n_8224), .A2 (n_8233));
INV_X1 i_8286 (.ZN (n_8222), .A (n_8607));
INV_X1 i_8285 (.ZN (n_8221), .A (n_8600));
OAI21_X1 i_8284 (.ZN (n_8220), .A (n_8221), .B1 (n_8222), .B2 (n_8609));
NAND3_X1 i_8283 (.ZN (n_8219), .A1 (n_8608), .A2 (n_8607), .A3 (n_8600));
NAND2_X1 i_8282 (.ZN (n_8218), .A1 (n_8219), .A2 (n_8220));
NAND2_X1 i_8281 (.ZN (n_8217), .A1 (n_8223), .A2 (n_8218));
NAND4_X1 i_8280 (.ZN (n_8216), .A1 (n_8224), .A2 (n_8219), .A3 (n_8220), .A4 (n_8233));
INV_X1 i_8279 (.ZN (n_8215), .A (n_8542));
INV_X1 i_8278 (.ZN (n_8214), .A (n_8536));
OAI21_X1 i_8277 (.ZN (n_8213), .A (n_8214), .B1 (n_8215), .B2 (n_8544));
NAND3_X1 i_8276 (.ZN (n_8212), .A1 (n_8543), .A2 (n_8542), .A3 (n_8536));
NAND2_X1 i_8275 (.ZN (n_8211), .A1 (n_8212), .A2 (n_8213));
NAND2_X1 i_8274 (.ZN (n_8210), .A1 (n_8216), .A2 (n_8211));
NAND2_X1 i_8273 (.ZN (n_8209), .A1 (n_8210), .A2 (n_8217));
AOI21_X1 i_8272 (.ZN (n_8208), .A (n_8235), .B1 (n_8209), .B2 (n_8234));
NAND2_X1 i_8271 (.ZN (n_8207), .A1 (n_8243), .A2 (n_8208));
AOI21_X1 i_8270 (.ZN (n_8206), .A (n_8668), .B1 (n_8687), .B2 (n_8686));
NAND3_X1 i_8269 (.ZN (n_8205), .A1 (n_8687), .A2 (n_8686), .A3 (n_8668));
INV_X1 i_8268 (.ZN (n_8204), .A (n_8205));
NOR2_X1 i_8267 (.ZN (n_8203), .A1 (n_8204), .A2 (n_8206));
NAND3_X1 i_8266 (.ZN (n_8202), .A1 (n_8207), .A2 (n_8203), .A3 (n_8245));
AOI22_X1 i_8265 (.ZN (n_8201), .A1 (n_8246), .A2 (n_8273), .B1 (n_8310), .B2 (n_8307));
NAND2_X1 i_8264 (.ZN (n_8200), .A1 (n_8239), .A2 (n_8242));
NAND2_X1 i_8263 (.ZN (n_8199), .A1 (n_8236), .A2 (n_8238));
NAND2_X1 i_8262 (.ZN (n_8198), .A1 (n_8199), .A2 (n_8200));
INV_X1 i_8261 (.ZN (n_8197), .A (n_8234));
INV_X1 i_8260 (.ZN (n_8196), .A (n_8209));
OAI21_X1 i_8259 (.ZN (n_8195), .A (n_8198), .B1 (n_8196), .B2 (n_8197));
OAI21_X1 i_8258 (.ZN (n_8194), .A (n_8245), .B1 (n_8201), .B2 (n_8195));
INV_X1 i_8257 (.ZN (n_8193), .A (n_8203));
NAND2_X2 i_8256 (.ZN (n_8192), .A1 (n_8194), .A2 (n_8193));
NAND3_X1 i_8255 (.ZN (n_8191), .A1 (n_8587), .A2 (n_8586), .A3 (n_8583));
NAND2_X1 i_8254 (.ZN (n_8190), .A1 (n_8587), .A2 (n_8586));
NAND2_X1 i_8253 (.ZN (n_8189), .A1 (n_8190), .A2 (n_8584));
NAND2_X1 i_8252 (.ZN (n_8188), .A1 (n_8189), .A2 (n_8191));
NAND2_X1 i_8251 (.ZN (n_8187), .A1 (n_8192), .A2 (n_8188));
NAND2_X1 i_8250 (.ZN (n_8186), .A1 (n_8187), .A2 (n_8202));
NAND3_X2 i_8249 (.ZN (n_8185), .A1 (n_8313), .A2 (n_8312), .A3 (n_8186));
INV_X1 i_8248 (.ZN (n_8184), .A (n_8312));
INV_X1 i_8247 (.ZN (n_8183), .A (n_8186));
OAI21_X2 i_8246 (.ZN (n_8182), .A (n_8183), .B1 (n_8184), .B2 (n_8314));
NAND3_X1 i_8245 (.ZN (n_8181), .A1 (n_8514), .A2 (n_8512), .A3 (n_8407));
AOI21_X1 i_8244 (.ZN (n_8180), .A (n_8513), .B1 (n_8516), .B2 (n_8550));
INV_X1 i_8243 (.ZN (n_8179), .A (n_8512));
OAI21_X1 i_8242 (.ZN (n_8178), .A (n_8406), .B1 (n_8180), .B2 (n_8179));
NAND3_X1 i_8241 (.ZN (n_8177), .A1 (n_8550), .A2 (n_8549), .A3 (n_8517));
INV_X1 i_8240 (.ZN (n_8176), .A (n_8177));
AOI21_X1 i_8239 (.ZN (n_8175), .A (n_8517), .B1 (n_8550), .B2 (n_8549));
NAND3_X1 i_8238 (.ZN (n_8174), .A1 (n_8625), .A2 (n_8628), .A3 (n_8594));
NAND2_X1 i_8237 (.ZN (n_8173), .A1 (n_8625), .A2 (n_8628));
NAND2_X1 i_8236 (.ZN (n_8172), .A1 (n_8173), .A2 (n_8595));
NAND2_X1 i_8235 (.ZN (n_8171), .A1 (n_8172), .A2 (n_8174));
OAI21_X1 i_8234 (.ZN (n_8170), .A (n_8171), .B1 (n_8176), .B2 (n_8175));
INV_X1 i_8233 (.ZN (n_8169), .A (n_8175));
NAND4_X1 i_8232 (.ZN (n_8168), .A1 (n_8169), .A2 (n_8177), .A3 (n_8174), .A4 (n_8172));
AOI21_X1 i_8231 (.ZN (n_8167), .A (n_8531), .B1 (n_8543), .B2 (n_8535));
OAI21_X1 i_8230 (.ZN (n_8166), .A (n_8519), .B1 (n_8167), .B2 (n_8529));
NAND3_X1 i_8229 (.ZN (n_8165), .A1 (n_8527), .A2 (n_8530), .A3 (n_8518));
NAND2_X1 i_8228 (.ZN (n_8164), .A1 (n_8165), .A2 (n_8166));
INV_X1 i_8227 (.ZN (n_8163), .A (n_8164));
OAI21_X1 i_8226 (.ZN (n_8162), .A (n_8554), .B1 (n_8556), .B2 (n_8559));
NAND3_X1 i_8225 (.ZN (n_8161), .A1 (n_8558), .A2 (n_8557), .A3 (n_8555));
NAND2_X1 i_8224 (.ZN (n_8160), .A1 (n_8162), .A2 (n_8161));
OAI22_X1 i_8223 (.ZN (n_8159), .A1 (n_8858), .A2 (n_8909), .B1 (n_8908), .B2 (n_8955));
NAND2_X1 i_8222 (.ZN (n_8158), .A1 (A_imm[23]), .A2 (B_imm[10]));
NAND4_X1 i_8221 (.ZN (n_8157), .A1 (A_imm[16]), .A2 (B_imm[17]), .A3 (B_imm[16]), .A4 (A_imm[17]));
NAND2_X1 i_8220 (.ZN (n_8156), .A1 (n_8157), .A2 (n_8158));
NAND2_X1 i_8219 (.ZN (n_8155), .A1 (n_8156), .A2 (n_8159));
OAI21_X1 i_8218 (.ZN (n_8154), .A (n_8155), .B1 (n_9006), .B2 (n_8293));
NAND4_X1 i_8217 (.ZN (n_8153), .A1 (n_8156), .A2 (B_imm[29]), .A3 (n_8159), .A4 (A_imm[5]));
NAND2_X1 i_8216 (.ZN (n_8152), .A1 (B_imm[12]), .A2 (A_imm[21]));
OAI21_X1 i_8215 (.ZN (n_8151), .A (n_8152), .B1 (n_8849), .B2 (n_8906));
NAND2_X1 i_8214 (.ZN (n_8150), .A1 (A_imm[26]), .A2 (B_imm[7]));
INV_X1 i_8213 (.ZN (n_8149), .A (n_8150));
NAND4_X1 i_8212 (.ZN (n_8148), .A1 (B_imm[11]), .A2 (B_imm[12]), .A3 (A_imm[22]), .A4 (A_imm[21]));
INV_X1 i_8211 (.ZN (n_8147), .A (n_8148));
OAI21_X1 i_8210 (.ZN (n_8146), .A (n_8151), .B1 (n_8147), .B2 (n_8149));
NAND2_X1 i_8209 (.ZN (n_8145), .A1 (n_8153), .A2 (n_8146));
AOI21_X1 i_8208 (.ZN (n_8144), .A (n_8604), .B1 (n_8605), .B2 (n_8602));
NAND3_X1 i_8207 (.ZN (n_8143), .A1 (n_8605), .A2 (n_8604), .A3 (n_8602));
INV_X1 i_8206 (.ZN (n_8142), .A (n_8143));
OAI211_X1 i_8205 (.ZN (n_8141), .A (n_8145), .B (n_8154), .C1 (n_8142), .C2 (n_8144));
NAND2_X1 i_8204 (.ZN (n_8140), .A1 (n_8145), .A2 (n_8154));
NOR2_X1 i_8203 (.ZN (n_8139), .A1 (n_8142), .A2 (n_8144));
NAND2_X1 i_8202 (.ZN (n_8138), .A1 (n_8140), .A2 (n_8139));
INV_X1 i_8201 (.ZN (n_8137), .A (n_8547));
NAND2_X1 i_8200 (.ZN (n_8136), .A1 (n_8548), .A2 (n_8546));
NAND2_X1 i_8199 (.ZN (n_8135), .A1 (n_8136), .A2 (n_8137));
NAND3_X1 i_8198 (.ZN (n_8134), .A1 (n_8548), .A2 (n_8547), .A3 (n_8546));
NAND2_X1 i_8197 (.ZN (n_8133), .A1 (n_8135), .A2 (n_8134));
NAND2_X1 i_8196 (.ZN (n_8132), .A1 (n_8138), .A2 (n_8133));
NAND2_X1 i_8195 (.ZN (n_8131), .A1 (n_8132), .A2 (n_8141));
NAND2_X1 i_8194 (.ZN (n_8130), .A1 (n_8131), .A2 (n_8160));
NAND4_X1 i_8193 (.ZN (n_8129), .A1 (n_8132), .A2 (n_8162), .A3 (n_8161), .A4 (n_8141));
NAND2_X1 i_8192 (.ZN (n_8128), .A1 (A_imm[28]), .A2 (B_imm[6]));
NAND2_X1 i_8191 (.ZN (n_8127), .A1 (A_imm[25]), .A2 (B_imm[8]));
OAI21_X1 i_8190 (.ZN (n_8126), .A (n_8127), .B1 (n_8423), .B2 (n_8946));
NAND2_X1 i_8189 (.ZN (n_8125), .A1 (B_imm[9]), .A2 (A_imm[24]));
INV_X1 i_8188 (.ZN (n_8124), .A (n_8125));
NAND4_X1 i_8187 (.ZN (n_8123), .A1 (B_imm[18]), .A2 (A_imm[25]), .A3 (B_imm[8]), .A4 (A_imm[15]));
INV_X1 i_8186 (.ZN (n_8122), .A (n_8123));
OAI21_X1 i_8185 (.ZN (n_8121), .A (n_8126), .B1 (n_8122), .B2 (n_8124));
NAND2_X1 i_8184 (.ZN (n_8120), .A1 (n_8121), .A2 (n_8128));
NAND2_X1 i_8183 (.ZN (n_8119), .A1 (n_8123), .A2 (n_8125));
NAND4_X1 i_8182 (.ZN (n_8118), .A1 (n_8119), .A2 (B_imm[6]), .A3 (A_imm[28]), .A4 (n_8126));
NAND2_X1 i_8181 (.ZN (n_8117), .A1 (A_imm[31]), .A2 (B_imm[2]));
OAI21_X1 i_8180 (.ZN (n_8116), .A (n_8117), .B1 (n_8948), .B2 (n_8645));
NAND2_X1 i_8179 (.ZN (n_8115), .A1 (B_imm[23]), .A2 (A_imm[10]));
INV_X1 i_8178 (.ZN (n_8114), .A (n_8115));
NAND4_X1 i_8177 (.ZN (n_8113), .A1 (B_imm[24]), .A2 (A_imm[31]), .A3 (B_imm[2]), .A4 (A_imm[9]));
INV_X1 i_8176 (.ZN (n_8112), .A (n_8113));
OAI21_X1 i_8175 (.ZN (n_8111), .A (n_8116), .B1 (n_8112), .B2 (n_8114));
NAND2_X1 i_8174 (.ZN (n_8110), .A1 (n_8118), .A2 (n_8111));
AOI21_X1 i_8173 (.ZN (n_8109), .A (n_8540), .B1 (n_8541), .B2 (n_8538));
NAND3_X1 i_8172 (.ZN (n_8108), .A1 (n_8541), .A2 (n_8540), .A3 (n_8538));
INV_X1 i_8171 (.ZN (n_8107), .A (n_8108));
OAI211_X1 i_8170 (.ZN (n_8106), .A (n_8110), .B (n_8120), .C1 (n_8109), .C2 (n_8107));
NAND2_X1 i_8169 (.ZN (n_8105), .A1 (n_8110), .A2 (n_8120));
NOR2_X1 i_8168 (.ZN (n_8104), .A1 (n_8109), .A2 (n_8107));
NAND2_X1 i_8167 (.ZN (n_8103), .A1 (n_8105), .A2 (n_8104));
NAND2_X1 i_8166 (.ZN (n_8102), .A1 (B_imm[21]), .A2 (A_imm[12]));
OAI21_X1 i_8165 (.ZN (n_8101), .A (n_8102), .B1 (n_8958), .B2 (n_8926));
NAND2_X1 i_8164 (.ZN (n_8100), .A1 (B_imm[15]), .A2 (A_imm[18]));
NAND4_X1 i_8163 (.ZN (n_8099), .A1 (B_imm[22]), .A2 (B_imm[21]), .A3 (A_imm[12]), .A4 (A_imm[11]));
NAND2_X1 i_8162 (.ZN (n_8098), .A1 (n_8099), .A2 (n_8100));
AOI22_X1 i_8161 (.ZN (n_8097), .A1 (n_8098), .A2 (n_8101), .B1 (A_imm[27]), .B2 (B_imm[7]));
INV_X1 i_8160 (.ZN (n_8096), .A (n_8097));
NAND4_X1 i_8159 (.ZN (n_8095), .A1 (n_8098), .A2 (B_imm[7]), .A3 (A_imm[27]), .A4 (n_8101));
INV_X1 i_8158 (.ZN (n_8094), .A (n_8095));
NAND2_X1 i_8157 (.ZN (n_8093), .A1 (B_imm[13]), .A2 (A_imm[20]));
OAI21_X1 i_8156 (.ZN (n_8092), .A (n_8093), .B1 (n_8974), .B2 (n_8511));
NAND2_X1 i_8155 (.ZN (n_8091), .A1 (B_imm[20]), .A2 (A_imm[13]));
INV_X1 i_8154 (.ZN (n_8090), .A (n_8091));
NAND4_X1 i_8153 (.ZN (n_8089), .A1 (B_imm[25]), .A2 (B_imm[13]), .A3 (A_imm[20]), .A4 (A_imm[8]));
INV_X1 i_8152 (.ZN (n_8088), .A (n_8089));
OAI21_X1 i_8151 (.ZN (n_8087), .A (n_8092), .B1 (n_8088), .B2 (n_8090));
INV_X1 i_8150 (.ZN (n_8086), .A (n_8087));
OAI21_X1 i_8149 (.ZN (n_8085), .A (n_8096), .B1 (n_8094), .B2 (n_8086));
INV_X1 i_8148 (.ZN (n_8084), .A (n_8085));
NAND2_X1 i_8147 (.ZN (n_8083), .A1 (n_8103), .A2 (n_8084));
NAND2_X1 i_8146 (.ZN (n_8082), .A1 (n_8083), .A2 (n_8106));
NAND2_X1 i_8145 (.ZN (n_8081), .A1 (n_8082), .A2 (n_8129));
NAND2_X1 i_8144 (.ZN (n_8080), .A1 (n_8081), .A2 (n_8130));
NAND2_X1 i_8143 (.ZN (n_8079), .A1 (n_8080), .A2 (n_8163));
NAND3_X1 i_8142 (.ZN (n_8078), .A1 (n_8164), .A2 (n_8130), .A3 (n_8081));
NAND3_X1 i_8141 (.ZN (n_8077), .A1 (n_8568), .A2 (n_8566), .A3 (n_8553));
INV_X1 i_8140 (.ZN (n_8076), .A (n_8553));
NAND2_X1 i_8139 (.ZN (n_8075), .A1 (n_8568), .A2 (n_8566));
NAND2_X1 i_8138 (.ZN (n_8074), .A1 (n_8075), .A2 (n_8076));
NAND2_X1 i_8137 (.ZN (n_8073), .A1 (n_8074), .A2 (n_8077));
NAND2_X1 i_8136 (.ZN (n_8072), .A1 (n_8078), .A2 (n_8073));
NAND2_X1 i_8135 (.ZN (n_8071), .A1 (n_8072), .A2 (n_8079));
NAND2_X1 i_8134 (.ZN (n_8070), .A1 (n_8071), .A2 (n_8168));
NAND2_X1 i_8133 (.ZN (n_8069), .A1 (n_8070), .A2 (n_8170));
NAND3_X1 i_8132 (.ZN (n_8068), .A1 (n_8069), .A2 (n_8181), .A3 (n_8178));
NAND2_X1 i_8131 (.ZN (n_8067), .A1 (n_8178), .A2 (n_8181));
NAND3_X1 i_8130 (.ZN (n_8066), .A1 (n_8067), .A2 (n_8170), .A3 (n_8070));
INV_X1 i_8129 (.ZN (n_8065), .A (n_8066));
NAND3_X1 i_8128 (.ZN (n_8064), .A1 (n_8358), .A2 (n_8357), .A3 (n_8356));
INV_X1 i_8127 (.ZN (n_8063), .A (n_8356));
NAND2_X1 i_8126 (.ZN (n_8062), .A1 (n_8358), .A2 (n_8357));
NAND2_X1 i_8125 (.ZN (n_8061), .A1 (n_8062), .A2 (n_8063));
NAND2_X1 i_8124 (.ZN (n_8060), .A1 (n_8061), .A2 (n_8064));
INV_X1 i_8123 (.ZN (n_8059), .A (n_8674));
OAI21_X1 i_8122 (.ZN (n_8058), .A (n_8669), .B1 (n_8673), .B2 (n_8059));
INV_X1 i_8121 (.ZN (n_8057), .A (n_8673));
INV_X1 i_8120 (.ZN (n_8056), .A (n_8669));
NAND3_X1 i_8119 (.ZN (n_8055), .A1 (n_8057), .A2 (n_8674), .A3 (n_8056));
INV_X1 i_8118 (.ZN (n_8054), .A (n_8703));
NAND2_X1 i_8117 (.ZN (n_8053), .A1 (n_8706), .A2 (n_8704));
NAND2_X1 i_8116 (.ZN (n_8052), .A1 (n_8053), .A2 (n_8054));
NAND3_X1 i_8115 (.ZN (n_8051), .A1 (n_8706), .A2 (n_8704), .A3 (n_8703));
NAND2_X1 i_8114 (.ZN (n_8050), .A1 (n_8052), .A2 (n_8051));
AOI21_X1 i_8113 (.ZN (n_8049), .A (n_8420), .B1 (n_8421), .B2 (n_8419));
NAND3_X1 i_8112 (.ZN (n_8048), .A1 (n_8421), .A2 (n_8420), .A3 (n_8419));
INV_X1 i_8111 (.ZN (n_8047), .A (n_8048));
OAI211_X2 i_8110 (.ZN (n_8046), .A (B_imm[7]), .B (A_imm[29]), .C1 (n_8047), .C2 (n_8049));
INV_X1 i_8109 (.ZN (n_8045), .A (n_8420));
NAND2_X1 i_8108 (.ZN (n_8044), .A1 (n_8421), .A2 (n_8419));
NAND2_X1 i_8107 (.ZN (n_8043), .A1 (n_8044), .A2 (n_8045));
OAI211_X1 i_8106 (.ZN (n_8042), .A (n_8043), .B (n_8048), .C1 (n_8994), .C2 (n_8573));
NAND2_X1 i_8105 (.ZN (n_8041), .A1 (B_imm[29]), .A2 (A_imm[6]));
NAND2_X1 i_8104 (.ZN (n_8040), .A1 (B_imm[12]), .A2 (A_imm[22]));
NAND2_X1 i_8103 (.ZN (n_8039), .A1 (B_imm[11]), .A2 (A_imm[23]));
NAND2_X1 i_8102 (.ZN (n_8038), .A1 (n_8039), .A2 (n_8040));
NAND2_X1 i_8101 (.ZN (n_8037), .A1 (B_imm[18]), .A2 (A_imm[16]));
NAND4_X1 i_8100 (.ZN (n_8036), .A1 (B_imm[11]), .A2 (B_imm[12]), .A3 (A_imm[23]), .A4 (A_imm[22]));
NAND2_X1 i_8099 (.ZN (n_8035), .A1 (n_8036), .A2 (n_8037));
NAND2_X1 i_8098 (.ZN (n_8034), .A1 (n_8035), .A2 (n_8038));
NAND2_X1 i_8097 (.ZN (n_8033), .A1 (n_8034), .A2 (n_8041));
INV_X1 i_8096 (.ZN (n_8032), .A (n_8041));
INV_X1 i_8095 (.ZN (n_8031), .A (n_8034));
NAND2_X1 i_8094 (.ZN (n_8030), .A1 (n_8031), .A2 (n_8032));
NAND2_X1 i_8093 (.ZN (n_8029), .A1 (A_imm[28]), .A2 (B_imm[7]));
NAND2_X1 i_8092 (.ZN (n_8028), .A1 (n_8030), .A2 (n_8029));
NAND3_X1 i_8091 (.ZN (n_8027), .A1 (n_8042), .A2 (n_8028), .A3 (n_8033));
NAND2_X1 i_8090 (.ZN (n_8026), .A1 (n_8027), .A2 (n_8046));
NAND2_X2 i_8089 (.ZN (n_8025), .A1 (n_8026), .A2 (n_8050));
NAND4_X2 i_8088 (.ZN (n_8024), .A1 (n_8027), .A2 (n_8052), .A3 (n_8051), .A4 (n_8046));
NAND2_X1 i_8087 (.ZN (n_8023), .A1 (n_8436), .A2 (n_8433));
NAND2_X1 i_8086 (.ZN (n_8022), .A1 (n_8023), .A2 (n_8434));
NAND3_X1 i_8085 (.ZN (n_8021), .A1 (n_8436), .A2 (n_8435), .A3 (n_8433));
NAND2_X1 i_8084 (.ZN (n_8020), .A1 (n_8022), .A2 (n_8021));
INV_X1 i_8083 (.ZN (n_8019), .A (n_8427));
NAND2_X1 i_8082 (.ZN (n_8018), .A1 (n_8428), .A2 (n_8426));
NAND2_X1 i_8081 (.ZN (n_8017), .A1 (n_8018), .A2 (n_8019));
NAND3_X1 i_8080 (.ZN (n_8016), .A1 (n_8428), .A2 (n_8427), .A3 (n_8426));
NAND2_X1 i_8079 (.ZN (n_8015), .A1 (n_8017), .A2 (n_8016));
NAND2_X1 i_8078 (.ZN (n_8014), .A1 (n_8020), .A2 (n_8015));
NAND4_X1 i_8077 (.ZN (n_8013), .A1 (n_8022), .A2 (n_8017), .A3 (n_8021), .A4 (n_8016));
NAND2_X1 i_8076 (.ZN (n_8012), .A1 (B_imm[9]), .A2 (A_imm[25]));
OAI21_X1 i_8075 (.ZN (n_8011), .A (n_8012), .B1 (n_8972), .B2 (n_8947));
NAND2_X1 i_8074 (.ZN (n_8010), .A1 (B_imm[24]), .A2 (A_imm[10]));
INV_X1 i_8073 (.ZN (n_8009), .A (n_8010));
NAND4_X1 i_8072 (.ZN (n_8008), .A1 (B_imm[9]), .A2 (A_imm[26]), .A3 (A_imm[25]), .A4 (B_imm[8]));
INV_X1 i_8071 (.ZN (n_8007), .A (n_8008));
OAI21_X1 i_8070 (.ZN (n_8006), .A (n_8011), .B1 (n_8007), .B2 (n_8009));
NAND2_X1 i_8069 (.ZN (n_8005), .A1 (A_imm[31]), .A2 (B_imm[3]));
OAI21_X1 i_8068 (.ZN (n_8004), .A (n_8005), .B1 (n_8821), .B2 (n_8926));
NAND2_X1 i_8067 (.ZN (n_8003), .A1 (B_imm[21]), .A2 (A_imm[13]));
INV_X1 i_8066 (.ZN (n_8002), .A (n_8003));
NAND4_X1 i_8065 (.ZN (n_8001), .A1 (B_imm[23]), .A2 (A_imm[31]), .A3 (B_imm[3]), .A4 (A_imm[11]));
INV_X1 i_8064 (.ZN (n_8000), .A (n_8001));
OAI21_X1 i_8063 (.ZN (n_7999), .A (n_8004), .B1 (n_8000), .B2 (n_8002));
NAND2_X1 i_8062 (.ZN (n_7998), .A1 (n_7999), .A2 (n_8006));
INV_X1 i_8061 (.ZN (n_7997), .A (n_8006));
INV_X1 i_8060 (.ZN (n_7996), .A (n_7999));
NAND2_X1 i_8059 (.ZN (n_7995), .A1 (n_7996), .A2 (n_7997));
OAI22_X1 i_8058 (.ZN (n_7994), .A1 (n_8829), .A2 (n_8892), .B1 (n_8958), .B2 (n_8752));
NAND2_X1 i_8057 (.ZN (n_7993), .A1 (B_imm[25]), .A2 (A_imm[9]));
INV_X1 i_8056 (.ZN (n_7992), .A (n_7993));
NAND4_X1 i_8055 (.ZN (n_7991), .A1 (B_imm[15]), .A2 (B_imm[22]), .A3 (A_imm[19]), .A4 (A_imm[12]));
INV_X1 i_8054 (.ZN (n_7990), .A (n_7991));
OAI21_X1 i_8053 (.ZN (n_7989), .A (n_7994), .B1 (n_7990), .B2 (n_7992));
NAND2_X1 i_8052 (.ZN (n_7988), .A1 (n_7995), .A2 (n_7989));
NAND3_X1 i_8051 (.ZN (n_7987), .A1 (n_8013), .A2 (n_7998), .A3 (n_7988));
NAND2_X1 i_8050 (.ZN (n_7986), .A1 (n_7987), .A2 (n_8014));
NAND2_X1 i_8049 (.ZN (n_7985), .A1 (n_7986), .A2 (n_8024));
NAND2_X1 i_8048 (.ZN (n_7984), .A1 (n_7985), .A2 (n_8025));
NAND3_X1 i_8047 (.ZN (n_7983), .A1 (n_7984), .A2 (n_8058), .A3 (n_8055));
NAND2_X1 i_8046 (.ZN (n_7982), .A1 (n_8058), .A2 (n_8055));
NAND3_X1 i_8045 (.ZN (n_7981), .A1 (n_7982), .A2 (n_8025), .A3 (n_7985));
NAND2_X1 i_8044 (.ZN (n_7980), .A1 (n_8415), .A2 (n_8431));
NAND2_X1 i_8043 (.ZN (n_7979), .A1 (n_7980), .A2 (n_8416));
INV_X1 i_8042 (.ZN (n_7978), .A (n_7979));
NAND2_X1 i_8041 (.ZN (n_7977), .A1 (B_imm[15]), .A2 (A_imm[23]));
OAI21_X1 i_8040 (.ZN (n_7976), .A (n_7977), .B1 (n_8974), .B2 (n_8927));
NAND4_X1 i_8039 (.ZN (n_7975), .A1 (B_imm[25]), .A2 (B_imm[15]), .A3 (A_imm[23]), .A4 (A_imm[13]));
NAND2_X1 i_8038 (.ZN (n_7974), .A1 (n_7976), .A2 (n_7975));
NAND3_X1 i_8037 (.ZN (n_7973), .A1 (n_7974), .A2 (B_imm[13]), .A3 (A_imm[25]));
NAND2_X1 i_8036 (.ZN (n_7972), .A1 (B_imm[13]), .A2 (A_imm[25]));
NAND3_X1 i_8035 (.ZN (n_7971), .A1 (n_7976), .A2 (n_7972), .A3 (n_7975));
NAND2_X1 i_8034 (.ZN (n_7970), .A1 (n_7973), .A2 (n_7971));
INV_X1 i_8033 (.ZN (n_7969), .A (n_8377));
OAI21_X1 i_8032 (.ZN (n_7968), .A (n_8375), .B1 (n_7969), .B2 (n_8373));
NAND3_X1 i_8031 (.ZN (n_7967), .A1 (n_8377), .A2 (n_8376), .A3 (n_8374));
NAND2_X1 i_8030 (.ZN (n_7966), .A1 (n_7968), .A2 (n_7967));
NAND2_X1 i_8029 (.ZN (n_7965), .A1 (n_7966), .A2 (n_7970));
NAND4_X1 i_8028 (.ZN (n_7964), .A1 (n_7968), .A2 (n_7973), .A3 (n_7971), .A4 (n_7967));
NAND2_X1 i_8027 (.ZN (n_7963), .A1 (n_7965), .A2 (n_7964));
NAND2_X1 i_8026 (.ZN (n_7962), .A1 (n_7963), .A2 (n_7978));
NAND3_X1 i_8025 (.ZN (n_7961), .A1 (n_7965), .A2 (n_7979), .A3 (n_7964));
NAND2_X1 i_8024 (.ZN (n_7960), .A1 (n_7962), .A2 (n_7961));
NAND2_X1 i_8023 (.ZN (n_7959), .A1 (n_7981), .A2 (n_7960));
NAND3_X1 i_8022 (.ZN (n_7958), .A1 (n_7959), .A2 (n_8060), .A3 (n_7983));
INV_X1 i_8021 (.ZN (n_7957), .A (n_7958));
AOI21_X1 i_8020 (.ZN (n_7956), .A (n_8060), .B1 (n_7959), .B2 (n_7983));
INV_X1 i_8019 (.ZN (n_7955), .A (n_7964));
OAI21_X1 i_8018 (.ZN (n_7954), .A (n_7965), .B1 (n_7979), .B2 (n_7955));
NAND2_X1 i_8017 (.ZN (n_7953), .A1 (B_imm[14]), .A2 (A_imm[25]));
INV_X1 i_8016 (.ZN (n_7952), .A (n_7953));
INV_X1 i_8015 (.ZN (n_7951), .A (n_8721));
OAI21_X1 i_8014 (.ZN (n_7950), .A (n_8722), .B1 (n_7951), .B2 (n_8724));
OAI21_X1 i_8013 (.ZN (n_7949), .A (n_7950), .B1 (n_9038), .B2 (n_8511));
NAND2_X1 i_8012 (.ZN (n_7948), .A1 (n_8721), .A2 (n_8725));
NAND4_X1 i_8011 (.ZN (n_7947), .A1 (n_7948), .A2 (B_imm[31]), .A3 (A_imm[8]), .A4 (n_8722));
NAND2_X1 i_8010 (.ZN (n_7946), .A1 (n_7949), .A2 (n_7947));
NAND2_X1 i_8009 (.ZN (n_7945), .A1 (n_7946), .A2 (n_7952));
NAND3_X1 i_8008 (.ZN (n_7944), .A1 (n_7949), .A2 (n_7953), .A3 (n_7947));
NAND2_X1 i_8007 (.ZN (n_7943), .A1 (n_7945), .A2 (n_7944));
NAND2_X1 i_8006 (.ZN (n_7942), .A1 (B_imm[30]), .A2 (A_imm[9]));
INV_X1 i_8005 (.ZN (n_7941), .A (n_7942));
NAND2_X1 i_8004 (.ZN (n_7940), .A1 (A_imm[27]), .A2 (B_imm[12]));
NAND2_X1 i_8003 (.ZN (n_7939), .A1 (n_7975), .A2 (n_7972));
NAND2_X1 i_8002 (.ZN (n_7938), .A1 (n_7939), .A2 (n_7976));
NAND2_X1 i_8001 (.ZN (n_7937), .A1 (n_7938), .A2 (n_7940));
NAND4_X1 i_8000 (.ZN (n_7936), .A1 (n_7939), .A2 (B_imm[12]), .A3 (A_imm[27]), .A4 (n_7976));
NAND2_X1 i_7999 (.ZN (n_7935), .A1 (n_7937), .A2 (n_7936));
NAND2_X1 i_7998 (.ZN (n_7934), .A1 (n_7935), .A2 (n_7941));
NAND3_X1 i_7997 (.ZN (n_7933), .A1 (n_7937), .A2 (n_7936), .A3 (n_7942));
NAND2_X1 i_7996 (.ZN (n_7932), .A1 (n_7934), .A2 (n_7933));
NAND2_X1 i_7995 (.ZN (n_7931), .A1 (n_7943), .A2 (n_7932));
NAND4_X1 i_7994 (.ZN (n_7930), .A1 (n_7945), .A2 (n_7934), .A3 (n_7944), .A4 (n_7933));
NAND2_X1 i_7993 (.ZN (n_7929), .A1 (n_7931), .A2 (n_7930));
OR2_X1 i_7992 (.ZN (n_7928), .A1 (n_7929), .A2 (n_7954));
NAND2_X1 i_7991 (.ZN (n_7927), .A1 (n_7929), .A2 (n_7954));
NAND2_X1 i_7990 (.ZN (n_7926), .A1 (n_7928), .A2 (n_7927));
INV_X1 i_7989 (.ZN (n_7925), .A (n_7926));
OAI21_X1 i_7988 (.ZN (n_7924), .A (n_7925), .B1 (n_7957), .B2 (n_7956));
NAND2_X1 i_7987 (.ZN (n_7923), .A1 (n_7959), .A2 (n_7983));
NAND3_X2 i_7986 (.ZN (n_7922), .A1 (n_7923), .A2 (n_8064), .A3 (n_8061));
NAND3_X1 i_7985 (.ZN (n_7921), .A1 (n_7922), .A2 (n_7958), .A3 (n_7926));
NAND2_X2 i_7984 (.ZN (n_7920), .A1 (n_7924), .A2 (n_7921));
OAI21_X2 i_7983 (.ZN (n_7919), .A (n_8068), .B1 (n_7920), .B2 (n_8065));
NAND2_X1 i_7982 (.ZN (n_7918), .A1 (n_7919), .A2 (n_8182));
NAND3_X1 i_7981 (.ZN (n_7917), .A1 (n_8317), .A2 (n_8185), .A3 (n_7918));
INV_X1 i_7980 (.ZN (n_7916), .A (n_8317));
NAND2_X1 i_7979 (.ZN (n_7915), .A1 (n_7918), .A2 (n_8185));
NAND2_X1 i_7978 (.ZN (n_7914), .A1 (n_7915), .A2 (n_7916));
INV_X4 i_7977 (.ZN (n_7913), .A (B_imm[14]));
INV_X2 i_7976 (.ZN (n_7912), .A (A_imm[27]));
OAI22_X1 i_7975 (.ZN (n_7911), .A1 (n_8994), .A2 (n_8795), .B1 (n_7913), .B2 (n_7912));
INV_X1 i_7974 (.ZN (n_7910), .A (n_7911));
NAND4_X1 i_7973 (.ZN (n_7909), .A1 (A_imm[29]), .A2 (B_imm[14]), .A3 (B_imm[12]), .A4 (A_imm[27]));
INV_X1 i_7972 (.ZN (n_7908), .A (n_7909));
NAND2_X1 i_7971 (.ZN (n_7907), .A1 (B_imm[18]), .A2 (A_imm[23]));
INV_X1 i_7970 (.ZN (n_7906), .A (n_7907));
OAI22_X1 i_7969 (.ZN (n_7905), .A1 (n_8794), .A2 (n_8908), .B1 (n_8767), .B2 (n_8909));
NAND4_X1 i_7968 (.ZN (n_7904), .A1 (A_imm[25]), .A2 (B_imm[17]), .A3 (B_imm[16]), .A4 (A_imm[24]));
NAND2_X1 i_7967 (.ZN (n_7903), .A1 (n_7905), .A2 (n_7904));
XNOR2_X1 i_7966 (.ZN (n_7902), .A (n_7903), .B (n_7906));
INV_X1 i_7965 (.ZN (n_7901), .A (n_7902));
OAI21_X1 i_7964 (.ZN (n_7900), .A (n_7901), .B1 (n_7910), .B2 (n_7908));
NAND3_X1 i_7963 (.ZN (n_7899), .A1 (n_7902), .A2 (n_7911), .A3 (n_7909));
NAND2_X1 i_7962 (.ZN (n_7898), .A1 (n_7900), .A2 (n_7899));
OAI21_X1 i_7961 (.ZN (n_7897), .A (n_8389), .B1 (n_8385), .B2 (n_8383));
NAND3_X1 i_7960 (.ZN (n_7896), .A1 (n_7898), .A2 (n_8391), .A3 (n_7897));
NAND2_X1 i_7959 (.ZN (n_7895), .A1 (n_7897), .A2 (n_8391));
NAND3_X1 i_7958 (.ZN (n_7894), .A1 (n_7895), .A2 (n_7900), .A3 (n_7899));
NAND2_X1 i_7957 (.ZN (n_7893), .A1 (n_7936), .A2 (n_7942));
NAND2_X1 i_7956 (.ZN (n_7892), .A1 (B_imm[28]), .A2 (A_imm[12]));
INV_X1 i_7955 (.ZN (n_7891), .A (n_7892));
NAND2_X1 i_7954 (.ZN (n_7890), .A1 (B_imm[25]), .A2 (A_imm[15]));
OAI21_X1 i_7953 (.ZN (n_7889), .A (n_7890), .B1 (n_8860), .B2 (n_8893));
NAND4_X1 i_7952 (.ZN (n_7888), .A1 (B_imm[20]), .A2 (B_imm[25]), .A3 (A_imm[20]), .A4 (A_imm[15]));
NAND2_X1 i_7951 (.ZN (n_7887), .A1 (n_7889), .A2 (n_7888));
NAND2_X1 i_7950 (.ZN (n_7886), .A1 (n_7887), .A2 (n_7891));
NAND3_X1 i_7949 (.ZN (n_7885), .A1 (n_7889), .A2 (n_7892), .A3 (n_7888));
NAND2_X1 i_7948 (.ZN (n_7884), .A1 (n_7886), .A2 (n_7885));
NAND3_X1 i_7947 (.ZN (n_7883), .A1 (n_7893), .A2 (n_7937), .A3 (n_7884));
AOI21_X1 i_7946 (.ZN (n_7882), .A (n_7884), .B1 (n_7937), .B2 (n_7893));
NAND2_X1 i_7945 (.ZN (n_7881), .A1 (A_imm[30]), .A2 (B_imm[10]));
OAI21_X1 i_7944 (.ZN (n_7880), .A (n_7883), .B1 (n_7882), .B2 (n_7881));
NAND3_X1 i_7943 (.ZN (n_7879), .A1 (n_7896), .A2 (n_7894), .A3 (n_7880));
NAND2_X1 i_7942 (.ZN (n_7878), .A1 (n_7896), .A2 (n_7894));
INV_X1 i_7941 (.ZN (n_7877), .A (n_7880));
NAND2_X1 i_7940 (.ZN (n_7876), .A1 (n_7878), .A2 (n_7877));
NAND2_X1 i_7939 (.ZN (n_7875), .A1 (n_7876), .A2 (n_7879));
NAND2_X1 i_7938 (.ZN (n_7874), .A1 (n_7930), .A2 (n_7954));
NAND2_X1 i_7937 (.ZN (n_7873), .A1 (n_7874), .A2 (n_7931));
INV_X1 i_7936 (.ZN (n_7872), .A (n_7883));
OAI21_X1 i_7935 (.ZN (n_7871), .A (n_7881), .B1 (n_7872), .B2 (n_7882));
NAND2_X1 i_7934 (.ZN (n_7870), .A1 (n_7893), .A2 (n_7937));
NAND3_X1 i_7933 (.ZN (n_7869), .A1 (n_7870), .A2 (n_7886), .A3 (n_7885));
INV_X1 i_7932 (.ZN (n_7868), .A (n_7881));
NAND3_X1 i_7931 (.ZN (n_7867), .A1 (n_7869), .A2 (n_7883), .A3 (n_7868));
NAND2_X1 i_7930 (.ZN (n_7866), .A1 (n_7871), .A2 (n_7867));
INV_X1 i_7929 (.ZN (n_7865), .A (n_7866));
NAND2_X1 i_7928 (.ZN (n_7864), .A1 (n_7873), .A2 (n_7865));
NAND3_X1 i_7927 (.ZN (n_7863), .A1 (n_7866), .A2 (n_7931), .A3 (n_7874));
NAND2_X1 i_7926 (.ZN (n_7862), .A1 (n_7947), .A2 (n_7953));
NAND2_X1 i_7925 (.ZN (n_7861), .A1 (n_8692), .A2 (n_8698));
NAND4_X2 i_7924 (.ZN (n_7860), .A1 (n_7861), .A2 (n_8696), .A3 (n_7949), .A4 (n_7862));
NAND2_X1 i_7923 (.ZN (n_7859), .A1 (n_7862), .A2 (n_7949));
NAND2_X1 i_7922 (.ZN (n_7858), .A1 (n_7861), .A2 (n_8696));
NAND2_X1 i_7921 (.ZN (n_7857), .A1 (n_7858), .A2 (n_7859));
NAND2_X1 i_7920 (.ZN (n_7856), .A1 (n_8900), .A2 (n_8898));
XNOR2_X1 i_7919 (.ZN (n_7855), .A (n_7856), .B (n_8899));
NAND3_X1 i_7918 (.ZN (n_7854), .A1 (n_7857), .A2 (n_7860), .A3 (n_7855));
NAND2_X1 i_7917 (.ZN (n_7853), .A1 (n_7857), .A2 (n_7860));
INV_X1 i_7916 (.ZN (n_7852), .A (n_7855));
NAND2_X1 i_7915 (.ZN (n_7851), .A1 (n_7853), .A2 (n_7852));
NAND2_X1 i_7914 (.ZN (n_7850), .A1 (n_7851), .A2 (n_7854));
NAND2_X1 i_7913 (.ZN (n_7849), .A1 (n_7863), .A2 (n_7850));
NAND3_X1 i_7912 (.ZN (n_7848), .A1 (n_7875), .A2 (n_7849), .A3 (n_7864));
NAND2_X1 i_7911 (.ZN (n_7847), .A1 (n_7849), .A2 (n_7864));
NAND3_X1 i_7910 (.ZN (n_7846), .A1 (n_7847), .A2 (n_7879), .A3 (n_7876));
AOI21_X1 i_7909 (.ZN (n_7845), .A (n_8367), .B1 (n_8372), .B2 (n_8365));
OAI21_X1 i_7908 (.ZN (n_7844), .A (n_8332), .B1 (n_7845), .B2 (n_8339));
NAND2_X1 i_7907 (.ZN (n_7843), .A1 (n_7844), .A2 (n_8338));
NAND2_X1 i_7906 (.ZN (n_7842), .A1 (n_7860), .A2 (n_7855));
NAND3_X1 i_7905 (.ZN (n_7841), .A1 (n_7843), .A2 (n_7842), .A3 (n_7857));
NAND2_X1 i_7904 (.ZN (n_7840), .A1 (n_7842), .A2 (n_7857));
NAND3_X1 i_7903 (.ZN (n_7839), .A1 (n_7840), .A2 (n_8338), .A3 (n_7844));
NAND2_X1 i_7902 (.ZN (n_7838), .A1 (n_8936), .A2 (n_8933));
NAND2_X1 i_7901 (.ZN (n_7837), .A1 (n_8965), .A2 (n_8962));
NAND4_X2 i_7900 (.ZN (n_7836), .A1 (n_7838), .A2 (n_7837), .A3 (n_8961), .A4 (n_8939));
NAND2_X1 i_7899 (.ZN (n_7835), .A1 (n_7838), .A2 (n_8939));
NAND2_X1 i_7898 (.ZN (n_7834), .A1 (n_7837), .A2 (n_8961));
NAND2_X1 i_7897 (.ZN (n_7833), .A1 (n_7835), .A2 (n_7834));
NAND2_X1 i_7896 (.ZN (n_7832), .A1 (B_imm[27]), .A2 (A_imm[14]));
OAI22_X1 i_7895 (.ZN (n_7831), .A1 (n_8525), .A2 (n_8906), .B1 (n_8993), .B2 (n_8946));
NAND4_X1 i_7894 (.ZN (n_7830), .A1 (B_imm[19]), .A2 (B_imm[26]), .A3 (A_imm[22]), .A4 (A_imm[15]));
NAND2_X1 i_7893 (.ZN (n_7829), .A1 (n_7831), .A2 (n_7830));
XNOR2_X1 i_7892 (.ZN (n_7828), .A (n_7829), .B (n_7832));
NAND3_X1 i_7891 (.ZN (n_7827), .A1 (n_7833), .A2 (n_7836), .A3 (n_7828));
NAND2_X1 i_7890 (.ZN (n_7826), .A1 (n_7833), .A2 (n_7836));
INV_X1 i_7889 (.ZN (n_7825), .A (n_7828));
NAND2_X1 i_7888 (.ZN (n_7824), .A1 (n_7826), .A2 (n_7825));
NAND4_X1 i_7887 (.ZN (n_7823), .A1 (n_7839), .A2 (n_7841), .A3 (n_7827), .A4 (n_7824));
NAND2_X1 i_7886 (.ZN (n_7822), .A1 (n_7839), .A2 (n_7841));
NAND2_X1 i_7885 (.ZN (n_7821), .A1 (n_7824), .A2 (n_7827));
NAND2_X1 i_7884 (.ZN (n_7820), .A1 (n_7822), .A2 (n_7821));
NAND2_X1 i_7883 (.ZN (n_7819), .A1 (n_7820), .A2 (n_7823));
NAND3_X1 i_7882 (.ZN (n_7818), .A1 (n_7846), .A2 (n_7819), .A3 (n_7848));
INV_X1 i_7881 (.ZN (n_7817), .A (n_7818));
AOI21_X1 i_7880 (.ZN (n_7816), .A (n_7819), .B1 (n_7846), .B2 (n_7848));
NAND2_X1 i_7879 (.ZN (n_7815), .A1 (n_8328), .A2 (n_8353));
NAND2_X1 i_7878 (.ZN (n_7814), .A1 (n_8769), .A2 (n_8738));
NAND4_X1 i_7877 (.ZN (n_7813), .A1 (n_7815), .A2 (n_8326), .A3 (n_8772), .A4 (n_7814));
NAND2_X1 i_7876 (.ZN (n_7812), .A1 (n_7815), .A2 (n_8326));
NAND2_X1 i_7875 (.ZN (n_7811), .A1 (n_7814), .A2 (n_8772));
NAND2_X1 i_7874 (.ZN (n_7810), .A1 (n_7812), .A2 (n_7811));
NAND2_X1 i_7873 (.ZN (n_7809), .A1 (B_imm[30]), .A2 (A_imm[11]));
INV_X1 i_7872 (.ZN (n_7808), .A (n_7809));
INV_X1 i_7871 (.ZN (n_7807), .A (n_8388));
INV_X1 i_7870 (.ZN (n_7806), .A (n_8386));
OAI21_X1 i_7869 (.ZN (n_7805), .A (n_8387), .B1 (n_7807), .B2 (n_7806));
OAI21_X1 i_7868 (.ZN (n_7804), .A (n_8346), .B1 (n_8348), .B2 (n_8343));
NAND2_X1 i_7867 (.ZN (n_7803), .A1 (n_7805), .A2 (n_7804));
INV_X1 i_7866 (.ZN (n_7802), .A (n_7805));
INV_X1 i_7865 (.ZN (n_7801), .A (n_7804));
NAND2_X1 i_7864 (.ZN (n_7800), .A1 (n_7802), .A2 (n_7801));
NAND2_X1 i_7863 (.ZN (n_7799), .A1 (n_7800), .A2 (n_7803));
NAND2_X1 i_7862 (.ZN (n_7798), .A1 (n_7799), .A2 (n_7808));
NAND3_X1 i_7861 (.ZN (n_7797), .A1 (n_7800), .A2 (n_7809), .A3 (n_7803));
NAND2_X1 i_7860 (.ZN (n_7796), .A1 (n_7798), .A2 (n_7797));
NAND2_X1 i_7859 (.ZN (n_7795), .A1 (A_imm[28]), .A2 (B_imm[13]));
INV_X1 i_7858 (.ZN (n_7794), .A (n_7795));
NAND2_X1 i_7857 (.ZN (n_7793), .A1 (n_8395), .A2 (n_8397));
NAND2_X1 i_7856 (.ZN (n_7792), .A1 (n_7793), .A2 (n_8396));
OAI21_X1 i_7855 (.ZN (n_7791), .A (n_7792), .B1 (n_9006), .B2 (n_8752));
INV_X1 i_7854 (.ZN (n_7790), .A (n_7792));
NAND3_X1 i_7853 (.ZN (n_7789), .A1 (n_7790), .A2 (B_imm[29]), .A3 (A_imm[12]));
NAND2_X1 i_7852 (.ZN (n_7788), .A1 (n_7789), .A2 (n_7791));
NAND2_X1 i_7851 (.ZN (n_7787), .A1 (n_7788), .A2 (n_7794));
NAND3_X1 i_7850 (.ZN (n_7786), .A1 (n_7789), .A2 (n_7795), .A3 (n_7791));
NAND2_X1 i_7849 (.ZN (n_7785), .A1 (n_7787), .A2 (n_7786));
NAND2_X1 i_7848 (.ZN (n_7784), .A1 (n_7796), .A2 (n_7785));
NAND4_X1 i_7847 (.ZN (n_7783), .A1 (n_7798), .A2 (n_7797), .A3 (n_7787), .A4 (n_7786));
INV_X1 i_7846 (.ZN (n_7782), .A (n_8334));
OAI21_X1 i_7845 (.ZN (n_7781), .A (n_8335), .B1 (n_8336), .B2 (n_7782));
INV_X1 i_7844 (.ZN (n_7780), .A (n_7781));
INV_X1 i_7843 (.ZN (n_7779), .A (n_7888));
OAI21_X1 i_7842 (.ZN (n_7778), .A (n_7889), .B1 (n_7779), .B2 (n_7891));
OAI21_X1 i_7841 (.ZN (n_7777), .A (n_7778), .B1 (n_9038), .B2 (n_8751));
INV_X1 i_7840 (.ZN (n_7776), .A (n_7778));
NAND3_X1 i_7839 (.ZN (n_7775), .A1 (n_7776), .A2 (B_imm[31]), .A3 (A_imm[10]));
NAND2_X1 i_7838 (.ZN (n_7774), .A1 (n_7775), .A2 (n_7777));
NAND2_X1 i_7837 (.ZN (n_7773), .A1 (n_7774), .A2 (n_7780));
NAND3_X1 i_7836 (.ZN (n_7772), .A1 (n_7775), .A2 (n_7781), .A3 (n_7777));
NAND2_X1 i_7835 (.ZN (n_7771), .A1 (n_7773), .A2 (n_7772));
AOI21_X1 i_7834 (.ZN (n_7770), .A (n_7771), .B1 (n_7784), .B2 (n_7783));
NAND3_X1 i_7833 (.ZN (n_7769), .A1 (n_7784), .A2 (n_7783), .A3 (n_7771));
INV_X1 i_7832 (.ZN (n_7768), .A (n_7769));
NOR2_X1 i_7831 (.ZN (n_7767), .A1 (n_7768), .A2 (n_7770));
NAND3_X1 i_7830 (.ZN (n_7766), .A1 (n_7810), .A2 (n_7813), .A3 (n_7767));
NAND2_X1 i_7829 (.ZN (n_7765), .A1 (n_7810), .A2 (n_7813));
INV_X1 i_7828 (.ZN (n_7764), .A (n_7767));
NAND2_X1 i_7827 (.ZN (n_7763), .A1 (n_7765), .A2 (n_7764));
NAND2_X1 i_7826 (.ZN (n_7762), .A1 (n_7763), .A2 (n_7766));
OAI21_X1 i_7825 (.ZN (n_7761), .A (n_7762), .B1 (n_7816), .B2 (n_7817));
INV_X1 i_7824 (.ZN (n_7760), .A (n_7816));
NAND4_X1 i_7823 (.ZN (n_7759), .A1 (n_7760), .A2 (n_7763), .A3 (n_7818), .A4 (n_7766));
NAND2_X1 i_7822 (.ZN (n_7758), .A1 (n_7761), .A2 (n_7759));
NAND3_X1 i_7821 (.ZN (n_7757), .A1 (n_7864), .A2 (n_7863), .A3 (n_7850));
INV_X1 i_7820 (.ZN (n_7756), .A (n_7850));
NAND2_X1 i_7819 (.ZN (n_7755), .A1 (n_7864), .A2 (n_7863));
NAND2_X1 i_7818 (.ZN (n_7754), .A1 (n_7755), .A2 (n_7756));
NAND2_X2 i_7817 (.ZN (n_7753), .A1 (n_7958), .A2 (n_7926));
NAND2_X1 i_7816 (.ZN (n_7752), .A1 (n_7753), .A2 (n_7922));
NAND3_X1 i_7815 (.ZN (n_7751), .A1 (n_7752), .A2 (n_7757), .A3 (n_7754));
NAND2_X1 i_7814 (.ZN (n_7750), .A1 (n_7754), .A2 (n_7757));
NAND3_X2 i_7813 (.ZN (n_7749), .A1 (n_7753), .A2 (n_7922), .A3 (n_7750));
INV_X1 i_7812 (.ZN (n_7748), .A (n_8911));
XNOR2_X1 i_7811 (.ZN (n_7747), .A (n_8661), .B (n_7748));
NAND3_X1 i_7810 (.ZN (n_7746), .A1 (n_8662), .A2 (n_7747), .A3 (n_8665));
NAND2_X1 i_7809 (.ZN (n_7745), .A1 (n_8662), .A2 (n_8665));
NAND2_X1 i_7808 (.ZN (n_7744), .A1 (n_7745), .A2 (n_8660));
NAND2_X1 i_7807 (.ZN (n_7743), .A1 (n_7744), .A2 (n_7746));
NAND2_X1 i_7806 (.ZN (n_7742), .A1 (n_7743), .A2 (n_7749));
NAND2_X1 i_7805 (.ZN (n_7741), .A1 (n_7742), .A2 (n_7751));
INV_X1 i_7804 (.ZN (n_7740), .A (n_7741));
NAND2_X1 i_7803 (.ZN (n_7739), .A1 (n_7758), .A2 (n_7740));
NAND3_X1 i_7802 (.ZN (n_7738), .A1 (n_7741), .A2 (n_7759), .A3 (n_7761));
NAND4_X1 i_7801 (.ZN (n_7737), .A1 (n_7914), .A2 (n_7917), .A3 (n_7739), .A4 (n_7738));
INV_X2 i_7800 (.ZN (n_7736), .A (n_7917));
AOI21_X1 i_7799 (.ZN (n_7735), .A (n_8317), .B1 (n_7918), .B2 (n_8185));
NAND2_X1 i_7798 (.ZN (n_7734), .A1 (n_7739), .A2 (n_7738));
OAI21_X2 i_7797 (.ZN (n_7733), .A (n_7734), .B1 (n_7736), .B2 (n_7735));
NAND2_X2 i_7796 (.ZN (n_7732), .A1 (n_7733), .A2 (n_7737));
AOI21_X1 i_7795 (.ZN (n_7731), .A (n_7750), .B1 (n_7922), .B2 (n_7753));
INV_X1 i_7794 (.ZN (n_7730), .A (n_7749));
INV_X1 i_7793 (.ZN (n_7729), .A (n_7743));
OAI21_X1 i_7792 (.ZN (n_7728), .A (n_7729), .B1 (n_7730), .B2 (n_7731));
NAND3_X1 i_7791 (.ZN (n_7727), .A1 (n_7751), .A2 (n_7743), .A3 (n_7749));
NAND2_X1 i_7790 (.ZN (n_7726), .A1 (n_7728), .A2 (n_7727));
INV_X1 i_7789 (.ZN (n_7725), .A (n_7726));
INV_X1 i_7788 (.ZN (n_7724), .A (n_8188));
NAND2_X1 i_7787 (.ZN (n_7723), .A1 (n_8192), .A2 (n_8202));
NAND2_X1 i_7786 (.ZN (n_7722), .A1 (n_7723), .A2 (n_7724));
NAND3_X1 i_7785 (.ZN (n_7721), .A1 (n_8188), .A2 (n_8192), .A3 (n_8202));
NAND3_X1 i_7784 (.ZN (n_7720), .A1 (n_8470), .A2 (n_8469), .A3 (n_8409));
NAND2_X1 i_7783 (.ZN (n_7719), .A1 (n_8470), .A2 (n_8469));
NAND3_X1 i_7782 (.ZN (n_7718), .A1 (n_7719), .A2 (n_8438), .A3 (n_8410));
NAND2_X1 i_7781 (.ZN (n_7717), .A1 (n_7718), .A2 (n_7720));
INV_X1 i_7780 (.ZN (n_7716), .A (n_7717));
AOI21_X1 i_7779 (.ZN (n_7715), .A (n_8411), .B1 (n_8438), .B2 (n_8437));
NAND3_X1 i_7778 (.ZN (n_7714), .A1 (n_8438), .A2 (n_8437), .A3 (n_8411));
INV_X1 i_7777 (.ZN (n_7713), .A (n_7714));
NOR2_X1 i_7776 (.ZN (n_7712), .A1 (n_7713), .A2 (n_7715));
NAND2_X1 i_7775 (.ZN (n_7711), .A1 (n_8455), .A2 (n_8458));
NAND2_X1 i_7774 (.ZN (n_7710), .A1 (n_7711), .A2 (n_8442));
NAND3_X1 i_7773 (.ZN (n_7709), .A1 (n_8441), .A2 (n_8458), .A3 (n_8455));
NAND2_X1 i_7772 (.ZN (n_7708), .A1 (n_8452), .A2 (n_8451));
NAND2_X1 i_7771 (.ZN (n_7707), .A1 (n_7708), .A2 (n_8443));
NAND3_X1 i_7770 (.ZN (n_7706), .A1 (n_8452), .A2 (n_8451), .A3 (n_8444));
NAND2_X1 i_7769 (.ZN (n_7705), .A1 (n_7707), .A2 (n_7706));
INV_X1 i_7768 (.ZN (n_7704), .A (n_8562));
NAND2_X1 i_7767 (.ZN (n_7703), .A1 (n_8563), .A2 (n_8561));
NAND2_X1 i_7766 (.ZN (n_7702), .A1 (n_7703), .A2 (n_7704));
NAND3_X1 i_7765 (.ZN (n_7701), .A1 (n_8563), .A2 (n_8561), .A3 (n_8562));
NAND2_X1 i_7764 (.ZN (n_7700), .A1 (n_7702), .A2 (n_7701));
NAND2_X1 i_7763 (.ZN (n_7699), .A1 (n_7705), .A2 (n_7700));
NAND4_X1 i_7762 (.ZN (n_7698), .A1 (n_7707), .A2 (n_7702), .A3 (n_7706), .A4 (n_7701));
NAND3_X1 i_7761 (.ZN (n_7697), .A1 (n_7698), .A2 (B_imm[5]), .A3 (A_imm[30]));
NAND2_X1 i_7760 (.ZN (n_7696), .A1 (n_7697), .A2 (n_7699));
NAND3_X1 i_7759 (.ZN (n_7695), .A1 (n_7696), .A2 (n_7710), .A3 (n_7709));
NAND2_X1 i_7758 (.ZN (n_7694), .A1 (n_7710), .A2 (n_7709));
NAND3_X1 i_7757 (.ZN (n_7693), .A1 (n_7694), .A2 (n_7699), .A3 (n_7697));
NAND2_X1 i_7756 (.ZN (n_7692), .A1 (B_imm[14]), .A2 (A_imm[20]));
INV_X2 i_7755 (.ZN (n_7691), .A (A_imm[6]));
NAND2_X1 i_7754 (.ZN (n_7690), .A1 (B_imm[19]), .A2 (A_imm[14]));
OAI21_X1 i_7753 (.ZN (n_7689), .A (n_7690), .B1 (n_9003), .B2 (n_7691));
NAND2_X1 i_7752 (.ZN (n_7688), .A1 (B_imm[29]), .A2 (A_imm[4]));
NAND4_X1 i_7751 (.ZN (n_7687), .A1 (B_imm[27]), .A2 (B_imm[19]), .A3 (A_imm[14]), .A4 (A_imm[6]));
NAND2_X1 i_7750 (.ZN (n_7686), .A1 (n_7687), .A2 (n_7688));
NAND2_X1 i_7749 (.ZN (n_7685), .A1 (n_7686), .A2 (n_7689));
NAND2_X1 i_7748 (.ZN (n_7684), .A1 (n_7685), .A2 (n_7692));
NAND4_X1 i_7747 (.ZN (n_7683), .A1 (n_7686), .A2 (B_imm[14]), .A3 (A_imm[20]), .A4 (n_7689));
INV_X1 i_7746 (.ZN (n_7682), .A (n_7683));
NAND2_X1 i_7745 (.ZN (n_7681), .A1 (B_imm[26]), .A2 (A_imm[7]));
NAND2_X1 i_7744 (.ZN (n_7680), .A1 (B_imm[28]), .A2 (A_imm[5]));
NAND2_X1 i_7743 (.ZN (n_7679), .A1 (n_7681), .A2 (n_7680));
OAI22_X1 i_7742 (.ZN (n_7678), .A1 (n_8906), .A2 (n_8880), .B1 (n_8946), .B2 (n_8909));
NAND2_X1 i_7741 (.ZN (n_7677), .A1 (A_imm[16]), .A2 (B_imm[16]));
NAND4_X1 i_7740 (.ZN (n_7676), .A1 (A_imm[22]), .A2 (B_imm[17]), .A3 (B_imm[10]), .A4 (A_imm[15]));
NAND2_X1 i_7739 (.ZN (n_7675), .A1 (n_7676), .A2 (n_7677));
NAND2_X1 i_7738 (.ZN (n_7674), .A1 (n_7675), .A2 (n_7678));
INV_X1 i_7737 (.ZN (n_7673), .A (n_7674));
NAND4_X1 i_7736 (.ZN (n_7672), .A1 (B_imm[28]), .A2 (B_imm[26]), .A3 (A_imm[7]), .A4 (A_imm[5]));
INV_X1 i_7735 (.ZN (n_7671), .A (n_7672));
OAI21_X1 i_7734 (.ZN (n_7670), .A (n_7679), .B1 (n_7671), .B2 (n_7673));
INV_X1 i_7733 (.ZN (n_7669), .A (n_7670));
OAI21_X1 i_7732 (.ZN (n_7668), .A (n_7684), .B1 (n_7682), .B2 (n_7669));
NAND4_X1 i_7731 (.ZN (n_7667), .A1 (B_imm[31]), .A2 (B_imm[30]), .A3 (A_imm[4]), .A4 (A_imm[3]));
NAND2_X1 i_7730 (.ZN (n_7666), .A1 (B_imm[30]), .A2 (A_imm[4]));
NAND2_X1 i_7729 (.ZN (n_7665), .A1 (B_imm[31]), .A2 (A_imm[3]));
NAND2_X1 i_7728 (.ZN (n_7664), .A1 (n_7665), .A2 (n_7666));
INV_X1 i_7727 (.ZN (n_7663), .A (n_8449));
OAI21_X1 i_7726 (.ZN (n_7662), .A (n_8447), .B1 (n_7663), .B2 (n_8445));
NAND3_X1 i_7725 (.ZN (n_7661), .A1 (n_8449), .A2 (n_8448), .A3 (n_8446));
NAND2_X1 i_7724 (.ZN (n_7660), .A1 (n_7662), .A2 (n_7661));
NAND2_X1 i_7723 (.ZN (n_7659), .A1 (n_7664), .A2 (n_7660));
NAND2_X1 i_7722 (.ZN (n_7658), .A1 (n_7659), .A2 (n_7667));
INV_X1 i_7721 (.ZN (n_7657), .A (n_7658));
NAND2_X1 i_7720 (.ZN (n_7656), .A1 (n_7668), .A2 (n_7657));
NAND2_X1 i_7719 (.ZN (n_7655), .A1 (n_7683), .A2 (n_7670));
NAND3_X1 i_7718 (.ZN (n_7654), .A1 (n_7655), .A2 (n_7658), .A3 (n_7684));
INV_X1 i_7717 (.ZN (n_7653), .A (n_8033));
INV_X1 i_7716 (.ZN (n_7652), .A (n_8030));
INV_X1 i_7715 (.ZN (n_7651), .A (n_8029));
OAI21_X1 i_7714 (.ZN (n_7650), .A (n_7651), .B1 (n_7652), .B2 (n_7653));
NAND3_X1 i_7713 (.ZN (n_7649), .A1 (n_8030), .A2 (n_8033), .A3 (n_8029));
NAND2_X1 i_7712 (.ZN (n_7648), .A1 (n_7650), .A2 (n_7649));
INV_X1 i_7711 (.ZN (n_7647), .A (n_7648));
NAND2_X1 i_7710 (.ZN (n_7646), .A1 (n_7654), .A2 (n_7647));
NAND3_X1 i_7709 (.ZN (n_7645), .A1 (n_7693), .A2 (n_7656), .A3 (n_7646));
NAND2_X1 i_7708 (.ZN (n_7644), .A1 (n_7645), .A2 (n_7695));
NAND2_X1 i_7707 (.ZN (n_7643), .A1 (n_7644), .A2 (n_7712));
INV_X1 i_7706 (.ZN (n_7642), .A (n_8411));
NAND2_X1 i_7705 (.ZN (n_7641), .A1 (n_8438), .A2 (n_8437));
NAND2_X1 i_7704 (.ZN (n_7640), .A1 (n_7641), .A2 (n_7642));
NAND2_X1 i_7703 (.ZN (n_7639), .A1 (n_7640), .A2 (n_7714));
NAND3_X1 i_7702 (.ZN (n_7638), .A1 (n_7639), .A2 (n_7695), .A3 (n_7645));
NAND2_X1 i_7701 (.ZN (n_7637), .A1 (n_8028), .A2 (n_8033));
NAND2_X1 i_7700 (.ZN (n_7636), .A1 (n_8046), .A2 (n_8042));
NAND2_X1 i_7699 (.ZN (n_7635), .A1 (n_7636), .A2 (n_7637));
NAND4_X1 i_7698 (.ZN (n_7634), .A1 (n_8042), .A2 (n_8046), .A3 (n_8033), .A4 (n_8028));
NAND2_X1 i_7697 (.ZN (n_7633), .A1 (n_7635), .A2 (n_7634));
INV_X1 i_7696 (.ZN (n_7632), .A (n_8285));
NAND2_X1 i_7695 (.ZN (n_7631), .A1 (n_8291), .A2 (n_8284));
NAND2_X1 i_7694 (.ZN (n_7630), .A1 (n_7631), .A2 (n_7632));
NAND3_X1 i_7693 (.ZN (n_7629), .A1 (n_8291), .A2 (n_8285), .A3 (n_8284));
NAND2_X1 i_7692 (.ZN (n_7628), .A1 (n_7630), .A2 (n_7629));
AOI21_X1 i_7691 (.ZN (n_7627), .A (n_8037), .B1 (n_8038), .B2 (n_8036));
NAND3_X1 i_7690 (.ZN (n_7626), .A1 (n_8038), .A2 (n_8036), .A3 (n_8037));
INV_X1 i_7689 (.ZN (n_7625), .A (n_7626));
OAI211_X1 i_7688 (.ZN (n_7624), .A (B_imm[5]), .B (A_imm[29]), .C1 (n_7625), .C2 (n_7627));
NAND2_X1 i_7687 (.ZN (n_7623), .A1 (A_imm[29]), .A2 (B_imm[5]));
NOR2_X1 i_7686 (.ZN (n_7622), .A1 (n_7625), .A2 (n_7627));
NAND2_X1 i_7685 (.ZN (n_7621), .A1 (n_7622), .A2 (n_7623));
NAND2_X1 i_7684 (.ZN (n_7620), .A1 (A_imm[28]), .A2 (B_imm[5]));
OAI22_X1 i_7683 (.ZN (n_7619), .A1 (n_8795), .A2 (n_8893), .B1 (n_8767), .B2 (n_8947));
NAND2_X1 i_7682 (.ZN (n_7618), .A1 (B_imm[11]), .A2 (A_imm[21]));
NAND4_X1 i_7681 (.ZN (n_7617), .A1 (B_imm[12]), .A2 (A_imm[24]), .A3 (B_imm[8]), .A4 (A_imm[20]));
NAND2_X1 i_7680 (.ZN (n_7616), .A1 (n_7617), .A2 (n_7618));
NAND2_X1 i_7679 (.ZN (n_7615), .A1 (n_7616), .A2 (n_7619));
NAND2_X1 i_7678 (.ZN (n_7614), .A1 (n_7615), .A2 (n_7620));
NAND4_X1 i_7677 (.ZN (n_7613), .A1 (n_7616), .A2 (n_7619), .A3 (B_imm[5]), .A4 (A_imm[28]));
NAND2_X1 i_7676 (.ZN (n_7612), .A1 (A_imm[25]), .A2 (B_imm[7]));
OAI21_X1 i_7675 (.ZN (n_7611), .A (n_7612), .B1 (n_8423), .B2 (n_8971));
NAND2_X1 i_7674 (.ZN (n_7610), .A1 (A_imm[26]), .A2 (B_imm[6]));
INV_X1 i_7673 (.ZN (n_7609), .A (n_7610));
NAND4_X1 i_7672 (.ZN (n_7608), .A1 (B_imm[18]), .A2 (A_imm[25]), .A3 (B_imm[7]), .A4 (A_imm[14]));
INV_X1 i_7671 (.ZN (n_7607), .A (n_7608));
OAI21_X1 i_7670 (.ZN (n_7606), .A (n_7611), .B1 (n_7607), .B2 (n_7609));
NAND2_X1 i_7669 (.ZN (n_7605), .A1 (n_7613), .A2 (n_7606));
NAND3_X1 i_7668 (.ZN (n_7604), .A1 (n_7621), .A2 (n_7614), .A3 (n_7605));
NAND2_X1 i_7667 (.ZN (n_7603), .A1 (n_7604), .A2 (n_7624));
NAND2_X1 i_7666 (.ZN (n_7602), .A1 (n_7603), .A2 (n_7628));
NAND4_X1 i_7665 (.ZN (n_7601), .A1 (n_7604), .A2 (n_7630), .A3 (n_7629), .A4 (n_7624));
AOI21_X1 i_7664 (.ZN (n_7600), .A (n_7989), .B1 (n_7995), .B2 (n_7998));
INV_X1 i_7663 (.ZN (n_7599), .A (n_7600));
NAND3_X1 i_7662 (.ZN (n_7598), .A1 (n_7995), .A2 (n_7998), .A3 (n_7989));
NAND2_X1 i_7661 (.ZN (n_7597), .A1 (n_7599), .A2 (n_7598));
NAND2_X1 i_7660 (.ZN (n_7596), .A1 (n_7601), .A2 (n_7597));
AOI21_X1 i_7659 (.ZN (n_7595), .A (n_7633), .B1 (n_7596), .B2 (n_7602));
INV_X1 i_7658 (.ZN (n_7594), .A (n_7595));
NAND3_X1 i_7657 (.ZN (n_7593), .A1 (n_7596), .A2 (n_7633), .A3 (n_7602));
NAND2_X1 i_7656 (.ZN (n_7592), .A1 (n_7988), .A2 (n_7998));
NAND3_X1 i_7655 (.ZN (n_7591), .A1 (n_7592), .A2 (n_8014), .A3 (n_8013));
NAND2_X1 i_7654 (.ZN (n_7590), .A1 (n_8014), .A2 (n_8013));
NAND3_X1 i_7653 (.ZN (n_7589), .A1 (n_7590), .A2 (n_7998), .A3 (n_7988));
NAND2_X1 i_7652 (.ZN (n_7588), .A1 (n_7589), .A2 (n_7591));
NAND2_X1 i_7651 (.ZN (n_7587), .A1 (n_7593), .A2 (n_7588));
NAND2_X1 i_7650 (.ZN (n_7586), .A1 (n_7587), .A2 (n_7594));
NAND2_X1 i_7649 (.ZN (n_7585), .A1 (n_7586), .A2 (n_7638));
NAND2_X1 i_7648 (.ZN (n_7584), .A1 (n_7585), .A2 (n_7643));
NAND2_X1 i_7647 (.ZN (n_7583), .A1 (n_7584), .A2 (n_7716));
NAND3_X1 i_7646 (.ZN (n_7582), .A1 (n_7585), .A2 (n_7717), .A3 (n_7643));
INV_X1 i_7645 (.ZN (n_7581), .A (n_7582));
NAND3_X1 i_7644 (.ZN (n_7580), .A1 (n_7983), .A2 (n_7981), .A3 (n_7960));
INV_X1 i_7643 (.ZN (n_7579), .A (n_7960));
NAND2_X1 i_7642 (.ZN (n_7578), .A1 (n_7983), .A2 (n_7981));
NAND2_X1 i_7641 (.ZN (n_7577), .A1 (n_7578), .A2 (n_7579));
NAND2_X2 i_7640 (.ZN (n_7576), .A1 (n_7577), .A2 (n_7580));
OAI21_X1 i_7639 (.ZN (n_7575), .A (n_7583), .B1 (n_7581), .B2 (n_7576));
NAND3_X2 i_7638 (.ZN (n_7574), .A1 (n_7575), .A2 (n_7722), .A3 (n_7721));
NAND2_X1 i_7637 (.ZN (n_7573), .A1 (n_7722), .A2 (n_7721));
INV_X1 i_7636 (.ZN (n_7572), .A (n_7575));
NAND2_X1 i_7635 (.ZN (n_7571), .A1 (n_7573), .A2 (n_7572));
NAND3_X1 i_7634 (.ZN (n_7570), .A1 (n_8243), .A2 (n_8245), .A3 (n_8195));
INV_X1 i_7633 (.ZN (n_7569), .A (n_8245));
OAI21_X1 i_7632 (.ZN (n_7568), .A (n_8208), .B1 (n_8201), .B2 (n_7569));
NAND2_X1 i_7631 (.ZN (n_7567), .A1 (n_7568), .A2 (n_7570));
INV_X1 i_7630 (.ZN (n_7566), .A (n_7567));
INV_X1 i_7629 (.ZN (n_7565), .A (n_8247));
NAND2_X1 i_7628 (.ZN (n_7564), .A1 (n_8273), .A2 (n_8272));
NAND2_X1 i_7627 (.ZN (n_7563), .A1 (n_7564), .A2 (n_7565));
NAND3_X1 i_7626 (.ZN (n_7562), .A1 (n_8273), .A2 (n_8247), .A3 (n_8272));
NAND3_X1 i_7625 (.ZN (n_7561), .A1 (n_8025), .A2 (n_7986), .A3 (n_8024));
NAND2_X1 i_7624 (.ZN (n_7560), .A1 (n_8025), .A2 (n_8024));
NAND3_X1 i_7623 (.ZN (n_7559), .A1 (n_7560), .A2 (n_8014), .A3 (n_7987));
NAND4_X1 i_7622 (.ZN (n_7558), .A1 (n_7563), .A2 (n_7559), .A3 (n_7562), .A4 (n_7561));
NAND2_X1 i_7621 (.ZN (n_7557), .A1 (n_7563), .A2 (n_7562));
NAND2_X1 i_7620 (.ZN (n_7556), .A1 (n_7559), .A2 (n_7561));
NAND2_X1 i_7619 (.ZN (n_7555), .A1 (n_7557), .A2 (n_7556));
NAND3_X1 i_7618 (.ZN (n_7554), .A1 (n_8295), .A2 (n_8294), .A3 (n_8282));
NAND2_X1 i_7617 (.ZN (n_7553), .A1 (n_8295), .A2 (n_8294));
NAND2_X1 i_7616 (.ZN (n_7552), .A1 (n_7553), .A2 (n_8281));
INV_X1 i_7615 (.ZN (n_7551), .A (n_8011));
OAI21_X1 i_7614 (.ZN (n_7550), .A (n_8009), .B1 (n_7551), .B2 (n_8007));
NAND3_X1 i_7613 (.ZN (n_7549), .A1 (n_8011), .A2 (n_8010), .A3 (n_8008));
NAND2_X1 i_7612 (.ZN (n_7548), .A1 (n_7550), .A2 (n_7549));
INV_X1 i_7611 (.ZN (n_7547), .A (n_8004));
OAI21_X1 i_7610 (.ZN (n_7546), .A (n_8002), .B1 (n_7547), .B2 (n_8000));
NAND3_X1 i_7609 (.ZN (n_7545), .A1 (n_8004), .A2 (n_8003), .A3 (n_8001));
NAND2_X1 i_7608 (.ZN (n_7544), .A1 (n_7546), .A2 (n_7545));
NAND2_X1 i_7607 (.ZN (n_7543), .A1 (n_7544), .A2 (n_7548));
NAND4_X1 i_7606 (.ZN (n_7542), .A1 (n_7546), .A2 (n_7550), .A3 (n_7549), .A4 (n_7545));
NAND2_X1 i_7605 (.ZN (n_7541), .A1 (n_7994), .A2 (n_7991));
NAND2_X1 i_7604 (.ZN (n_7540), .A1 (n_7541), .A2 (n_7992));
NAND3_X1 i_7603 (.ZN (n_7539), .A1 (n_7994), .A2 (n_7993), .A3 (n_7991));
NAND2_X1 i_7602 (.ZN (n_7538), .A1 (n_7540), .A2 (n_7539));
NAND2_X1 i_7601 (.ZN (n_7537), .A1 (n_7542), .A2 (n_7538));
NAND2_X1 i_7600 (.ZN (n_7536), .A1 (n_7537), .A2 (n_7543));
NAND3_X1 i_7599 (.ZN (n_7535), .A1 (n_8230), .A2 (n_8233), .A3 (n_8226));
NAND2_X1 i_7598 (.ZN (n_7534), .A1 (n_8230), .A2 (n_8233));
NAND2_X1 i_7597 (.ZN (n_7533), .A1 (n_7534), .A2 (n_8225));
NAND2_X1 i_7596 (.ZN (n_7532), .A1 (n_7533), .A2 (n_7535));
NAND2_X1 i_7595 (.ZN (n_7531), .A1 (n_7532), .A2 (n_7536));
NAND4_X1 i_7594 (.ZN (n_7530), .A1 (n_7533), .A2 (n_7537), .A3 (n_7543), .A4 (n_7535));
NAND2_X1 i_7593 (.ZN (n_7529), .A1 (B_imm[9]), .A2 (A_imm[23]));
OAI21_X1 i_7592 (.ZN (n_7528), .A (n_7529), .B1 (n_8948), .B2 (n_8511));
NAND2_X1 i_7591 (.ZN (n_7527), .A1 (A_imm[31]), .A2 (B_imm[1]));
INV_X1 i_7590 (.ZN (n_7526), .A (n_7527));
NAND4_X1 i_7589 (.ZN (n_7525), .A1 (B_imm[24]), .A2 (B_imm[9]), .A3 (A_imm[23]), .A4 (A_imm[8]));
INV_X1 i_7588 (.ZN (n_7524), .A (n_7525));
OAI21_X1 i_7587 (.ZN (n_7523), .A (n_7528), .B1 (n_7524), .B2 (n_7526));
OAI22_X1 i_7586 (.ZN (n_7522), .A1 (n_8829), .A2 (n_8955), .B1 (n_8958), .B2 (n_8751));
NAND2_X1 i_7585 (.ZN (n_7521), .A1 (B_imm[25]), .A2 (A_imm[7]));
NAND4_X1 i_7584 (.ZN (n_7520), .A1 (B_imm[15]), .A2 (B_imm[22]), .A3 (A_imm[17]), .A4 (A_imm[10]));
NAND2_X1 i_7583 (.ZN (n_7519), .A1 (n_7520), .A2 (n_7521));
NAND2_X1 i_7582 (.ZN (n_7518), .A1 (n_7519), .A2 (n_7522));
NAND2_X1 i_7581 (.ZN (n_7517), .A1 (n_7518), .A2 (n_7523));
INV_X1 i_7580 (.ZN (n_7516), .A (n_7523));
NAND3_X1 i_7579 (.ZN (n_7515), .A1 (n_7516), .A2 (n_7522), .A3 (n_7519));
NAND2_X1 i_7578 (.ZN (n_7514), .A1 (A_imm[27]), .A2 (B_imm[6]));
NAND2_X1 i_7577 (.ZN (n_7513), .A1 (n_7515), .A2 (n_7514));
AOI21_X1 i_7576 (.ZN (n_7512), .A (n_8254), .B1 (n_8255), .B2 (n_8252));
INV_X1 i_7575 (.ZN (n_7511), .A (n_7512));
NAND3_X1 i_7574 (.ZN (n_7510), .A1 (n_8255), .A2 (n_8254), .A3 (n_8252));
NAND2_X1 i_7573 (.ZN (n_7509), .A1 (n_7511), .A2 (n_7510));
NAND3_X1 i_7572 (.ZN (n_7508), .A1 (n_7513), .A2 (n_7509), .A3 (n_7517));
INV_X1 i_7571 (.ZN (n_7507), .A (n_7508));
NAND2_X1 i_7570 (.ZN (n_7506), .A1 (n_7513), .A2 (n_7517));
INV_X1 i_7569 (.ZN (n_7505), .A (n_7509));
AOI21_X1 i_7568 (.ZN (n_7504), .A (n_8289), .B1 (n_8290), .B2 (n_8287));
NAND3_X1 i_7567 (.ZN (n_7503), .A1 (n_8290), .A2 (n_8289), .A3 (n_8287));
INV_X1 i_7566 (.ZN (n_7502), .A (n_7503));
NOR2_X1 i_7565 (.ZN (n_7501), .A1 (n_7504), .A2 (n_7502));
AOI21_X1 i_7564 (.ZN (n_7500), .A (n_7501), .B1 (n_7506), .B2 (n_7505));
OAI21_X1 i_7563 (.ZN (n_7499), .A (n_7530), .B1 (n_7507), .B2 (n_7500));
AOI22_X1 i_7562 (.ZN (n_7498), .A1 (n_7499), .A2 (n_7531), .B1 (n_7554), .B2 (n_7552));
INV_X1 i_7561 (.ZN (n_7497), .A (n_7498));
NAND2_X1 i_7560 (.ZN (n_7496), .A1 (n_7552), .A2 (n_7554));
INV_X1 i_7559 (.ZN (n_7495), .A (n_7496));
NAND3_X1 i_7558 (.ZN (n_7494), .A1 (n_7499), .A2 (n_7495), .A3 (n_7531));
AOI21_X1 i_7557 (.ZN (n_7493), .A (n_8249), .B1 (n_8265), .B2 (n_8268));
NAND3_X1 i_7556 (.ZN (n_7492), .A1 (n_8265), .A2 (n_8268), .A3 (n_8249));
INV_X1 i_7555 (.ZN (n_7491), .A (n_7492));
NOR2_X1 i_7554 (.ZN (n_7490), .A1 (n_7491), .A2 (n_7493));
NAND2_X1 i_7553 (.ZN (n_7489), .A1 (n_7494), .A2 (n_7490));
NAND2_X1 i_7552 (.ZN (n_7488), .A1 (n_7489), .A2 (n_7497));
NAND2_X2 i_7551 (.ZN (n_7487), .A1 (n_7488), .A2 (n_7555));
NAND2_X1 i_7550 (.ZN (n_7486), .A1 (n_7487), .A2 (n_7558));
NAND2_X4 i_7549 (.ZN (n_7485), .A1 (n_7486), .A2 (n_7566));
NAND3_X2 i_7548 (.ZN (n_7484), .A1 (n_7487), .A2 (n_7567), .A3 (n_7558));
NAND3_X1 i_7547 (.ZN (n_7483), .A1 (n_8168), .A2 (n_8071), .A3 (n_8170));
NAND2_X1 i_7546 (.ZN (n_7482), .A1 (n_8168), .A2 (n_8170));
NAND3_X1 i_7545 (.ZN (n_7481), .A1 (n_7482), .A2 (n_8079), .A3 (n_8072));
NAND3_X1 i_7544 (.ZN (n_7480), .A1 (n_7484), .A2 (n_7483), .A3 (n_7481));
NAND2_X1 i_7543 (.ZN (n_7479), .A1 (n_7480), .A2 (n_7485));
NAND2_X1 i_7542 (.ZN (n_7478), .A1 (n_7571), .A2 (n_7479));
NAND2_X1 i_7541 (.ZN (n_7477), .A1 (n_7478), .A2 (n_7574));
NAND2_X2 i_7540 (.ZN (n_7476), .A1 (n_7477), .A2 (n_7725));
NAND3_X2 i_7539 (.ZN (n_7475), .A1 (n_7726), .A2 (n_7478), .A3 (n_7574));
INV_X1 i_7538 (.ZN (n_7474), .A (n_7919));
NAND2_X1 i_7537 (.ZN (n_7473), .A1 (n_8182), .A2 (n_8185));
NAND2_X2 i_7536 (.ZN (n_7472), .A1 (n_7473), .A2 (n_7474));
NAND3_X1 i_7535 (.ZN (n_7471), .A1 (n_7919), .A2 (n_8185), .A3 (n_8182));
NAND2_X2 i_7534 (.ZN (n_7470), .A1 (n_7472), .A2 (n_7471));
INV_X1 i_7533 (.ZN (n_7469), .A (n_7470));
NAND2_X1 i_7532 (.ZN (n_7468), .A1 (n_7469), .A2 (n_7475));
NAND2_X1 i_7531 (.ZN (n_7467), .A1 (n_7468), .A2 (n_7476));
INV_X1 i_7530 (.ZN (n_7466), .A (n_7467));
NAND2_X4 i_7529 (.ZN (n_7465), .A1 (n_7732), .A2 (n_7466));
OAI22_X1 i_7528 (.ZN (n_7464), .A1 (n_9021), .A2 (n_8971), .B1 (n_8860), .B2 (n_8906));
NAND2_X1 i_7527 (.ZN (n_7463), .A1 (B_imm[26]), .A2 (A_imm[16]));
INV_X1 i_7526 (.ZN (n_7462), .A (n_7463));
NAND4_X1 i_7525 (.ZN (n_7461), .A1 (B_imm[28]), .A2 (B_imm[20]), .A3 (A_imm[22]), .A4 (A_imm[14]));
INV_X1 i_7524 (.ZN (n_7460), .A (n_7461));
OAI21_X1 i_7523 (.ZN (n_7459), .A (n_7464), .B1 (n_7462), .B2 (n_7460));
INV_X1 i_7522 (.ZN (n_7458), .A (n_7459));
OAI22_X1 i_7521 (.ZN (n_7457), .A1 (n_9004), .A2 (n_8927), .B1 (n_7912), .B2 (n_8908));
INV_X1 i_7520 (.ZN (n_7456), .A (n_7457));
NAND4_X1 i_7519 (.ZN (n_7455), .A1 (B_imm[30]), .A2 (A_imm[27]), .A3 (B_imm[16]), .A4 (A_imm[13]));
INV_X1 i_7518 (.ZN (n_7454), .A (n_7455));
OAI21_X1 i_7517 (.ZN (n_7453), .A (n_7458), .B1 (n_7456), .B2 (n_7454));
NAND3_X1 i_7516 (.ZN (n_7452), .A1 (n_7457), .A2 (n_7459), .A3 (n_7455));
NAND2_X1 i_7515 (.ZN (n_7451), .A1 (n_7453), .A2 (n_7452));
OAI22_X1 i_7514 (.ZN (n_7450), .A1 (n_8958), .A2 (n_8893), .B1 (n_8957), .B2 (n_8859));
NAND2_X1 i_7513 (.ZN (n_7449), .A1 (B_imm[25]), .A2 (A_imm[17]));
INV_X1 i_7512 (.ZN (n_7448), .A (n_7449));
NAND4_X1 i_7511 (.ZN (n_7447), .A1 (B_imm[22]), .A2 (B_imm[21]), .A3 (A_imm[21]), .A4 (A_imm[20]));
INV_X1 i_7510 (.ZN (n_7446), .A (n_7447));
OAI21_X1 i_7509 (.ZN (n_7445), .A (n_7450), .B1 (n_7448), .B2 (n_7446));
INV_X1 i_7508 (.ZN (n_7444), .A (n_7445));
OAI22_X1 i_7507 (.ZN (n_7443), .A1 (n_8948), .A2 (n_8956), .B1 (n_9037), .B2 (n_8849));
NAND2_X1 i_7506 (.ZN (n_7442), .A1 (B_imm[23]), .A2 (A_imm[19]));
INV_X1 i_7505 (.ZN (n_7441), .A (n_7442));
NAND4_X1 i_7504 (.ZN (n_7440), .A1 (B_imm[24]), .A2 (opt_ipoPP_0), .A3 (B_imm[11]), .A4 (A_imm[18]));
INV_X1 i_7503 (.ZN (n_7439), .A (n_7440));
OAI21_X1 i_7502 (.ZN (n_7438), .A (n_7443), .B1 (n_7441), .B2 (n_7439));
OAI22_X1 i_7501 (.ZN (n_7437), .A1 (n_8909), .A2 (n_8794), .B1 (n_8972), .B2 (n_8908));
NAND2_X1 i_7500 (.ZN (n_7436), .A1 (B_imm[18]), .A2 (A_imm[24]));
INV_X1 i_7499 (.ZN (n_7435), .A (n_7436));
NAND4_X1 i_7498 (.ZN (n_7434), .A1 (A_imm[26]), .A2 (A_imm[25]), .A3 (B_imm[17]), .A4 (B_imm[16]));
INV_X1 i_7497 (.ZN (n_7433), .A (n_7434));
OAI21_X1 i_7496 (.ZN (n_7432), .A (n_7437), .B1 (n_7435), .B2 (n_7433));
NAND2_X1 i_7495 (.ZN (n_7431), .A1 (n_7438), .A2 (n_7432));
INV_X1 i_7494 (.ZN (n_7430), .A (n_7438));
INV_X1 i_7493 (.ZN (n_7429), .A (n_7432));
NAND2_X1 i_7492 (.ZN (n_7428), .A1 (n_7430), .A2 (n_7429));
NAND2_X1 i_7491 (.ZN (n_7427), .A1 (n_7428), .A2 (n_7431));
NAND2_X1 i_7490 (.ZN (n_7426), .A1 (n_7427), .A2 (n_7444));
NAND3_X1 i_7489 (.ZN (n_7425), .A1 (n_7428), .A2 (n_7445), .A3 (n_7431));
NAND2_X1 i_7488 (.ZN (n_7424), .A1 (n_7426), .A2 (n_7425));
NAND2_X1 i_7487 (.ZN (n_7423), .A1 (n_7451), .A2 (n_7424));
NAND4_X1 i_7486 (.ZN (n_7422), .A1 (n_7453), .A2 (n_7426), .A3 (n_7452), .A4 (n_7425));
NAND2_X1 i_7485 (.ZN (n_7421), .A1 (n_7437), .A2 (n_7434));
XNOR2_X1 i_7484 (.ZN (n_7420), .A (n_7421), .B (n_7435));
NAND3_X1 i_7483 (.ZN (n_7419), .A1 (n_7420), .A2 (B_imm[13]), .A3 (A_imm[29]));
XNOR2_X1 i_7482 (.ZN (n_7418), .A (n_7421), .B (n_7436));
OAI21_X1 i_7481 (.ZN (n_7417), .A (n_7418), .B1 (n_8973), .B2 (n_8994));
INV_X1 i_7480 (.ZN (n_7416), .A (n_7417));
INV_X1 i_7479 (.ZN (n_7415), .A (n_7789));
OAI21_X1 i_7478 (.ZN (n_7414), .A (n_7791), .B1 (n_7415), .B2 (n_7794));
OAI21_X1 i_7477 (.ZN (n_7413), .A (n_7419), .B1 (n_7416), .B2 (n_7414));
NAND2_X1 i_7476 (.ZN (n_7412), .A1 (n_7413), .A2 (n_7422));
NAND2_X1 i_7475 (.ZN (n_7411), .A1 (n_7412), .A2 (n_7423));
NAND2_X1 i_7474 (.ZN (n_7410), .A1 (B_imm[23]), .A2 (A_imm[21]));
OAI22_X1 i_7473 (.ZN (n_7409), .A1 (n_8423), .A2 (n_8972), .B1 (n_8948), .B2 (n_8893));
NAND4_X1 i_7472 (.ZN (n_7408), .A1 (B_imm[24]), .A2 (B_imm[18]), .A3 (A_imm[26]), .A4 (A_imm[20]));
NAND2_X1 i_7471 (.ZN (n_7407), .A1 (n_7409), .A2 (n_7408));
XNOR2_X1 i_7470 (.ZN (n_7406), .A (n_7407), .B (n_7410));
OAI22_X1 i_7469 (.ZN (n_7405), .A1 (n_9006), .A2 (n_8971), .B1 (n_9003), .B2 (n_8858));
NAND2_X1 i_7468 (.ZN (n_7404), .A1 (A_imm[28]), .A2 (B_imm[15]));
INV_X1 i_7467 (.ZN (n_7403), .A (n_7404));
NAND4_X1 i_7466 (.ZN (n_7402), .A1 (B_imm[29]), .A2 (B_imm[27]), .A3 (A_imm[16]), .A4 (A_imm[14]));
INV_X1 i_7465 (.ZN (n_7401), .A (n_7402));
OAI21_X1 i_7464 (.ZN (n_7400), .A (n_7405), .B1 (n_7403), .B2 (n_7401));
INV_X1 i_7463 (.ZN (n_7399), .A (n_7400));
NAND3_X1 i_7462 (.ZN (n_7398), .A1 (n_7399), .A2 (B_imm[15]), .A3 (A_imm[29]));
OAI21_X1 i_7461 (.ZN (n_7397), .A (n_7400), .B1 (n_8829), .B2 (n_8994));
NAND3_X1 i_7460 (.ZN (n_7396), .A1 (n_7406), .A2 (n_7398), .A3 (n_7397));
INV_X1 i_7459 (.ZN (n_7395), .A (n_7406));
INV_X1 i_7458 (.ZN (n_7394), .A (n_7398));
INV_X1 i_7457 (.ZN (n_7393), .A (n_7397));
OAI21_X1 i_7456 (.ZN (n_7392), .A (n_7395), .B1 (n_7394), .B2 (n_7393));
NAND2_X1 i_7455 (.ZN (n_7391), .A1 (n_7392), .A2 (n_7396));
NAND2_X1 i_7454 (.ZN (n_7390), .A1 (A_imm[30]), .A2 (B_imm[13]));
INV_X1 i_7453 (.ZN (n_7389), .A (n_7390));
NAND2_X1 i_7452 (.ZN (n_7388), .A1 (B_imm[31]), .A2 (A_imm[11]));
INV_X1 i_7451 (.ZN (n_7387), .A (n_7832));
INV_X1 i_7450 (.ZN (n_7386), .A (n_7830));
OAI21_X1 i_7449 (.ZN (n_7385), .A (n_7831), .B1 (n_7387), .B2 (n_7386));
NAND2_X1 i_7448 (.ZN (n_7384), .A1 (n_7385), .A2 (n_7388));
NAND2_X1 i_7447 (.ZN (n_7383), .A1 (B_imm[14]), .A2 (A_imm[28]));
OAI21_X1 i_7446 (.ZN (n_7382), .A (n_7383), .B1 (n_7385), .B2 (n_7388));
NAND2_X1 i_7445 (.ZN (n_7381), .A1 (n_7382), .A2 (n_7384));
INV_X1 i_7444 (.ZN (n_7380), .A (n_7381));
NAND2_X1 i_7443 (.ZN (n_7379), .A1 (n_7380), .A2 (n_7389));
NOR2_X1 i_7442 (.ZN (n_7378), .A1 (n_7380), .A2 (n_7389));
INV_X1 i_7441 (.ZN (n_7377), .A (n_7378));
NAND2_X1 i_7440 (.ZN (n_7376), .A1 (n_7405), .A2 (n_7402));
XNOR2_X1 i_7439 (.ZN (n_7375), .A (n_7376), .B (n_7404));
INV_X1 i_7438 (.ZN (n_7374), .A (n_7375));
NAND2_X1 i_7437 (.ZN (n_7373), .A1 (n_7377), .A2 (n_7374));
NAND2_X1 i_7436 (.ZN (n_7372), .A1 (n_7373), .A2 (n_7379));
NAND2_X1 i_7435 (.ZN (n_7371), .A1 (n_7372), .A2 (n_7391));
NAND4_X1 i_7434 (.ZN (n_7370), .A1 (n_7373), .A2 (n_7392), .A3 (n_7396), .A4 (n_7379));
NAND3_X1 i_7433 (.ZN (n_7369), .A1 (n_7371), .A2 (n_7411), .A3 (n_7370));
NAND2_X1 i_7432 (.ZN (n_7368), .A1 (n_7371), .A2 (n_7370));
NAND3_X1 i_7431 (.ZN (n_7367), .A1 (n_7368), .A2 (n_7423), .A3 (n_7412));
OAI21_X1 i_7430 (.ZN (n_7366), .A (n_8857), .B1 (n_8861), .B2 (n_8854));
OAI22_X1 i_7429 (.ZN (n_7365), .A1 (n_9004), .A2 (n_8752), .B1 (n_7912), .B2 (n_8829));
NAND4_X1 i_7428 (.ZN (n_7364), .A1 (B_imm[30]), .A2 (A_imm[27]), .A3 (B_imm[15]), .A4 (A_imm[12]));
NAND2_X1 i_7427 (.ZN (n_7363), .A1 (n_7365), .A2 (n_7364));
XNOR2_X1 i_7426 (.ZN (n_7362), .A (n_7363), .B (n_7366));
INV_X1 i_7425 (.ZN (n_7361), .A (n_7362));
NAND2_X1 i_7424 (.ZN (n_7360), .A1 (n_8870), .A2 (n_8885));
NAND2_X1 i_7423 (.ZN (n_7359), .A1 (n_7360), .A2 (n_8883));
NAND2_X1 i_7422 (.ZN (n_7358), .A1 (n_7361), .A2 (n_7359));
NAND3_X1 i_7421 (.ZN (n_7357), .A1 (n_7362), .A2 (n_8883), .A3 (n_7360));
INV_X1 i_7420 (.ZN (n_7356), .A (n_7385));
NAND3_X1 i_7419 (.ZN (n_7355), .A1 (n_7356), .A2 (B_imm[31]), .A3 (A_imm[11]));
AOI21_X1 i_7418 (.ZN (n_7354), .A (n_7383), .B1 (n_7355), .B2 (n_7384));
INV_X1 i_7417 (.ZN (n_7353), .A (n_7354));
NAND2_X1 i_7416 (.ZN (n_7352), .A1 (n_7355), .A2 (n_7384));
INV_X1 i_7415 (.ZN (n_7351), .A (n_7352));
NAND2_X1 i_7414 (.ZN (n_7350), .A1 (n_7351), .A2 (n_7383));
NAND2_X1 i_7413 (.ZN (n_7349), .A1 (n_7353), .A2 (n_7350));
NAND2_X1 i_7412 (.ZN (n_7348), .A1 (n_7357), .A2 (n_7349));
NAND2_X1 i_7411 (.ZN (n_7347), .A1 (n_7348), .A2 (n_7358));
INV_X1 i_7410 (.ZN (n_7346), .A (n_7366));
INV_X1 i_7409 (.ZN (n_7345), .A (n_7364));
OAI21_X1 i_7408 (.ZN (n_7344), .A (n_7365), .B1 (n_7346), .B2 (n_7345));
INV_X1 i_7407 (.ZN (n_7343), .A (n_7344));
NAND2_X1 i_7406 (.ZN (n_7342), .A1 (n_8878), .A2 (n_8881));
NAND2_X1 i_7405 (.ZN (n_7341), .A1 (n_7342), .A2 (n_8879));
NAND2_X1 i_7404 (.ZN (n_7340), .A1 (n_7904), .A2 (n_7907));
NAND2_X1 i_7403 (.ZN (n_7339), .A1 (n_7340), .A2 (n_7905));
NAND2_X1 i_7402 (.ZN (n_7338), .A1 (n_7341), .A2 (n_7339));
OAI21_X1 i_7401 (.ZN (n_7337), .A (n_8891), .B1 (n_8894), .B2 (n_8888));
NAND4_X1 i_7400 (.ZN (n_7336), .A1 (n_7342), .A2 (n_8879), .A3 (n_7905), .A4 (n_7340));
NAND2_X1 i_7399 (.ZN (n_7335), .A1 (n_7336), .A2 (n_7337));
NAND2_X1 i_7398 (.ZN (n_7334), .A1 (B_imm[19]), .A2 (A_imm[24]));
OAI22_X1 i_7397 (.ZN (n_7333), .A1 (n_9021), .A2 (n_8946), .B1 (n_8993), .B2 (n_8955));
NAND4_X1 i_7396 (.ZN (n_7332), .A1 (B_imm[28]), .A2 (B_imm[26]), .A3 (A_imm[17]), .A4 (A_imm[15]));
NAND2_X1 i_7395 (.ZN (n_7331), .A1 (n_7333), .A2 (n_7332));
XNOR2_X1 i_7394 (.ZN (n_7330), .A (n_7331), .B (n_7334));
INV_X1 i_7393 (.ZN (n_7329), .A (n_7330));
NAND3_X1 i_7392 (.ZN (n_7328), .A1 (n_7329), .A2 (n_7338), .A3 (n_7335));
NAND2_X1 i_7391 (.ZN (n_7327), .A1 (n_7335), .A2 (n_7338));
NAND2_X1 i_7390 (.ZN (n_7326), .A1 (n_7330), .A2 (n_7327));
NAND2_X1 i_7389 (.ZN (n_7325), .A1 (n_7328), .A2 (n_7326));
NAND2_X1 i_7388 (.ZN (n_7324), .A1 (n_7325), .A2 (n_7343));
NAND3_X1 i_7387 (.ZN (n_7323), .A1 (n_7328), .A2 (n_7344), .A3 (n_7326));
NAND2_X1 i_7386 (.ZN (n_7322), .A1 (n_7324), .A2 (n_7323));
NAND2_X1 i_7385 (.ZN (n_7321), .A1 (n_7347), .A2 (n_7322));
NAND4_X1 i_7384 (.ZN (n_7320), .A1 (n_7348), .A2 (n_7358), .A3 (n_7323), .A4 (n_7324));
NAND2_X2 i_7383 (.ZN (n_7319), .A1 (n_7836), .A2 (n_7828));
NAND2_X1 i_7382 (.ZN (n_7318), .A1 (n_7319), .A2 (n_7833));
NAND2_X1 i_7381 (.ZN (n_7317), .A1 (n_8863), .A2 (n_8850));
NAND2_X1 i_7380 (.ZN (n_7316), .A1 (n_7317), .A2 (n_8848));
NAND2_X2 i_7379 (.ZN (n_7315), .A1 (n_7318), .A2 (n_7316));
NAND4_X2 i_7378 (.ZN (n_7314), .A1 (n_7319), .A2 (n_7317), .A3 (n_8848), .A4 (n_7833));
INV_X1 i_7377 (.ZN (n_7313), .A (n_7314));
INV_X1 i_7376 (.ZN (n_7312), .A (n_7414));
NAND2_X1 i_7375 (.ZN (n_7311), .A1 (n_7417), .A2 (n_7419));
NAND2_X1 i_7374 (.ZN (n_7310), .A1 (n_7311), .A2 (n_7312));
NAND3_X1 i_7373 (.ZN (n_7309), .A1 (n_7417), .A2 (n_7419), .A3 (n_7414));
NAND2_X1 i_7372 (.ZN (n_7308), .A1 (n_7310), .A2 (n_7309));
OAI21_X1 i_7371 (.ZN (n_7307), .A (n_7315), .B1 (n_7313), .B2 (n_7308));
INV_X1 i_7370 (.ZN (n_7306), .A (n_7307));
NAND2_X1 i_7369 (.ZN (n_7305), .A1 (n_7320), .A2 (n_7306));
NAND2_X1 i_7368 (.ZN (n_7304), .A1 (n_7305), .A2 (n_7321));
NAND3_X1 i_7367 (.ZN (n_7303), .A1 (n_7304), .A2 (n_7369), .A3 (n_7367));
NAND2_X1 i_7366 (.ZN (n_7302), .A1 (n_7367), .A2 (n_7369));
NAND3_X1 i_7365 (.ZN (n_7301), .A1 (n_7302), .A2 (n_7321), .A3 (n_7305));
INV_X1 i_7364 (.ZN (n_7300), .A (n_7443));
OAI21_X1 i_7363 (.ZN (n_7299), .A (n_7441), .B1 (n_7300), .B2 (n_7439));
NAND3_X1 i_7362 (.ZN (n_7298), .A1 (n_7443), .A2 (n_7442), .A3 (n_7440));
NAND2_X1 i_7361 (.ZN (n_7297), .A1 (n_7299), .A2 (n_7298));
INV_X1 i_7360 (.ZN (n_7296), .A (n_7450));
OAI21_X1 i_7359 (.ZN (n_7295), .A (n_7448), .B1 (n_7296), .B2 (n_7446));
NAND3_X1 i_7358 (.ZN (n_7294), .A1 (n_7450), .A2 (n_7449), .A3 (n_7447));
NAND2_X1 i_7357 (.ZN (n_7293), .A1 (n_7295), .A2 (n_7294));
NAND2_X1 i_7356 (.ZN (n_7292), .A1 (n_7293), .A2 (n_7297));
NAND4_X1 i_7355 (.ZN (n_7291), .A1 (n_7295), .A2 (n_7299), .A3 (n_7298), .A4 (n_7294));
NAND2_X1 i_7354 (.ZN (n_7290), .A1 (n_7464), .A2 (n_7461));
XNOR2_X1 i_7353 (.ZN (n_7289), .A (n_7290), .B (n_7462));
NAND2_X1 i_7352 (.ZN (n_7288), .A1 (n_7289), .A2 (n_7291));
NAND2_X1 i_7351 (.ZN (n_7287), .A1 (n_7288), .A2 (n_7292));
NAND2_X1 i_7350 (.ZN (n_7286), .A1 (n_7800), .A2 (n_7809));
NAND2_X1 i_7349 (.ZN (n_7285), .A1 (B_imm[29]), .A2 (A_imm[13]));
OAI22_X1 i_7348 (.ZN (n_7284), .A1 (CLOCK_opt_ipo_n433), .A2 (n_8946), .B1 (n_8525), .B2 (n_8907));
NAND4_X1 i_7347 (.ZN (n_7283), .A1 (B_imm[27]), .A2 (B_imm[19]), .A3 (A_imm[23]), .A4 (A_imm[15]));
NAND2_X1 i_7346 (.ZN (n_7282), .A1 (n_7284), .A2 (n_7283));
XNOR2_X1 i_7345 (.ZN (n_7281), .A (n_7282), .B (n_7285));
INV_X1 i_7344 (.ZN (n_7280), .A (n_7281));
NAND3_X1 i_7343 (.ZN (n_7279), .A1 (n_7280), .A2 (n_7803), .A3 (n_7286));
NAND2_X1 i_7342 (.ZN (n_7278), .A1 (A_imm[30]), .A2 (B_imm[12]));
NAND2_X1 i_7341 (.ZN (n_7277), .A1 (n_7286), .A2 (n_7803));
NAND2_X1 i_7340 (.ZN (n_7276), .A1 (n_7277), .A2 (n_7281));
INV_X1 i_7339 (.ZN (n_7275), .A (n_7276));
OAI21_X1 i_7338 (.ZN (n_7274), .A (n_7279), .B1 (n_7275), .B2 (n_7278));
NAND2_X1 i_7337 (.ZN (n_7273), .A1 (n_7274), .A2 (n_7287));
INV_X1 i_7336 (.ZN (n_7272), .A (n_7287));
OAI211_X1 i_7335 (.ZN (n_7271), .A (n_7272), .B (n_7279), .C1 (n_7275), .C2 (n_7278));
NAND2_X1 i_7334 (.ZN (n_7270), .A1 (A_imm[29]), .A2 (B_imm[14]));
INV_X1 i_7333 (.ZN (n_7269), .A (n_7270));
NAND2_X1 i_7332 (.ZN (n_7268), .A1 (n_7283), .A2 (n_7285));
NAND2_X1 i_7331 (.ZN (n_7267), .A1 (n_7268), .A2 (n_7284));
OAI21_X1 i_7330 (.ZN (n_7266), .A (n_7267), .B1 (n_9038), .B2 (n_8752));
INV_X1 i_7329 (.ZN (n_7265), .A (n_7267));
NAND3_X1 i_7328 (.ZN (n_7264), .A1 (n_7265), .A2 (B_imm[31]), .A3 (A_imm[12]));
NAND2_X1 i_7327 (.ZN (n_7263), .A1 (n_7264), .A2 (n_7266));
XNOR2_X1 i_7326 (.ZN (n_7262), .A (n_7263), .B (n_7269));
INV_X1 i_7325 (.ZN (n_7261), .A (n_7262));
NAND3_X1 i_7324 (.ZN (n_7260), .A1 (n_7273), .A2 (n_7271), .A3 (n_7261));
INV_X1 i_7323 (.ZN (n_7259), .A (n_7260));
AOI21_X1 i_7322 (.ZN (n_7258), .A (n_7261), .B1 (n_7273), .B2 (n_7271));
NAND3_X1 i_7321 (.ZN (n_7257), .A1 (n_7413), .A2 (n_7423), .A3 (n_7422));
INV_X1 i_7320 (.ZN (n_7256), .A (n_7413));
NAND2_X1 i_7319 (.ZN (n_7255), .A1 (n_7423), .A2 (n_7422));
NAND2_X1 i_7318 (.ZN (n_7254), .A1 (n_7255), .A2 (n_7256));
NAND2_X1 i_7317 (.ZN (n_7253), .A1 (n_7254), .A2 (n_7257));
INV_X1 i_7316 (.ZN (n_7252), .A (n_7253));
OAI21_X2 i_7315 (.ZN (n_7251), .A (n_7252), .B1 (n_7259), .B2 (n_7258));
NAND2_X1 i_7314 (.ZN (n_7250), .A1 (n_7273), .A2 (n_7271));
NAND2_X1 i_7313 (.ZN (n_7249), .A1 (n_7250), .A2 (n_7262));
NAND3_X1 i_7312 (.ZN (n_7248), .A1 (n_7249), .A2 (n_7260), .A3 (n_7253));
NAND2_X1 i_7311 (.ZN (n_7247), .A1 (n_7783), .A2 (n_7771));
NAND2_X1 i_7310 (.ZN (n_7246), .A1 (n_7247), .A2 (n_7784));
INV_X1 i_7309 (.ZN (n_7245), .A (n_7289));
NAND2_X1 i_7308 (.ZN (n_7244), .A1 (n_7292), .A2 (n_7291));
NAND2_X1 i_7307 (.ZN (n_7243), .A1 (n_7244), .A2 (n_7245));
NAND3_X1 i_7306 (.ZN (n_7242), .A1 (n_7289), .A2 (n_7292), .A3 (n_7291));
NAND3_X1 i_7305 (.ZN (n_7241), .A1 (n_7246), .A2 (n_7243), .A3 (n_7242));
NAND2_X1 i_7304 (.ZN (n_7240), .A1 (n_7243), .A2 (n_7242));
NAND3_X1 i_7303 (.ZN (n_7239), .A1 (n_7247), .A2 (n_7784), .A3 (n_7240));
NAND2_X1 i_7302 (.ZN (n_7238), .A1 (n_7896), .A2 (n_7880));
NAND2_X1 i_7301 (.ZN (n_7237), .A1 (n_7238), .A2 (n_7894));
NAND2_X1 i_7300 (.ZN (n_7236), .A1 (n_7237), .A2 (n_7239));
NAND2_X1 i_7299 (.ZN (n_7235), .A1 (n_7236), .A2 (n_7241));
NAND2_X1 i_7298 (.ZN (n_7234), .A1 (n_7248), .A2 (n_7235));
NAND2_X1 i_7297 (.ZN (n_7233), .A1 (n_7234), .A2 (n_7251));
NAND3_X1 i_7296 (.ZN (n_7232), .A1 (n_7233), .A2 (n_7303), .A3 (n_7301));
NAND2_X1 i_7295 (.ZN (n_7231), .A1 (n_7303), .A2 (n_7301));
INV_X1 i_7294 (.ZN (n_7230), .A (n_7233));
NAND2_X1 i_7293 (.ZN (n_7229), .A1 (n_7231), .A2 (n_7230));
NAND2_X1 i_7292 (.ZN (n_7228), .A1 (n_7229), .A2 (n_7232));
NAND3_X1 i_7291 (.ZN (n_7227), .A1 (n_7251), .A2 (n_7248), .A3 (n_7235));
INV_X1 i_7290 (.ZN (n_7226), .A (n_7235));
NAND2_X1 i_7289 (.ZN (n_7225), .A1 (n_7251), .A2 (n_7248));
NAND2_X1 i_7288 (.ZN (n_7224), .A1 (n_7225), .A2 (n_7226));
NAND3_X1 i_7287 (.ZN (n_7223), .A1 (n_7321), .A2 (n_7320), .A3 (n_7307));
NAND2_X1 i_7286 (.ZN (n_7222), .A1 (n_7321), .A2 (n_7320));
NAND2_X1 i_7285 (.ZN (n_7221), .A1 (n_7222), .A2 (n_7306));
NAND2_X1 i_7284 (.ZN (n_7220), .A1 (n_7221), .A2 (n_7223));
NAND3_X1 i_7283 (.ZN (n_7219), .A1 (n_7224), .A2 (n_7220), .A3 (n_7227));
NAND2_X1 i_7282 (.ZN (n_7218), .A1 (n_7224), .A2 (n_7227));
INV_X1 i_7281 (.ZN (n_7217), .A (n_7220));
NAND2_X1 i_7280 (.ZN (n_7216), .A1 (n_7218), .A2 (n_7217));
NAND3_X1 i_7279 (.ZN (n_7215), .A1 (n_7241), .A2 (n_7239), .A3 (n_7237));
NAND2_X1 i_7278 (.ZN (n_7214), .A1 (n_7241), .A2 (n_7239));
NAND3_X1 i_7277 (.ZN (n_7213), .A1 (n_7214), .A2 (n_7894), .A3 (n_7238));
NAND2_X1 i_7276 (.ZN (n_7212), .A1 (n_7213), .A2 (n_7215));
INV_X1 i_7275 (.ZN (n_7211), .A (n_7212));
NAND2_X1 i_7274 (.ZN (n_7210), .A1 (n_7813), .A2 (n_7767));
NAND2_X1 i_7273 (.ZN (n_7209), .A1 (n_7210), .A2 (n_7810));
NAND2_X1 i_7272 (.ZN (n_7208), .A1 (n_7209), .A2 (n_7211));
NAND3_X1 i_7271 (.ZN (n_7207), .A1 (n_7212), .A2 (n_7810), .A3 (n_7210));
NAND2_X1 i_7270 (.ZN (n_7206), .A1 (n_7819), .A2 (n_7848));
NAND2_X1 i_7269 (.ZN (n_7205), .A1 (n_7206), .A2 (n_7846));
NAND2_X1 i_7268 (.ZN (n_7204), .A1 (n_7207), .A2 (n_7205));
NAND2_X1 i_7267 (.ZN (n_7203), .A1 (n_7204), .A2 (n_7208));
NAND2_X1 i_7266 (.ZN (n_7202), .A1 (n_7216), .A2 (n_7203));
AOI21_X1 i_7265 (.ZN (n_7201), .A (n_7228), .B1 (n_7202), .B2 (n_7219));
INV_X1 i_7264 (.ZN (n_7200), .A (n_7201));
NAND3_X1 i_7263 (.ZN (n_7199), .A1 (n_7202), .A2 (n_7228), .A3 (n_7219));
OAI21_X1 i_7262 (.ZN (n_7198), .A (n_7457), .B1 (n_7458), .B2 (n_7454));
INV_X1 i_7261 (.ZN (n_7197), .A (n_7198));
NAND2_X1 i_7260 (.ZN (n_7196), .A1 (B_imm[28]), .A2 (A_imm[16]));
INV_X1 i_7259 (.ZN (n_7195), .A (n_7196));
OAI22_X1 i_7258 (.ZN (n_7194), .A1 (n_8860), .A2 (n_8767), .B1 (n_8973), .B2 (n_9037));
NAND4_X1 i_7257 (.ZN (n_7193), .A1 (B_imm[20]), .A2 (B_imm[13]), .A3 (A_imm[31]), .A4 (A_imm[24]));
NAND2_X1 i_7256 (.ZN (n_7192), .A1 (n_7194), .A2 (n_7193));
XNOR2_X1 i_7255 (.ZN (n_7191), .A (n_7192), .B (n_7195));
INV_X1 i_7254 (.ZN (n_7190), .A (n_7191));
OAI21_X1 i_7253 (.ZN (n_7189), .A (n_7190), .B1 (n_7913), .B2 (n_9005));
NAND3_X1 i_7252 (.ZN (n_7188), .A1 (n_7191), .A2 (B_imm[14]), .A3 (A_imm[30]));
AOI21_X1 i_7251 (.ZN (n_7187), .A (n_7197), .B1 (n_7189), .B2 (n_7188));
NAND3_X1 i_7250 (.ZN (n_7186), .A1 (n_7189), .A2 (n_7188), .A3 (n_7197));
INV_X1 i_7249 (.ZN (n_7185), .A (n_7186));
NOR2_X1 i_7248 (.ZN (n_7184), .A1 (n_7185), .A2 (n_7187));
NAND2_X1 i_7247 (.ZN (n_7183), .A1 (B_imm[27]), .A2 (A_imm[17]));
OAI22_X1 i_7246 (.ZN (n_7182), .A1 (n_8525), .A2 (n_8794), .B1 (n_8993), .B2 (n_8956));
NAND4_X1 i_7245 (.ZN (n_7181), .A1 (B_imm[19]), .A2 (B_imm[26]), .A3 (A_imm[25]), .A4 (A_imm[18]));
NAND2_X1 i_7244 (.ZN (n_7180), .A1 (n_7182), .A2 (n_7181));
XNOR2_X1 i_7243 (.ZN (n_7179), .A (n_7180), .B (n_7183));
NAND2_X1 i_7242 (.ZN (n_7178), .A1 (n_7428), .A2 (n_7445));
NAND2_X1 i_7241 (.ZN (n_7177), .A1 (B_imm[25]), .A2 (A_imm[19]));
OAI22_X1 i_7240 (.ZN (n_7176), .A1 (n_8958), .A2 (n_8906), .B1 (n_8957), .B2 (n_8907));
NAND4_X1 i_7239 (.ZN (n_7175), .A1 (B_imm[22]), .A2 (B_imm[21]), .A3 (A_imm[23]), .A4 (A_imm[22]));
NAND2_X1 i_7238 (.ZN (n_7174), .A1 (n_7176), .A2 (n_7175));
XNOR2_X1 i_7237 (.ZN (n_7173), .A (n_7174), .B (n_7177));
INV_X1 i_7236 (.ZN (n_7172), .A (n_7173));
NAND3_X1 i_7235 (.ZN (n_7171), .A1 (n_7172), .A2 (n_7431), .A3 (n_7178));
NAND2_X1 i_7234 (.ZN (n_7170), .A1 (n_7178), .A2 (n_7431));
NAND2_X1 i_7233 (.ZN (n_7169), .A1 (n_7170), .A2 (n_7173));
NAND3_X1 i_7232 (.ZN (n_7168), .A1 (n_7171), .A2 (n_7169), .A3 (n_7179));
INV_X1 i_7231 (.ZN (n_7167), .A (n_7179));
INV_X1 i_7230 (.ZN (n_7166), .A (n_7171));
INV_X1 i_7229 (.ZN (n_7165), .A (n_7169));
OAI21_X1 i_7228 (.ZN (n_7164), .A (n_7167), .B1 (n_7165), .B2 (n_7166));
NAND2_X1 i_7227 (.ZN (n_7163), .A1 (n_7164), .A2 (n_7168));
NAND2_X1 i_7226 (.ZN (n_7162), .A1 (n_7163), .A2 (n_7184));
OAI211_X1 i_7225 (.ZN (n_7161), .A (n_7164), .B (n_7168), .C1 (n_7187), .C2 (n_7185));
NAND2_X1 i_7224 (.ZN (n_7160), .A1 (n_7271), .A2 (n_7262));
NAND4_X1 i_7223 (.ZN (n_7159), .A1 (n_7162), .A2 (n_7161), .A3 (n_7160), .A4 (n_7273));
NAND2_X1 i_7222 (.ZN (n_7158), .A1 (n_7161), .A2 (n_7162));
NAND2_X1 i_7221 (.ZN (n_7157), .A1 (n_7160), .A2 (n_7273));
NAND2_X1 i_7220 (.ZN (n_7156), .A1 (n_7158), .A2 (n_7157));
NAND2_X1 i_7219 (.ZN (n_7155), .A1 (n_7156), .A2 (n_7159));
NAND2_X1 i_7218 (.ZN (n_7154), .A1 (n_7326), .A2 (n_7343));
NAND2_X1 i_7217 (.ZN (n_7153), .A1 (n_7154), .A2 (n_7328));
NAND2_X1 i_7216 (.ZN (n_7152), .A1 (n_7332), .A2 (n_7334));
NAND2_X1 i_7215 (.ZN (n_7151), .A1 (n_7152), .A2 (n_7333));
INV_X1 i_7214 (.ZN (n_7150), .A (n_7151));
OAI22_X1 i_7213 (.ZN (n_7149), .A1 (n_9038), .A2 (n_8927), .B1 (n_9004), .B2 (n_8971));
NAND4_X1 i_7212 (.ZN (n_7148), .A1 (B_imm[31]), .A2 (B_imm[30]), .A3 (A_imm[14]), .A4 (A_imm[13]));
NAND2_X1 i_7211 (.ZN (n_7147), .A1 (n_7149), .A2 (n_7148));
XNOR2_X1 i_7210 (.ZN (n_7146), .A (n_7147), .B (n_7150));
NAND2_X1 i_7209 (.ZN (n_7145), .A1 (B_imm[21]), .A2 (A_imm[22]));
INV_X1 i_7208 (.ZN (n_7144), .A (n_7145));
OAI22_X1 i_7207 (.ZN (n_7143), .A1 (n_8821), .A2 (n_8893), .B1 (n_9037), .B2 (n_8795));
INV_X1 i_7206 (.ZN (n_7142), .A (n_7143));
NAND4_X1 i_7205 (.ZN (n_7141), .A1 (B_imm[23]), .A2 (A_imm[31]), .A3 (B_imm[12]), .A4 (A_imm[20]));
INV_X1 i_7204 (.ZN (n_7140), .A (n_7141));
OAI21_X1 i_7203 (.ZN (n_7139), .A (n_7144), .B1 (n_7142), .B2 (n_7140));
NAND3_X1 i_7202 (.ZN (n_7138), .A1 (n_7143), .A2 (n_7145), .A3 (n_7141));
NAND2_X1 i_7201 (.ZN (n_7137), .A1 (n_7139), .A2 (n_7138));
NAND2_X1 i_7200 (.ZN (n_7136), .A1 (B_imm[24]), .A2 (A_imm[19]));
INV_X1 i_7199 (.ZN (n_7135), .A (n_7136));
OAI22_X1 i_7198 (.ZN (n_7134), .A1 (n_8423), .A2 (n_8794), .B1 (n_8972), .B2 (n_8909));
INV_X1 i_7197 (.ZN (n_7133), .A (n_7134));
NAND4_X1 i_7196 (.ZN (n_7132), .A1 (B_imm[18]), .A2 (A_imm[26]), .A3 (A_imm[25]), .A4 (B_imm[17]));
INV_X1 i_7195 (.ZN (n_7131), .A (n_7132));
OAI21_X1 i_7194 (.ZN (n_7130), .A (n_7135), .B1 (n_7133), .B2 (n_7131));
NAND3_X1 i_7193 (.ZN (n_7129), .A1 (n_7134), .A2 (n_7136), .A3 (n_7132));
NAND2_X1 i_7192 (.ZN (n_7128), .A1 (n_7130), .A2 (n_7129));
NAND2_X1 i_7191 (.ZN (n_7127), .A1 (n_7137), .A2 (n_7128));
NAND4_X1 i_7190 (.ZN (n_7126), .A1 (n_7139), .A2 (n_7130), .A3 (n_7138), .A4 (n_7129));
INV_X1 i_7189 (.ZN (n_7125), .A (n_7126));
NAND2_X1 i_7188 (.ZN (n_7124), .A1 (B_imm[20]), .A2 (A_imm[23]));
OAI22_X1 i_7187 (.ZN (n_7123), .A1 (n_8974), .A2 (n_8956), .B1 (n_8958), .B2 (n_8859));
NAND4_X1 i_7186 (.ZN (n_7122), .A1 (B_imm[25]), .A2 (B_imm[22]), .A3 (A_imm[21]), .A4 (A_imm[18]));
NAND2_X1 i_7185 (.ZN (n_7121), .A1 (n_7123), .A2 (n_7122));
XNOR2_X1 i_7184 (.ZN (n_7120), .A (n_7121), .B (n_7124));
OAI21_X1 i_7183 (.ZN (n_7119), .A (n_7127), .B1 (n_7120), .B2 (n_7125));
NAND2_X1 i_7182 (.ZN (n_7118), .A1 (n_7146), .A2 (n_7119));
INV_X1 i_7181 (.ZN (n_7117), .A (n_7146));
INV_X1 i_7180 (.ZN (n_7116), .A (n_7119));
NAND2_X1 i_7179 (.ZN (n_7115), .A1 (n_7117), .A2 (n_7116));
NAND3_X1 i_7178 (.ZN (n_7114), .A1 (n_7115), .A2 (n_7153), .A3 (n_7118));
NAND2_X1 i_7177 (.ZN (n_7113), .A1 (n_7115), .A2 (n_7118));
NAND3_X1 i_7176 (.ZN (n_7112), .A1 (n_7113), .A2 (n_7328), .A3 (n_7154));
INV_X1 i_7175 (.ZN (n_7111), .A (n_7124));
INV_X1 i_7174 (.ZN (n_7110), .A (n_7122));
OAI21_X1 i_7173 (.ZN (n_7109), .A (n_7123), .B1 (n_7111), .B2 (n_7110));
INV_X1 i_7172 (.ZN (n_7108), .A (n_7109));
OAI21_X1 i_7171 (.ZN (n_7107), .A (n_7143), .B1 (n_7144), .B2 (n_7140));
OAI21_X1 i_7170 (.ZN (n_7106), .A (n_7107), .B1 (n_8909), .B2 (n_7912));
INV_X1 i_7169 (.ZN (n_7105), .A (n_7107));
NAND3_X1 i_7168 (.ZN (n_7104), .A1 (n_7105), .A2 (B_imm[17]), .A3 (A_imm[27]));
NAND2_X1 i_7167 (.ZN (n_7103), .A1 (n_7104), .A2 (n_7106));
NAND2_X1 i_7166 (.ZN (n_7102), .A1 (n_7103), .A2 (n_7108));
NAND3_X1 i_7165 (.ZN (n_7101), .A1 (n_7104), .A2 (n_7109), .A3 (n_7106));
OAI21_X1 i_7164 (.ZN (n_7100), .A (n_7134), .B1 (n_7131), .B2 (n_7135));
INV_X1 i_7163 (.ZN (n_7099), .A (n_7100));
OAI22_X1 i_7162 (.ZN (n_7098), .A1 (n_9020), .A2 (n_8908), .B1 (n_9006), .B2 (n_8946));
NAND4_X1 i_7161 (.ZN (n_7097), .A1 (A_imm[28]), .A2 (B_imm[29]), .A3 (B_imm[16]), .A4 (A_imm[15]));
NAND2_X1 i_7160 (.ZN (n_7096), .A1 (n_7098), .A2 (n_7097));
XNOR2_X1 i_7159 (.ZN (n_7095), .A (n_7096), .B (n_7099));
INV_X1 i_7158 (.ZN (n_7094), .A (n_7264));
OAI21_X1 i_7157 (.ZN (n_7093), .A (n_7266), .B1 (n_7094), .B2 (n_7269));
INV_X1 i_7156 (.ZN (n_7092), .A (n_7093));
NAND2_X1 i_7155 (.ZN (n_7091), .A1 (n_7092), .A2 (n_7095));
INV_X1 i_7154 (.ZN (n_7090), .A (n_7095));
NAND2_X1 i_7153 (.ZN (n_7089), .A1 (n_7090), .A2 (n_7093));
NAND4_X1 i_7152 (.ZN (n_7088), .A1 (n_7089), .A2 (n_7091), .A3 (n_7102), .A4 (n_7101));
NAND2_X1 i_7151 (.ZN (n_7087), .A1 (n_7102), .A2 (n_7101));
NAND2_X1 i_7150 (.ZN (n_7086), .A1 (n_7089), .A2 (n_7091));
NAND2_X1 i_7149 (.ZN (n_7085), .A1 (n_7086), .A2 (n_7087));
NAND2_X1 i_7148 (.ZN (n_7084), .A1 (n_7085), .A2 (n_7088));
NAND3_X1 i_7147 (.ZN (n_7083), .A1 (n_7112), .A2 (n_7084), .A3 (n_7114));
NAND2_X1 i_7146 (.ZN (n_7082), .A1 (n_7112), .A2 (n_7114));
INV_X1 i_7145 (.ZN (n_7081), .A (n_7084));
NAND2_X1 i_7144 (.ZN (n_7080), .A1 (n_7082), .A2 (n_7081));
INV_X1 i_7143 (.ZN (n_7079), .A (n_7127));
OAI21_X1 i_7142 (.ZN (n_7078), .A (n_7120), .B1 (n_7079), .B2 (n_7125));
INV_X1 i_7141 (.ZN (n_7077), .A (n_7120));
NAND3_X1 i_7140 (.ZN (n_7076), .A1 (n_7077), .A2 (n_7127), .A3 (n_7126));
INV_X1 i_7139 (.ZN (n_7075), .A (n_7775));
OAI21_X1 i_7138 (.ZN (n_7074), .A (n_7777), .B1 (n_7075), .B2 (n_7780));
INV_X1 i_7137 (.ZN (n_7073), .A (n_7074));
INV_X1 i_7136 (.ZN (n_7072), .A (n_7337));
NAND2_X1 i_7135 (.ZN (n_7071), .A1 (n_7336), .A2 (n_7338));
NAND2_X1 i_7134 (.ZN (n_7070), .A1 (n_7071), .A2 (n_7072));
NAND3_X1 i_7133 (.ZN (n_7069), .A1 (n_7338), .A2 (n_7336), .A3 (n_7337));
NAND2_X1 i_7132 (.ZN (n_7068), .A1 (n_7070), .A2 (n_7069));
NAND2_X1 i_7131 (.ZN (n_7067), .A1 (n_7073), .A2 (n_7068));
NAND3_X1 i_7130 (.ZN (n_7066), .A1 (n_7074), .A2 (n_7069), .A3 (n_7070));
AOI21_X1 i_7129 (.ZN (n_7065), .A (n_7908), .B1 (n_7902), .B2 (n_7911));
INV_X1 i_7128 (.ZN (n_7064), .A (n_7065));
NAND2_X1 i_7127 (.ZN (n_7063), .A1 (n_7066), .A2 (n_7064));
NAND2_X1 i_7126 (.ZN (n_7062), .A1 (n_7063), .A2 (n_7067));
NAND3_X1 i_7125 (.ZN (n_7061), .A1 (n_7062), .A2 (n_7078), .A3 (n_7076));
NAND2_X1 i_7124 (.ZN (n_7060), .A1 (n_7078), .A2 (n_7076));
NAND3_X1 i_7123 (.ZN (n_7059), .A1 (n_7063), .A2 (n_7060), .A3 (n_7067));
NAND3_X1 i_7122 (.ZN (n_7058), .A1 (n_7377), .A2 (n_7379), .A3 (n_7375));
INV_X1 i_7121 (.ZN (n_7057), .A (n_7379));
OAI21_X1 i_7120 (.ZN (n_7056), .A (n_7374), .B1 (n_7378), .B2 (n_7057));
NAND2_X1 i_7119 (.ZN (n_7055), .A1 (n_7056), .A2 (n_7058));
NAND2_X1 i_7118 (.ZN (n_7054), .A1 (n_7055), .A2 (n_7059));
NAND2_X1 i_7117 (.ZN (n_7053), .A1 (n_7054), .A2 (n_7061));
NAND3_X1 i_7116 (.ZN (n_7052), .A1 (n_7080), .A2 (n_7083), .A3 (n_7053));
NAND2_X1 i_7115 (.ZN (n_7051), .A1 (n_7080), .A2 (n_7083));
INV_X1 i_7114 (.ZN (n_7050), .A (n_7053));
NAND2_X1 i_7113 (.ZN (n_7049), .A1 (n_7051), .A2 (n_7050));
NAND3_X1 i_7112 (.ZN (n_7048), .A1 (n_7049), .A2 (n_7155), .A3 (n_7052));
AOI21_X1 i_7111 (.ZN (n_7047), .A (n_7155), .B1 (n_7052), .B2 (n_7049));
INV_X1 i_7110 (.ZN (n_7046), .A (n_7047));
NAND3_X1 i_7109 (.ZN (n_7045), .A1 (n_7061), .A2 (n_7059), .A3 (n_7055));
NAND2_X1 i_7108 (.ZN (n_7044), .A1 (n_7061), .A2 (n_7059));
NAND3_X1 i_7107 (.ZN (n_7043), .A1 (n_7044), .A2 (n_7058), .A3 (n_7056));
NAND2_X1 i_7106 (.ZN (n_7042), .A1 (n_7043), .A2 (n_7045));
INV_X1 i_7105 (.ZN (n_7041), .A (n_7042));
INV_X1 i_7104 (.ZN (n_7040), .A (n_7349));
NAND3_X1 i_7103 (.ZN (n_7039), .A1 (n_7358), .A2 (n_7357), .A3 (n_7040));
INV_X1 i_7102 (.ZN (n_7038), .A (n_7039));
AOI21_X1 i_7101 (.ZN (n_7037), .A (n_7040), .B1 (n_7357), .B2 (n_7358));
INV_X1 i_7100 (.ZN (n_7036), .A (n_7278));
NAND2_X1 i_7099 (.ZN (n_7035), .A1 (n_7279), .A2 (n_7276));
NAND2_X1 i_7098 (.ZN (n_7034), .A1 (n_7035), .A2 (n_7036));
NAND3_X1 i_7097 (.ZN (n_7033), .A1 (n_7279), .A2 (n_7276), .A3 (n_7278));
NAND2_X1 i_7096 (.ZN (n_7032), .A1 (n_7034), .A2 (n_7033));
OAI21_X1 i_7095 (.ZN (n_7031), .A (n_7032), .B1 (n_7038), .B2 (n_7037));
INV_X1 i_7094 (.ZN (n_7030), .A (n_7037));
NAND4_X1 i_7093 (.ZN (n_7029), .A1 (n_7030), .A2 (n_7039), .A3 (n_7034), .A4 (n_7033));
AOI21_X1 i_7092 (.ZN (n_7028), .A (n_7064), .B1 (n_7066), .B2 (n_7067));
NAND3_X1 i_7091 (.ZN (n_7027), .A1 (n_7067), .A2 (n_7066), .A3 (n_7064));
INV_X1 i_7090 (.ZN (n_7026), .A (n_7027));
NOR2_X1 i_7089 (.ZN (n_7025), .A1 (n_7026), .A2 (n_7028));
NAND2_X1 i_7088 (.ZN (n_7024), .A1 (n_7029), .A2 (n_7025));
NAND2_X1 i_7087 (.ZN (n_7023), .A1 (n_7024), .A2 (n_7031));
NAND2_X1 i_7086 (.ZN (n_7022), .A1 (n_7023), .A2 (n_7041));
NAND3_X1 i_7085 (.ZN (n_7021), .A1 (n_7042), .A2 (n_7031), .A3 (n_7024));
AOI21_X1 i_7084 (.ZN (n_7020), .A (n_7308), .B1 (n_7314), .B2 (n_7315));
NAND3_X1 i_7083 (.ZN (n_7019), .A1 (n_7315), .A2 (n_7308), .A3 (n_7314));
INV_X1 i_7082 (.ZN (n_7018), .A (n_7019));
NAND3_X1 i_7081 (.ZN (n_7017), .A1 (n_7841), .A2 (n_7827), .A3 (n_7824));
NAND2_X1 i_7080 (.ZN (n_7016), .A1 (n_7017), .A2 (n_7839));
OAI21_X1 i_7079 (.ZN (n_7015), .A (n_7016), .B1 (n_7018), .B2 (n_7020));
INV_X1 i_7078 (.ZN (n_7014), .A (n_7020));
NAND4_X1 i_7077 (.ZN (n_7013), .A1 (n_7014), .A2 (n_7839), .A3 (n_7019), .A4 (n_7017));
INV_X1 i_7076 (.ZN (n_7012), .A (n_8867));
OAI21_X1 i_7075 (.ZN (n_7011), .A (n_8865), .B1 (n_7012), .B2 (n_8841));
INV_X1 i_7074 (.ZN (n_7010), .A (n_7011));
NAND2_X1 i_7073 (.ZN (n_7009), .A1 (n_7013), .A2 (n_7010));
NAND2_X1 i_7072 (.ZN (n_7008), .A1 (n_7009), .A2 (n_7015));
INV_X1 i_7071 (.ZN (n_7007), .A (n_7008));
NAND2_X1 i_7070 (.ZN (n_7006), .A1 (n_7007), .A2 (n_7021));
NAND2_X2 i_7069 (.ZN (n_7005), .A1 (n_7006), .A2 (n_7022));
NAND3_X1 i_7068 (.ZN (n_7004), .A1 (n_7005), .A2 (n_7046), .A3 (n_7048));
INV_X1 i_7067 (.ZN (n_7003), .A (n_7048));
OAI211_X1 i_7066 (.ZN (n_7002), .A (n_7022), .B (n_7006), .C1 (n_7003), .C2 (n_7047));
NAND2_X1 i_7065 (.ZN (n_7001), .A1 (n_7002), .A2 (n_7004));
NAND3_X1 i_7064 (.ZN (n_7000), .A1 (n_7200), .A2 (n_7199), .A3 (n_7001));
INV_X1 i_7063 (.ZN (n_6999), .A (n_7199));
INV_X1 i_7062 (.ZN (n_6998), .A (n_7001));
OAI21_X1 i_7061 (.ZN (n_6997), .A (n_6998), .B1 (n_6999), .B2 (n_7201));
NAND3_X1 i_7060 (.ZN (n_6996), .A1 (n_7022), .A2 (n_7008), .A3 (n_7021));
NAND2_X1 i_7059 (.ZN (n_6995), .A1 (n_7022), .A2 (n_7021));
NAND2_X1 i_7058 (.ZN (n_6994), .A1 (n_6995), .A2 (n_7007));
NAND3_X1 i_7057 (.ZN (n_6993), .A1 (n_7015), .A2 (n_7013), .A3 (n_7010));
INV_X1 i_7056 (.ZN (n_6992), .A (n_6993));
AOI21_X1 i_7055 (.ZN (n_6991), .A (n_7010), .B1 (n_7013), .B2 (n_7015));
NAND3_X1 i_7054 (.ZN (n_6990), .A1 (n_7029), .A2 (n_7031), .A3 (n_7025));
INV_X1 i_7053 (.ZN (n_6989), .A (n_6990));
AOI21_X1 i_7052 (.ZN (n_6988), .A (n_7025), .B1 (n_7031), .B2 (n_7029));
NOR2_X1 i_7051 (.ZN (n_6987), .A1 (n_6989), .A2 (n_6988));
OAI21_X2 i_7050 (.ZN (n_6986), .A (n_6987), .B1 (n_6992), .B2 (n_6991));
NAND2_X1 i_7049 (.ZN (n_6985), .A1 (n_7013), .A2 (n_7015));
NAND2_X1 i_7048 (.ZN (n_6984), .A1 (n_6985), .A2 (n_7011));
INV_X1 i_7047 (.ZN (n_6983), .A (n_6988));
NAND2_X1 i_7046 (.ZN (n_6982), .A1 (n_6983), .A2 (n_6990));
NAND3_X1 i_7045 (.ZN (n_6981), .A1 (n_6982), .A2 (n_6984), .A3 (n_6993));
INV_X1 i_7044 (.ZN (n_6980), .A (n_8404));
OAI21_X1 i_7043 (.ZN (n_6979), .A (n_8658), .B1 (n_6980), .B2 (n_8323));
NAND2_X1 i_7042 (.ZN (n_6978), .A1 (n_6979), .A2 (n_8656));
NAND2_X2 i_7041 (.ZN (n_6977), .A1 (n_6978), .A2 (n_6981));
AOI22_X2 i_7040 (.ZN (n_6976), .A1 (n_6977), .A2 (n_6986), .B1 (n_6996), .B2 (n_6994));
INV_X1 i_7039 (.ZN (n_6975), .A (n_6976));
NAND2_X1 i_7038 (.ZN (n_6974), .A1 (n_6994), .A2 (n_6996));
INV_X1 i_7037 (.ZN (n_6973), .A (n_6974));
NAND3_X1 i_7036 (.ZN (n_6972), .A1 (n_6977), .A2 (n_6973), .A3 (n_6986));
NAND3_X1 i_7035 (.ZN (n_6971), .A1 (n_7216), .A2 (n_7219), .A3 (n_7203));
INV_X1 i_7034 (.ZN (n_6970), .A (n_7203));
NAND2_X1 i_7033 (.ZN (n_6969), .A1 (n_7216), .A2 (n_7219));
NAND2_X1 i_7032 (.ZN (n_6968), .A1 (n_6969), .A2 (n_6970));
NAND2_X1 i_7031 (.ZN (n_6967), .A1 (n_6968), .A2 (n_6971));
INV_X1 i_7030 (.ZN (n_6966), .A (n_6967));
NAND2_X1 i_7029 (.ZN (n_6965), .A1 (n_6966), .A2 (n_6972));
NAND4_X2 i_7028 (.ZN (n_6964), .A1 (n_6997), .A2 (n_7000), .A3 (n_6975), .A4 (n_6965));
NAND3_X1 i_7027 (.ZN (n_6963), .A1 (n_6975), .A2 (n_6972), .A3 (n_6967));
INV_X1 i_7026 (.ZN (n_6962), .A (n_6972));
OAI21_X2 i_7025 (.ZN (n_6961), .A (n_6966), .B1 (n_6962), .B2 (n_6976));
NAND3_X1 i_7024 (.ZN (n_6960), .A1 (n_7208), .A2 (n_7207), .A3 (n_7205));
INV_X1 i_7023 (.ZN (n_6959), .A (n_7205));
NAND2_X1 i_7022 (.ZN (n_6958), .A1 (n_7208), .A2 (n_7207));
NAND2_X1 i_7021 (.ZN (n_6957), .A1 (n_6958), .A2 (n_6959));
NAND2_X1 i_7020 (.ZN (n_6956), .A1 (n_7741), .A2 (n_7761));
NAND2_X1 i_7019 (.ZN (n_6955), .A1 (n_6956), .A2 (n_7759));
NAND3_X1 i_7018 (.ZN (n_6954), .A1 (n_6955), .A2 (n_6960), .A3 (n_6957));
NAND2_X1 i_7017 (.ZN (n_6953), .A1 (n_6957), .A2 (n_6960));
NAND3_X1 i_7016 (.ZN (n_6952), .A1 (n_6953), .A2 (n_6956), .A3 (n_7759));
INV_X1 i_7015 (.ZN (n_6951), .A (n_6952));
NAND3_X1 i_7014 (.ZN (n_6950), .A1 (n_6978), .A2 (n_6986), .A3 (n_6981));
INV_X1 i_7013 (.ZN (n_6949), .A (n_6978));
NAND2_X1 i_7012 (.ZN (n_6948), .A1 (n_6986), .A2 (n_6981));
NAND2_X1 i_7011 (.ZN (n_6947), .A1 (n_6948), .A2 (n_6949));
NAND2_X1 i_7010 (.ZN (n_6946), .A1 (n_6947), .A2 (n_6950));
OAI21_X1 i_7009 (.ZN (n_6945), .A (n_6954), .B1 (n_6951), .B2 (n_6946));
INV_X1 i_7008 (.ZN (n_6944), .A (n_6945));
NAND3_X2 i_7007 (.ZN (n_6943), .A1 (n_6944), .A2 (n_6961), .A3 (n_6963));
NAND3_X1 i_7006 (.ZN (n_6942), .A1 (n_6954), .A2 (n_6952), .A3 (n_6946));
INV_X1 i_7005 (.ZN (n_6941), .A (n_6946));
NAND2_X1 i_7004 (.ZN (n_6940), .A1 (n_6954), .A2 (n_6952));
NAND2_X1 i_7003 (.ZN (n_6939), .A1 (n_6940), .A2 (n_6941));
OAI21_X1 i_7002 (.ZN (n_6938), .A (n_7914), .B1 (n_7736), .B2 (n_7734));
INV_X1 i_7001 (.ZN (n_6937), .A (n_6938));
NAND3_X2 i_7000 (.ZN (n_6936), .A1 (n_6937), .A2 (n_6939), .A3 (n_6942));
NAND4_X1 i_6999 (.ZN (n_6935), .A1 (n_7465), .A2 (n_6936), .A3 (n_6964), .A4 (n_6943));
INV_X2 i_6998 (.ZN (n_6934), .A (n_6935));
NAND3_X1 i_6997 (.ZN (n_6933), .A1 (n_7586), .A2 (n_7643), .A3 (n_7638));
INV_X1 i_6996 (.ZN (n_6932), .A (n_7586));
NAND2_X1 i_6995 (.ZN (n_6931), .A1 (n_7643), .A2 (n_7638));
NAND2_X1 i_6994 (.ZN (n_6930), .A1 (n_6931), .A2 (n_6932));
NAND2_X1 i_6993 (.ZN (n_6929), .A1 (n_6930), .A2 (n_6933));
NAND3_X1 i_6992 (.ZN (n_6928), .A1 (n_8130), .A2 (n_8082), .A3 (n_8129));
INV_X1 i_6991 (.ZN (n_6927), .A (n_8082));
NAND2_X1 i_6990 (.ZN (n_6926), .A1 (n_8130), .A2 (n_8129));
NAND2_X1 i_6989 (.ZN (n_6925), .A1 (n_6926), .A2 (n_6927));
NAND3_X1 i_6988 (.ZN (n_6924), .A1 (n_7647), .A2 (n_7656), .A3 (n_7654));
NAND2_X1 i_6987 (.ZN (n_6923), .A1 (n_7656), .A2 (n_7654));
NAND2_X1 i_6986 (.ZN (n_6922), .A1 (n_6923), .A2 (n_7648));
NAND2_X1 i_6985 (.ZN (n_6921), .A1 (n_6922), .A2 (n_6924));
NAND2_X1 i_6984 (.ZN (n_6920), .A1 (A_imm[30]), .A2 (B_imm[5]));
AOI21_X1 i_6983 (.ZN (n_6919), .A (n_6920), .B1 (n_7699), .B2 (n_7698));
NAND3_X1 i_6982 (.ZN (n_6918), .A1 (n_7699), .A2 (n_7698), .A3 (n_6920));
INV_X1 i_6981 (.ZN (n_6917), .A (n_6918));
OAI21_X2 i_6980 (.ZN (n_6916), .A (n_6921), .B1 (n_6919), .B2 (n_6917));
NOR2_X1 i_6979 (.ZN (n_6915), .A1 (n_6917), .A2 (n_6919));
NAND3_X2 i_6978 (.ZN (n_6914), .A1 (n_6922), .A2 (n_6915), .A3 (n_6924));
NAND2_X1 i_6977 (.ZN (n_6913), .A1 (n_7679), .A2 (n_7672));
NAND2_X1 i_6976 (.ZN (n_6912), .A1 (n_6913), .A2 (n_7673));
NAND3_X1 i_6975 (.ZN (n_6911), .A1 (n_7679), .A2 (n_7672), .A3 (n_7674));
NAND2_X1 i_6974 (.ZN (n_6910), .A1 (n_8092), .A2 (n_8089));
NAND2_X1 i_6973 (.ZN (n_6909), .A1 (n_6910), .A2 (n_8090));
NAND3_X1 i_6972 (.ZN (n_6908), .A1 (n_8092), .A2 (n_8091), .A3 (n_8089));
NAND4_X1 i_6971 (.ZN (n_6907), .A1 (n_6912), .A2 (n_6909), .A3 (n_6911), .A4 (n_6908));
NAND2_X1 i_6970 (.ZN (n_6906), .A1 (n_6912), .A2 (n_6911));
NAND2_X1 i_6969 (.ZN (n_6905), .A1 (n_6909), .A2 (n_6908));
NAND2_X1 i_6968 (.ZN (n_6904), .A1 (n_6906), .A2 (n_6905));
AOI21_X1 i_6967 (.ZN (n_6903), .A (n_7688), .B1 (n_7689), .B2 (n_7687));
NAND3_X1 i_6966 (.ZN (n_6902), .A1 (n_7689), .A2 (n_7688), .A3 (n_7687));
INV_X1 i_6965 (.ZN (n_6901), .A (n_6902));
NOR2_X1 i_6964 (.ZN (n_6900), .A1 (n_6901), .A2 (n_6903));
NAND2_X1 i_6963 (.ZN (n_6899), .A1 (n_6904), .A2 (n_6900));
NAND2_X1 i_6962 (.ZN (n_6898), .A1 (B_imm[29]), .A2 (A_imm[3]));
NAND2_X1 i_6961 (.ZN (n_6897), .A1 (A_imm[24]), .A2 (B_imm[7]));
OAI21_X1 i_6960 (.ZN (n_6896), .A (n_6897), .B1 (n_8907), .B2 (n_8947));
NAND2_X1 i_6959 (.ZN (n_6895), .A1 (B_imm[12]), .A2 (A_imm[19]));
NAND4_X1 i_6958 (.ZN (n_6894), .A1 (A_imm[23]), .A2 (A_imm[24]), .A3 (B_imm[8]), .A4 (B_imm[7]));
NAND2_X1 i_6957 (.ZN (n_6893), .A1 (n_6894), .A2 (n_6895));
NAND2_X1 i_6956 (.ZN (n_6892), .A1 (n_6893), .A2 (n_6896));
NAND2_X1 i_6955 (.ZN (n_6891), .A1 (n_6892), .A2 (n_6898));
NAND2_X1 i_6954 (.ZN (n_6890), .A1 (A_imm[28]), .A2 (B_imm[4]));
NAND4_X1 i_6953 (.ZN (n_6889), .A1 (n_6893), .A2 (B_imm[29]), .A3 (A_imm[3]), .A4 (n_6896));
NAND2_X1 i_6952 (.ZN (n_6888), .A1 (n_6889), .A2 (n_6890));
NAND2_X1 i_6951 (.ZN (n_6887), .A1 (n_8126), .A2 (n_8123));
NAND2_X1 i_6950 (.ZN (n_6886), .A1 (n_6887), .A2 (n_8124));
NAND3_X1 i_6949 (.ZN (n_6885), .A1 (n_8126), .A2 (n_8125), .A3 (n_8123));
NAND2_X1 i_6948 (.ZN (n_6884), .A1 (n_6886), .A2 (n_6885));
NAND3_X1 i_6947 (.ZN (n_6883), .A1 (n_6884), .A2 (n_6888), .A3 (n_6891));
INV_X1 i_6946 (.ZN (n_6882), .A (n_6883));
INV_X1 i_6945 (.ZN (n_6881), .A (n_6890));
INV_X1 i_6944 (.ZN (n_6880), .A (n_6889));
OAI21_X1 i_6943 (.ZN (n_6879), .A (n_6891), .B1 (n_6880), .B2 (n_6881));
INV_X1 i_6942 (.ZN (n_6878), .A (n_6884));
NAND2_X1 i_6941 (.ZN (n_6877), .A1 (n_8101), .A2 (n_8099));
NAND3_X1 i_6940 (.ZN (n_6876), .A1 (n_6877), .A2 (B_imm[15]), .A3 (A_imm[18]));
NAND3_X1 i_6939 (.ZN (n_6875), .A1 (n_8101), .A2 (n_8100), .A3 (n_8099));
AOI22_X1 i_6938 (.ZN (n_6874), .A1 (n_6879), .A2 (n_6878), .B1 (n_6876), .B2 (n_6875));
OAI211_X1 i_6937 (.ZN (n_6873), .A (n_6899), .B (n_6907), .C1 (n_6874), .C2 (n_6882));
NAND2_X1 i_6936 (.ZN (n_6872), .A1 (n_6899), .A2 (n_6907));
NOR2_X1 i_6935 (.ZN (n_6871), .A1 (n_6874), .A2 (n_6882));
NAND2_X1 i_6934 (.ZN (n_6870), .A1 (n_6872), .A2 (n_6871));
NAND2_X1 i_6933 (.ZN (n_6869), .A1 (n_7684), .A2 (n_7683));
NAND2_X1 i_6932 (.ZN (n_6868), .A1 (n_6869), .A2 (n_7669));
NAND3_X1 i_6931 (.ZN (n_6867), .A1 (n_7684), .A2 (n_7683), .A3 (n_7670));
NAND2_X1 i_6930 (.ZN (n_6866), .A1 (n_6868), .A2 (n_6867));
NAND2_X1 i_6929 (.ZN (n_6865), .A1 (n_6870), .A2 (n_6866));
NAND2_X1 i_6928 (.ZN (n_6864), .A1 (n_6865), .A2 (n_6873));
NAND2_X1 i_6927 (.ZN (n_6863), .A1 (n_6864), .A2 (n_6914));
NAND2_X1 i_6926 (.ZN (n_6862), .A1 (n_6863), .A2 (n_6916));
NAND3_X1 i_6925 (.ZN (n_6861), .A1 (n_6862), .A2 (n_6928), .A3 (n_6925));
NAND2_X1 i_6924 (.ZN (n_6860), .A1 (n_6925), .A2 (n_6928));
NAND3_X1 i_6923 (.ZN (n_6859), .A1 (n_6863), .A2 (n_6916), .A3 (n_6860));
NAND2_X1 i_6922 (.ZN (n_6858), .A1 (n_7646), .A2 (n_7656));
NAND3_X1 i_6921 (.ZN (n_6857), .A1 (n_6858), .A2 (n_7695), .A3 (n_7693));
NAND2_X1 i_6920 (.ZN (n_6856), .A1 (n_7695), .A2 (n_7693));
NAND3_X1 i_6919 (.ZN (n_6855), .A1 (n_6856), .A2 (n_7656), .A3 (n_7646));
NAND2_X1 i_6918 (.ZN (n_6854), .A1 (n_6855), .A2 (n_6857));
NAND2_X1 i_6917 (.ZN (n_6853), .A1 (n_6859), .A2 (n_6854));
NAND3_X1 i_6916 (.ZN (n_6852), .A1 (n_6929), .A2 (n_6861), .A3 (n_6853));
INV_X1 i_6915 (.ZN (n_6851), .A (n_6929));
NAND2_X1 i_6914 (.ZN (n_6850), .A1 (n_6853), .A2 (n_6861));
NAND2_X1 i_6913 (.ZN (n_6849), .A1 (n_6850), .A2 (n_6851));
NAND3_X1 i_6912 (.ZN (n_6848), .A1 (n_7594), .A2 (n_7593), .A3 (n_7588));
INV_X1 i_6911 (.ZN (n_6847), .A (n_7593));
INV_X1 i_6910 (.ZN (n_6846), .A (n_7588));
OAI21_X1 i_6909 (.ZN (n_6845), .A (n_6846), .B1 (n_6847), .B2 (n_7595));
NAND2_X1 i_6908 (.ZN (n_6844), .A1 (n_6845), .A2 (n_6848));
INV_X1 i_6907 (.ZN (n_6843), .A (n_6844));
NAND2_X1 i_6906 (.ZN (n_6842), .A1 (n_7605), .A2 (n_7614));
NAND2_X1 i_6905 (.ZN (n_6841), .A1 (n_7621), .A2 (n_7624));
NAND2_X1 i_6904 (.ZN (n_6840), .A1 (n_6841), .A2 (n_6842));
NAND4_X1 i_6903 (.ZN (n_6839), .A1 (n_7621), .A2 (n_7624), .A3 (n_7614), .A4 (n_7605));
NAND2_X1 i_6902 (.ZN (n_6838), .A1 (n_6840), .A2 (n_6839));
NAND2_X1 i_6901 (.ZN (n_6837), .A1 (A_imm[30]), .A2 (B_imm[3]));
INV_X2 i_6900 (.ZN (n_6836), .A (A_imm[1]));
NAND2_X1 i_6899 (.ZN (n_6835), .A1 (B_imm[13]), .A2 (A_imm[18]));
OAI21_X1 i_6898 (.ZN (n_6834), .A (n_6835), .B1 (n_8860), .B2 (n_8926));
NAND2_X1 i_6897 (.ZN (n_6833), .A1 (B_imm[28]), .A2 (A_imm[3]));
NAND4_X1 i_6896 (.ZN (n_6832), .A1 (B_imm[20]), .A2 (B_imm[13]), .A3 (A_imm[18]), .A4 (A_imm[11]));
NAND2_X1 i_6895 (.ZN (n_6831), .A1 (n_6832), .A2 (n_6833));
NAND2_X1 i_6894 (.ZN (n_6830), .A1 (n_6831), .A2 (n_6834));
OAI21_X1 i_6893 (.ZN (n_6829), .A (n_6830), .B1 (n_9038), .B2 (n_6836));
NAND4_X1 i_6892 (.ZN (n_6828), .A1 (n_6831), .A2 (B_imm[31]), .A3 (A_imm[1]), .A4 (n_6834));
NAND2_X1 i_6891 (.ZN (n_6827), .A1 (n_7678), .A2 (n_7676));
NAND3_X1 i_6890 (.ZN (n_6826), .A1 (n_6827), .A2 (B_imm[16]), .A3 (A_imm[16]));
NAND3_X1 i_6889 (.ZN (n_6825), .A1 (n_7678), .A2 (n_7677), .A3 (n_7676));
NAND2_X1 i_6888 (.ZN (n_6824), .A1 (n_6826), .A2 (n_6825));
INV_X1 i_6887 (.ZN (n_6823), .A (n_6824));
NAND2_X1 i_6886 (.ZN (n_6822), .A1 (n_6828), .A2 (n_6823));
NAND2_X1 i_6885 (.ZN (n_6821), .A1 (n_6822), .A2 (n_6829));
NAND2_X1 i_6884 (.ZN (n_6820), .A1 (n_6821), .A2 (n_6837));
NAND4_X1 i_6883 (.ZN (n_6819), .A1 (n_6822), .A2 (n_6829), .A3 (B_imm[3]), .A4 (A_imm[30]));
INV_X1 i_6882 (.ZN (n_6818), .A (n_6819));
INV_X1 i_6881 (.ZN (n_6817), .A (B_imm[3]));
OAI22_X1 i_6880 (.ZN (n_6816), .A1 (n_8994), .A2 (n_6817), .B1 (n_7913), .B2 (n_8956));
OAI22_X1 i_6879 (.ZN (n_6815), .A1 (n_8908), .A2 (n_8971), .B1 (n_8927), .B2 (n_8909));
NAND2_X1 i_6878 (.ZN (n_6814), .A1 (A_imm[20]), .A2 (B_imm[10]));
NAND4_X1 i_6877 (.ZN (n_6813), .A1 (B_imm[16]), .A2 (A_imm[13]), .A3 (B_imm[17]), .A4 (A_imm[14]));
NAND2_X1 i_6876 (.ZN (n_6812), .A1 (n_6813), .A2 (n_6814));
NAND2_X1 i_6875 (.ZN (n_6811), .A1 (n_6812), .A2 (n_6815));
OAI21_X1 i_6874 (.ZN (n_6810), .A (n_6811), .B1 (n_8993), .B2 (n_8293));
NAND2_X1 i_6873 (.ZN (n_6809), .A1 (B_imm[19]), .A2 (A_imm[12]));
INV_X1 i_6872 (.ZN (n_6808), .A (n_6809));
NAND4_X1 i_6871 (.ZN (n_6807), .A1 (n_6812), .A2 (B_imm[26]), .A3 (n_6815), .A4 (A_imm[5]));
INV_X1 i_6870 (.ZN (n_6806), .A (n_6807));
OAI21_X1 i_6869 (.ZN (n_6805), .A (n_6810), .B1 (n_6806), .B2 (n_6808));
NAND4_X1 i_6868 (.ZN (n_6804), .A1 (A_imm[29]), .A2 (B_imm[14]), .A3 (B_imm[3]), .A4 (A_imm[18]));
NAND2_X1 i_6867 (.ZN (n_6803), .A1 (n_6804), .A2 (n_6805));
NAND2_X1 i_6866 (.ZN (n_6802), .A1 (n_6803), .A2 (n_6816));
INV_X1 i_6865 (.ZN (n_6801), .A (n_6802));
OAI21_X1 i_6864 (.ZN (n_6800), .A (n_6820), .B1 (n_6818), .B2 (n_6801));
NAND2_X1 i_6863 (.ZN (n_6799), .A1 (n_6800), .A2 (n_6838));
NAND2_X1 i_6862 (.ZN (n_6798), .A1 (n_7542), .A2 (n_7543));
NAND3_X1 i_6861 (.ZN (n_6797), .A1 (n_6798), .A2 (n_7540), .A3 (n_7539));
NAND3_X1 i_6860 (.ZN (n_6796), .A1 (n_7543), .A2 (n_7542), .A3 (n_7538));
NAND2_X1 i_6859 (.ZN (n_6795), .A1 (n_6797), .A2 (n_6796));
OAI21_X1 i_6858 (.ZN (n_6794), .A (n_6795), .B1 (n_6800), .B2 (n_6838));
NAND2_X1 i_6857 (.ZN (n_6793), .A1 (n_7602), .A2 (n_7601));
NAND3_X1 i_6856 (.ZN (n_6792), .A1 (n_6793), .A2 (n_7599), .A3 (n_7598));
NAND3_X1 i_6855 (.ZN (n_6791), .A1 (n_7602), .A2 (n_7601), .A3 (n_7597));
NAND4_X2 i_6854 (.ZN (n_6790), .A1 (n_6794), .A2 (n_6792), .A3 (n_6799), .A4 (n_6791));
NAND2_X1 i_6853 (.ZN (n_6789), .A1 (n_6794), .A2 (n_6799));
NAND2_X1 i_6852 (.ZN (n_6788), .A1 (n_6792), .A2 (n_6791));
NAND2_X1 i_6851 (.ZN (n_6787), .A1 (n_6789), .A2 (n_6788));
NOR2_X1 i_6850 (.ZN (n_6786), .A1 (n_7500), .A2 (n_7507));
NAND2_X1 i_6849 (.ZN (n_6785), .A1 (n_7530), .A2 (n_7531));
NAND2_X1 i_6848 (.ZN (n_6784), .A1 (n_6785), .A2 (n_6786));
OAI211_X1 i_6847 (.ZN (n_6783), .A (n_7531), .B (n_7530), .C1 (n_7507), .C2 (n_7500));
NAND2_X1 i_6846 (.ZN (n_6782), .A1 (n_6783), .A2 (n_6784));
INV_X1 i_6845 (.ZN (n_6781), .A (n_6782));
NAND2_X1 i_6844 (.ZN (n_6780), .A1 (n_6787), .A2 (n_6781));
NAND2_X1 i_6843 (.ZN (n_6779), .A1 (n_6780), .A2 (n_6790));
NAND2_X4 i_6842 (.ZN (n_6778), .A1 (n_6779), .A2 (n_6843));
NAND3_X2 i_6841 (.ZN (n_6777), .A1 (n_6780), .A2 (n_6844), .A3 (n_6790));
INV_X1 i_6840 (.ZN (n_6776), .A (n_7490));
NAND3_X1 i_6839 (.ZN (n_6775), .A1 (n_7497), .A2 (n_7494), .A3 (n_6776));
INV_X1 i_6838 (.ZN (n_6774), .A (n_7494));
OAI21_X1 i_6837 (.ZN (n_6773), .A (n_7490), .B1 (n_7498), .B2 (n_6774));
NAND2_X2 i_6836 (.ZN (n_6772), .A1 (n_6773), .A2 (n_6775));
NAND2_X1 i_6835 (.ZN (n_6771), .A1 (n_6777), .A2 (n_6772));
NAND2_X1 i_6834 (.ZN (n_6770), .A1 (n_6771), .A2 (n_6778));
NAND3_X1 i_6833 (.ZN (n_6769), .A1 (n_6770), .A2 (n_6852), .A3 (n_6849));
NAND2_X1 i_6832 (.ZN (n_6768), .A1 (n_6849), .A2 (n_6852));
NAND3_X1 i_6831 (.ZN (n_6767), .A1 (n_6768), .A2 (n_6778), .A3 (n_6771));
NAND2_X1 i_6830 (.ZN (n_6766), .A1 (n_6767), .A2 (n_6769));
NAND3_X1 i_6829 (.ZN (n_6765), .A1 (n_6778), .A2 (n_6777), .A3 (n_6772));
INV_X1 i_6828 (.ZN (n_6764), .A (n_6765));
AOI21_X2 i_6827 (.ZN (n_6763), .A (n_6772), .B1 (n_6778), .B2 (n_6777));
NOR2_X1 i_6826 (.ZN (n_6762), .A1 (n_6764), .A2 (n_6763));
OAI21_X1 i_6825 (.ZN (n_6761), .A (n_8086), .B1 (n_8094), .B2 (n_8097));
NAND3_X1 i_6824 (.ZN (n_6760), .A1 (n_8096), .A2 (n_8095), .A3 (n_8087));
AOI21_X1 i_6823 (.ZN (n_6759), .A (n_7660), .B1 (n_7664), .B2 (n_7667));
NAND3_X1 i_6822 (.ZN (n_6758), .A1 (n_7664), .A2 (n_7667), .A3 (n_7660));
INV_X1 i_6821 (.ZN (n_6757), .A (n_6758));
OAI211_X1 i_6820 (.ZN (n_6756), .A (n_6761), .B (n_6760), .C1 (n_6759), .C2 (n_6757));
NAND2_X1 i_6819 (.ZN (n_6755), .A1 (n_6761), .A2 (n_6760));
NOR2_X1 i_6818 (.ZN (n_6754), .A1 (n_6757), .A2 (n_6759));
NAND2_X1 i_6817 (.ZN (n_6753), .A1 (n_6755), .A2 (n_6754));
OAI22_X1 i_6816 (.ZN (n_6752), .A1 (n_8347), .A2 (n_8906), .B1 (n_8794), .B2 (n_8232));
NAND2_X1 i_6815 (.ZN (n_6751), .A1 (B_imm[24]), .A2 (A_imm[7]));
NAND4_X1 i_6814 (.ZN (n_6750), .A1 (B_imm[9]), .A2 (A_imm[25]), .A3 (B_imm[6]), .A4 (A_imm[22]));
NAND2_X1 i_6813 (.ZN (n_6749), .A1 (n_6750), .A2 (n_6751));
NAND2_X1 i_6812 (.ZN (n_6748), .A1 (n_6749), .A2 (n_6752));
NAND2_X1 i_6811 (.ZN (n_6747), .A1 (B_imm[11]), .A2 (A_imm[20]));
OAI21_X1 i_6810 (.ZN (n_6746), .A (n_6747), .B1 (n_8972), .B2 (n_8429));
NAND2_X1 i_6809 (.ZN (n_6745), .A1 (B_imm[18]), .A2 (A_imm[13]));
NAND4_X1 i_6808 (.ZN (n_6744), .A1 (A_imm[26]), .A2 (B_imm[11]), .A3 (B_imm[5]), .A4 (A_imm[20]));
NAND2_X1 i_6807 (.ZN (n_6743), .A1 (n_6744), .A2 (n_6745));
NAND2_X1 i_6806 (.ZN (n_6742), .A1 (n_6743), .A2 (n_6746));
NAND2_X1 i_6805 (.ZN (n_6741), .A1 (n_6748), .A2 (n_6742));
INV_X1 i_6804 (.ZN (n_6740), .A (B_imm[0]));
OAI22_X1 i_6803 (.ZN (n_6739), .A1 (n_8821), .A2 (n_8511), .B1 (n_9037), .B2 (n_6740));
NAND2_X1 i_6802 (.ZN (n_6738), .A1 (B_imm[21]), .A2 (A_imm[10]));
INV_X1 i_6801 (.ZN (n_6737), .A (n_6738));
NAND4_X1 i_6800 (.ZN (n_6736), .A1 (B_imm[23]), .A2 (A_imm[31]), .A3 (B_imm[0]), .A4 (A_imm[8]));
INV_X1 i_6799 (.ZN (n_6735), .A (n_6736));
OAI21_X1 i_6798 (.ZN (n_6734), .A (n_6739), .B1 (n_6737), .B2 (n_6735));
NAND4_X1 i_6797 (.ZN (n_6733), .A1 (n_6752), .A2 (n_6749), .A3 (n_6743), .A4 (n_6746));
NAND2_X1 i_6796 (.ZN (n_6732), .A1 (n_6733), .A2 (n_6734));
NAND2_X1 i_6795 (.ZN (n_6731), .A1 (n_6732), .A2 (n_6741));
INV_X1 i_6794 (.ZN (n_6730), .A (n_8116));
OAI21_X1 i_6793 (.ZN (n_6729), .A (n_8114), .B1 (n_6730), .B2 (n_8112));
NAND3_X1 i_6792 (.ZN (n_6728), .A1 (n_8116), .A2 (n_8115), .A3 (n_8113));
NAND3_X1 i_6791 (.ZN (n_6727), .A1 (n_6731), .A2 (n_6729), .A3 (n_6728));
NAND2_X1 i_6790 (.ZN (n_6726), .A1 (n_6729), .A2 (n_6728));
NAND3_X1 i_6789 (.ZN (n_6725), .A1 (n_6732), .A2 (n_6741), .A3 (n_6726));
NAND2_X1 i_6788 (.ZN (n_6724), .A1 (A_imm[27]), .A2 (B_imm[5]));
NAND2_X1 i_6787 (.ZN (n_6723), .A1 (B_imm[22]), .A2 (A_imm[9]));
OAI21_X1 i_6786 (.ZN (n_6722), .A (n_6723), .B1 (n_8829), .B2 (n_8858));
NAND2_X1 i_6785 (.ZN (n_6721), .A1 (B_imm[25]), .A2 (A_imm[6]));
NAND4_X1 i_6784 (.ZN (n_6720), .A1 (B_imm[15]), .A2 (B_imm[22]), .A3 (A_imm[16]), .A4 (A_imm[9]));
NAND2_X1 i_6783 (.ZN (n_6719), .A1 (n_6720), .A2 (n_6721));
NAND2_X1 i_6782 (.ZN (n_6718), .A1 (n_6719), .A2 (n_6722));
NAND2_X1 i_6781 (.ZN (n_6717), .A1 (n_6718), .A2 (n_6724));
NAND2_X1 i_6780 (.ZN (n_6716), .A1 (B_imm[30]), .A2 (A_imm[2]));
INV_X1 i_6779 (.ZN (n_6715), .A (n_6716));
NAND4_X1 i_6778 (.ZN (n_6714), .A1 (n_6719), .A2 (B_imm[5]), .A3 (A_imm[27]), .A4 (n_6722));
INV_X1 i_6777 (.ZN (n_6713), .A (n_6714));
OAI21_X1 i_6776 (.ZN (n_6712), .A (n_6717), .B1 (n_6713), .B2 (n_6715));
NAND2_X1 i_6775 (.ZN (n_6711), .A1 (n_6725), .A2 (n_6712));
NAND2_X1 i_6774 (.ZN (n_6710), .A1 (n_6711), .A2 (n_6727));
NAND2_X1 i_6773 (.ZN (n_6709), .A1 (n_6710), .A2 (n_6753));
AOI21_X1 i_6772 (.ZN (n_6708), .A (n_8133), .B1 (n_8138), .B2 (n_8141));
NAND3_X1 i_6771 (.ZN (n_6707), .A1 (n_8138), .A2 (n_8141), .A3 (n_8133));
INV_X1 i_6770 (.ZN (n_6706), .A (n_6707));
NOR2_X1 i_6769 (.ZN (n_6705), .A1 (n_6706), .A2 (n_6708));
AOI21_X1 i_6768 (.ZN (n_6704), .A (n_6705), .B1 (n_6709), .B2 (n_6756));
INV_X1 i_6767 (.ZN (n_6703), .A (n_6704));
NAND3_X1 i_6766 (.ZN (n_6702), .A1 (n_6709), .A2 (n_6756), .A3 (n_6705));
NAND2_X1 i_6765 (.ZN (n_6701), .A1 (n_8106), .A2 (n_8103));
NAND2_X1 i_6764 (.ZN (n_6700), .A1 (n_6701), .A2 (n_8085));
NAND3_X1 i_6763 (.ZN (n_6699), .A1 (n_8103), .A2 (n_8106), .A3 (n_8084));
NAND4_X1 i_6762 (.ZN (n_6698), .A1 (n_6703), .A2 (n_6702), .A3 (n_6700), .A4 (n_6699));
INV_X1 i_6761 (.ZN (n_6697), .A (n_6702));
NAND2_X1 i_6760 (.ZN (n_6696), .A1 (n_6700), .A2 (n_6699));
OAI21_X1 i_6759 (.ZN (n_6695), .A (n_6696), .B1 (n_6697), .B2 (n_6704));
NAND2_X1 i_6758 (.ZN (n_6694), .A1 (n_6698), .A2 (n_6695));
INV_X1 i_6757 (.ZN (n_6693), .A (n_6694));
AOI21_X1 i_6756 (.ZN (n_6692), .A (n_6866), .B1 (n_6873), .B2 (n_6870));
NAND3_X1 i_6755 (.ZN (n_6691), .A1 (n_6870), .A2 (n_6873), .A3 (n_6866));
INV_X1 i_6754 (.ZN (n_6690), .A (n_6691));
NOR2_X1 i_6753 (.ZN (n_6689), .A1 (n_6690), .A2 (n_6692));
NAND2_X1 i_6752 (.ZN (n_6688), .A1 (n_6879), .A2 (n_6878));
INV_X1 i_6751 (.ZN (n_6687), .A (n_6688));
NAND2_X1 i_6750 (.ZN (n_6686), .A1 (n_6876), .A2 (n_6875));
INV_X1 i_6749 (.ZN (n_6685), .A (n_6686));
OAI21_X1 i_6748 (.ZN (n_6684), .A (n_6685), .B1 (n_6687), .B2 (n_6882));
NAND3_X1 i_6747 (.ZN (n_6683), .A1 (n_6688), .A2 (n_6883), .A3 (n_6686));
AOI22_X1 i_6746 (.ZN (n_6682), .A1 (n_6893), .A2 (n_6896), .B1 (B_imm[29]), .B2 (A_imm[3]));
OAI21_X1 i_6745 (.ZN (n_6681), .A (n_6881), .B1 (n_6880), .B2 (n_6682));
NAND3_X1 i_6744 (.ZN (n_6680), .A1 (n_6891), .A2 (n_6889), .A3 (n_6890));
NAND2_X1 i_6743 (.ZN (n_6679), .A1 (n_6681), .A2 (n_6680));
INV_X2 i_6742 (.ZN (n_6678), .A (A_imm[4]));
INV_X4 i_6741 (.ZN (n_6677), .A (A_imm[2]));
OAI22_X1 i_6740 (.ZN (n_6676), .A1 (n_9021), .A2 (n_6677), .B1 (n_8993), .B2 (n_6678));
NAND2_X1 i_6739 (.ZN (n_6675), .A1 (B_imm[19]), .A2 (A_imm[11]));
NAND4_X1 i_6738 (.ZN (n_6674), .A1 (B_imm[28]), .A2 (B_imm[26]), .A3 (A_imm[4]), .A4 (A_imm[2]));
NAND2_X1 i_6737 (.ZN (n_6673), .A1 (n_6674), .A2 (n_6675));
OAI22_X2 i_6736 (.ZN (n_6672), .A1 (n_8908), .A2 (n_8946), .B1 (n_8909), .B2 (n_8971));
NAND4_X1 i_6735 (.ZN (n_6671), .A1 (B_imm[16]), .A2 (B_imm[17]), .A3 (A_imm[15]), .A4 (A_imm[14]));
NAND2_X1 i_6734 (.ZN (n_6670), .A1 (n_6672), .A2 (n_6671));
NAND3_X1 i_6733 (.ZN (n_6669), .A1 (n_6670), .A2 (B_imm[10]), .A3 (A_imm[21]));
NAND2_X1 i_6732 (.ZN (n_6668), .A1 (A_imm[21]), .A2 (B_imm[10]));
NAND3_X1 i_6731 (.ZN (n_6667), .A1 (n_6672), .A2 (n_6668), .A3 (n_6671));
NAND2_X1 i_6730 (.ZN (n_6666), .A1 (n_6669), .A2 (n_6667));
NAND3_X1 i_6729 (.ZN (n_6665), .A1 (n_6673), .A2 (n_6676), .A3 (n_6666));
NAND2_X1 i_6728 (.ZN (n_6664), .A1 (B_imm[14]), .A2 (A_imm[17]));
AOI21_X1 i_6727 (.ZN (n_6663), .A (n_6666), .B1 (n_6676), .B2 (n_6673));
OAI21_X1 i_6726 (.ZN (n_6662), .A (n_6665), .B1 (n_6663), .B2 (n_6664));
NAND2_X1 i_6725 (.ZN (n_6661), .A1 (n_6662), .A2 (n_6679));
INV_X1 i_6724 (.ZN (n_6660), .A (n_6679));
INV_X1 i_6723 (.ZN (n_6659), .A (n_6662));
NAND2_X1 i_6722 (.ZN (n_6658), .A1 (n_6659), .A2 (n_6660));
NAND2_X1 i_6721 (.ZN (n_6657), .A1 (A_imm[29]), .A2 (B_imm[2]));
INV_X1 i_6720 (.ZN (n_6656), .A (n_6657));
OAI22_X1 i_6719 (.ZN (n_6655), .A1 (n_8947), .A2 (n_8859), .B1 (n_8752), .B2 (n_8909));
NAND2_X1 i_6718 (.ZN (n_6654), .A1 (A_imm[24]), .A2 (B_imm[5]));
NAND4_X1 i_6717 (.ZN (n_6653), .A1 (B_imm[8]), .A2 (B_imm[17]), .A3 (A_imm[21]), .A4 (A_imm[12]));
NAND2_X1 i_6716 (.ZN (n_6652), .A1 (n_6653), .A2 (n_6654));
AOI22_X1 i_6715 (.ZN (n_6651), .A1 (n_6652), .A2 (n_6655), .B1 (B_imm[27]), .B2 (A_imm[3]));
INV_X1 i_6714 (.ZN (n_6650), .A (n_6651));
NAND2_X1 i_6713 (.ZN (n_6649), .A1 (B_imm[29]), .A2 (A_imm[1]));
NAND4_X1 i_6712 (.ZN (n_6648), .A1 (n_6652), .A2 (n_6655), .A3 (B_imm[27]), .A4 (A_imm[3]));
NAND2_X1 i_6711 (.ZN (n_6647), .A1 (n_6648), .A2 (n_6649));
NAND3_X1 i_6710 (.ZN (n_6646), .A1 (n_6656), .A2 (n_6650), .A3 (n_6647));
NAND2_X1 i_6709 (.ZN (n_6645), .A1 (n_6647), .A2 (n_6650));
NAND2_X1 i_6708 (.ZN (n_6644), .A1 (n_6645), .A2 (n_6657));
INV_X1 i_6707 (.ZN (n_6643), .A (n_6644));
NAND2_X1 i_6706 (.ZN (n_6642), .A1 (n_6896), .A2 (n_6894));
INV_X1 i_6705 (.ZN (n_6641), .A (n_6642));
NOR2_X1 i_6704 (.ZN (n_6640), .A1 (n_6641), .A2 (n_6895));
NAND2_X1 i_6703 (.ZN (n_6639), .A1 (n_6641), .A2 (n_6895));
INV_X1 i_6702 (.ZN (n_6638), .A (n_6639));
NOR2_X1 i_6701 (.ZN (n_6637), .A1 (n_6638), .A2 (n_6640));
OAI21_X1 i_6700 (.ZN (n_6636), .A (n_6646), .B1 (n_6643), .B2 (n_6637));
NAND2_X1 i_6699 (.ZN (n_6635), .A1 (n_6658), .A2 (n_6636));
NAND2_X1 i_6698 (.ZN (n_6634), .A1 (n_6635), .A2 (n_6661));
NAND3_X1 i_6697 (.ZN (n_6633), .A1 (n_6634), .A2 (n_6684), .A3 (n_6683));
NAND2_X1 i_6696 (.ZN (n_6632), .A1 (n_6684), .A2 (n_6683));
NAND3_X1 i_6695 (.ZN (n_6631), .A1 (n_6635), .A2 (n_6632), .A3 (n_6661));
NAND3_X1 i_6694 (.ZN (n_6630), .A1 (n_6727), .A2 (n_6725), .A3 (n_6712));
INV_X1 i_6693 (.ZN (n_6629), .A (n_6712));
NAND2_X1 i_6692 (.ZN (n_6628), .A1 (n_6727), .A2 (n_6725));
NAND2_X1 i_6691 (.ZN (n_6627), .A1 (n_6628), .A2 (n_6629));
NAND2_X1 i_6690 (.ZN (n_6626), .A1 (n_6627), .A2 (n_6630));
NAND2_X1 i_6689 (.ZN (n_6625), .A1 (n_6631), .A2 (n_6626));
NAND2_X1 i_6688 (.ZN (n_6624), .A1 (n_6625), .A2 (n_6633));
NAND2_X1 i_6687 (.ZN (n_6623), .A1 (n_6624), .A2 (n_6689));
INV_X1 i_6686 (.ZN (n_6622), .A (n_6623));
INV_X1 i_6685 (.ZN (n_6621), .A (n_6689));
INV_X1 i_6684 (.ZN (n_6620), .A (n_6624));
NAND3_X1 i_6683 (.ZN (n_6619), .A1 (n_6710), .A2 (n_6753), .A3 (n_6756));
NAND2_X1 i_6682 (.ZN (n_6618), .A1 (n_6756), .A2 (n_6753));
NAND3_X1 i_6681 (.ZN (n_6617), .A1 (n_6618), .A2 (n_6727), .A3 (n_6711));
NAND2_X1 i_6680 (.ZN (n_6616), .A1 (n_6617), .A2 (n_6619));
INV_X1 i_6679 (.ZN (n_6615), .A (n_6616));
AOI21_X1 i_6678 (.ZN (n_6614), .A (n_6615), .B1 (n_6620), .B2 (n_6621));
OAI21_X1 i_6677 (.ZN (n_6613), .A (n_6693), .B1 (n_6614), .B2 (n_6622));
NAND2_X1 i_6676 (.ZN (n_6612), .A1 (n_6620), .A2 (n_6621));
NAND2_X1 i_6675 (.ZN (n_6611), .A1 (n_6612), .A2 (n_6616));
NAND3_X1 i_6674 (.ZN (n_6610), .A1 (n_6611), .A2 (n_6694), .A3 (n_6623));
NAND3_X1 i_6673 (.ZN (n_6609), .A1 (n_6916), .A2 (n_6914), .A3 (n_6864));
NAND2_X1 i_6672 (.ZN (n_6608), .A1 (n_6916), .A2 (n_6914));
NAND3_X1 i_6671 (.ZN (n_6607), .A1 (n_6608), .A2 (n_6873), .A3 (n_6865));
NAND2_X1 i_6670 (.ZN (n_6606), .A1 (n_6607), .A2 (n_6609));
INV_X1 i_6669 (.ZN (n_6605), .A (n_6606));
NAND2_X1 i_6668 (.ZN (n_6604), .A1 (n_6610), .A2 (n_6605));
NAND2_X1 i_6667 (.ZN (n_6603), .A1 (n_6604), .A2 (n_6613));
NAND2_X1 i_6666 (.ZN (n_6602), .A1 (n_6762), .A2 (n_6603));
OAI211_X1 i_6665 (.ZN (n_6601), .A (n_6613), .B (n_6604), .C1 (n_6764), .C2 (n_6763));
NAND3_X1 i_6664 (.ZN (n_6600), .A1 (n_6787), .A2 (n_6790), .A3 (n_6781));
NAND2_X1 i_6663 (.ZN (n_6599), .A1 (n_6787), .A2 (n_6790));
NAND2_X1 i_6662 (.ZN (n_6598), .A1 (n_6599), .A2 (n_6782));
NAND2_X1 i_6661 (.ZN (n_6597), .A1 (n_6598), .A2 (n_6600));
INV_X1 i_6660 (.ZN (n_6596), .A (n_6597));
INV_X1 i_6659 (.ZN (n_6595), .A (n_6734));
NAND2_X1 i_6658 (.ZN (n_6594), .A1 (n_6733), .A2 (n_6741));
NAND2_X1 i_6657 (.ZN (n_6593), .A1 (n_6594), .A2 (n_6595));
NAND3_X1 i_6656 (.ZN (n_6592), .A1 (n_6741), .A2 (n_6733), .A3 (n_6734));
NAND2_X1 i_6655 (.ZN (n_6591), .A1 (n_6593), .A2 (n_6592));
NAND2_X1 i_6654 (.ZN (n_6590), .A1 (n_6717), .A2 (n_6714));
NAND2_X1 i_6653 (.ZN (n_6589), .A1 (n_6590), .A2 (n_6715));
NAND3_X1 i_6652 (.ZN (n_6588), .A1 (n_6717), .A2 (n_6714), .A3 (n_6716));
NAND2_X1 i_6651 (.ZN (n_6587), .A1 (n_6589), .A2 (n_6588));
NAND2_X1 i_6650 (.ZN (n_6586), .A1 (n_6587), .A2 (n_6591));
NAND4_X1 i_6649 (.ZN (n_6585), .A1 (n_6589), .A2 (n_6593), .A3 (n_6592), .A4 (n_6588));
INV_X2 i_6648 (.ZN (n_6584), .A (B_imm[2]));
OAI22_X1 i_6647 (.ZN (n_6583), .A1 (n_8795), .A2 (n_8955), .B1 (n_8907), .B2 (n_8232));
NAND2_X1 i_6646 (.ZN (n_6582), .A1 (B_imm[11]), .A2 (A_imm[18]));
NAND4_X1 i_6645 (.ZN (n_6581), .A1 (B_imm[12]), .A2 (A_imm[23]), .A3 (B_imm[6]), .A4 (A_imm[17]));
NAND2_X1 i_6644 (.ZN (n_6580), .A1 (n_6581), .A2 (n_6582));
NAND2_X1 i_6643 (.ZN (n_6579), .A1 (n_6580), .A2 (n_6583));
OAI21_X1 i_6642 (.ZN (n_6578), .A (n_6579), .B1 (n_6584), .B2 (n_9020));
INV_X2 i_6641 (.ZN (n_6577), .A (B_imm[4]));
OAI22_X1 i_6640 (.ZN (n_6576), .A1 (n_6577), .A2 (n_8794), .B1 (n_8972), .B2 (n_6817));
NAND2_X1 i_6639 (.ZN (n_6575), .A1 (B_imm[18]), .A2 (A_imm[11]));
INV_X1 i_6638 (.ZN (n_6574), .A (n_6575));
NAND4_X1 i_6637 (.ZN (n_6573), .A1 (A_imm[26]), .A2 (A_imm[25]), .A3 (B_imm[4]), .A4 (B_imm[3]));
INV_X1 i_6636 (.ZN (n_6572), .A (n_6573));
OAI21_X2 i_6635 (.ZN (n_6571), .A (n_6576), .B1 (n_6574), .B2 (n_6572));
NAND4_X1 i_6634 (.ZN (n_6570), .A1 (n_6580), .A2 (n_6583), .A3 (B_imm[2]), .A4 (A_imm[28]));
NAND2_X1 i_6633 (.ZN (n_6569), .A1 (n_6570), .A2 (n_6571));
INV_X1 i_6632 (.ZN (n_6568), .A (n_6745));
NAND2_X1 i_6631 (.ZN (n_6567), .A1 (n_6746), .A2 (n_6744));
NAND2_X1 i_6630 (.ZN (n_6566), .A1 (n_6567), .A2 (n_6568));
NAND3_X1 i_6629 (.ZN (n_6565), .A1 (n_6746), .A2 (n_6745), .A3 (n_6744));
NAND2_X1 i_6628 (.ZN (n_6564), .A1 (n_6566), .A2 (n_6565));
NAND3_X1 i_6627 (.ZN (n_6563), .A1 (n_6569), .A2 (n_6578), .A3 (n_6564));
AOI21_X1 i_6626 (.ZN (n_6562), .A (n_6564), .B1 (n_6578), .B2 (n_6569));
NAND2_X1 i_6625 (.ZN (n_6561), .A1 (n_6752), .A2 (n_6750));
XNOR2_X1 i_6624 (.ZN (n_6560), .A (n_6561), .B (n_6751));
OAI21_X1 i_6623 (.ZN (n_6559), .A (n_6563), .B1 (n_6562), .B2 (n_6560));
NAND2_X1 i_6622 (.ZN (n_6558), .A1 (n_6585), .A2 (n_6559));
NAND2_X1 i_6621 (.ZN (n_6557), .A1 (n_6558), .A2 (n_6586));
NAND3_X1 i_6620 (.ZN (n_6556), .A1 (n_6820), .A2 (n_6819), .A3 (n_6802));
NAND2_X1 i_6619 (.ZN (n_6555), .A1 (n_6820), .A2 (n_6819));
NAND2_X1 i_6618 (.ZN (n_6554), .A1 (n_6555), .A2 (n_6801));
NAND2_X1 i_6617 (.ZN (n_6553), .A1 (n_6554), .A2 (n_6556));
NAND2_X1 i_6616 (.ZN (n_6552), .A1 (n_6553), .A2 (n_6557));
NAND4_X1 i_6615 (.ZN (n_6551), .A1 (n_6558), .A2 (n_6554), .A3 (n_6586), .A4 (n_6556));
INV_X1 i_6614 (.ZN (n_6550), .A (n_6551));
NAND2_X1 i_6613 (.ZN (n_6549), .A1 (n_6904), .A2 (n_6907));
XNOR2_X1 i_6612 (.ZN (n_6548), .A (n_6549), .B (n_6900));
OAI21_X1 i_6611 (.ZN (n_6547), .A (n_6552), .B1 (n_6550), .B2 (n_6548));
AOI21_X1 i_6610 (.ZN (n_6546), .A (n_7606), .B1 (n_7613), .B2 (n_7614));
NAND3_X1 i_6609 (.ZN (n_6545), .A1 (n_7614), .A2 (n_7613), .A3 (n_7606));
INV_X1 i_6608 (.ZN (n_6544), .A (n_6545));
NOR2_X1 i_6607 (.ZN (n_6543), .A1 (n_6544), .A2 (n_6546));
NAND2_X1 i_6606 (.ZN (n_6542), .A1 (B_imm[8]), .A2 (A_imm[22]));
OAI21_X1 i_6605 (.ZN (n_6541), .A (n_6542), .B1 (n_8907), .B2 (n_8573));
NAND2_X1 i_6604 (.ZN (n_6540), .A1 (A_imm[24]), .A2 (B_imm[6]));
NAND4_X1 i_6603 (.ZN (n_6539), .A1 (A_imm[23]), .A2 (B_imm[8]), .A3 (B_imm[7]), .A4 (A_imm[22]));
NAND2_X1 i_6602 (.ZN (n_6538), .A1 (n_6539), .A2 (n_6540));
NAND2_X1 i_6601 (.ZN (n_6537), .A1 (n_6538), .A2 (n_6541));
OAI21_X1 i_6600 (.ZN (n_6536), .A (n_6537), .B1 (CLOCK_opt_ipo_n433), .B2 (n_6678));
NAND2_X1 i_6599 (.ZN (n_6535), .A1 (B_imm[29]), .A2 (A_imm[2]));
NAND4_X1 i_6598 (.ZN (n_6534), .A1 (n_6538), .A2 (B_imm[27]), .A3 (A_imm[4]), .A4 (n_6541));
NAND2_X1 i_6597 (.ZN (n_6533), .A1 (n_6534), .A2 (n_6535));
INV_X1 i_6596 (.ZN (n_6532), .A (n_7611));
OAI21_X1 i_6595 (.ZN (n_6531), .A (n_7609), .B1 (n_6532), .B2 (n_7607));
NAND3_X1 i_6594 (.ZN (n_6530), .A1 (n_7611), .A2 (n_7610), .A3 (n_7608));
NAND2_X1 i_6593 (.ZN (n_6529), .A1 (n_6531), .A2 (n_6530));
NAND3_X1 i_6592 (.ZN (n_6528), .A1 (n_6529), .A2 (n_6536), .A3 (n_6533));
INV_X1 i_6591 (.ZN (n_6527), .A (n_6535));
INV_X1 i_6590 (.ZN (n_6526), .A (n_6534));
OAI21_X1 i_6589 (.ZN (n_6525), .A (n_6536), .B1 (n_6526), .B2 (n_6527));
AOI21_X1 i_6588 (.ZN (n_6524), .A (n_7610), .B1 (n_7611), .B2 (n_7608));
INV_X1 i_6587 (.ZN (n_6523), .A (n_6530));
NOR2_X1 i_6586 (.ZN (n_6522), .A1 (n_6523), .A2 (n_6524));
NAND2_X1 i_6585 (.ZN (n_6521), .A1 (n_6525), .A2 (n_6522));
AOI21_X1 i_6584 (.ZN (n_6520), .A (n_7618), .B1 (n_7619), .B2 (n_7617));
NAND3_X1 i_6583 (.ZN (n_6519), .A1 (n_7619), .A2 (n_7618), .A3 (n_7617));
INV_X1 i_6582 (.ZN (n_6518), .A (n_6519));
NOR2_X1 i_6581 (.ZN (n_6517), .A1 (n_6520), .A2 (n_6518));
INV_X1 i_6580 (.ZN (n_6516), .A (n_6517));
NAND2_X1 i_6579 (.ZN (n_6515), .A1 (n_6521), .A2 (n_6516));
NAND3_X1 i_6578 (.ZN (n_6514), .A1 (n_6543), .A2 (n_6515), .A3 (n_6528));
INV_X1 i_6577 (.ZN (n_6513), .A (n_6528));
AOI21_X1 i_6576 (.ZN (n_6512), .A (n_6517), .B1 (n_6525), .B2 (n_6522));
OAI22_X1 i_6575 (.ZN (n_6511), .A1 (n_6512), .A2 (n_6513), .B1 (n_6546), .B2 (n_6544));
NAND2_X1 i_6574 (.ZN (n_6510), .A1 (n_6511), .A2 (n_6514));
NAND2_X1 i_6573 (.ZN (n_6509), .A1 (n_7515), .A2 (n_7517));
NAND3_X1 i_6572 (.ZN (n_6508), .A1 (n_6509), .A2 (B_imm[6]), .A3 (A_imm[27]));
NAND3_X1 i_6571 (.ZN (n_6507), .A1 (n_7515), .A2 (n_7517), .A3 (n_7514));
NAND2_X1 i_6570 (.ZN (n_6506), .A1 (n_6508), .A2 (n_6507));
INV_X1 i_6569 (.ZN (n_6505), .A (n_6506));
NAND2_X1 i_6568 (.ZN (n_6504), .A1 (n_6510), .A2 (n_6505));
NAND3_X1 i_6567 (.ZN (n_6503), .A1 (n_6511), .A2 (n_6514), .A3 (n_6506));
INV_X1 i_6566 (.ZN (n_6502), .A (n_6805));
NAND2_X1 i_6565 (.ZN (n_6501), .A1 (n_6816), .A2 (n_6804));
NAND2_X1 i_6564 (.ZN (n_6500), .A1 (n_6501), .A2 (n_6502));
NAND3_X1 i_6563 (.ZN (n_6499), .A1 (n_6816), .A2 (n_6805), .A3 (n_6804));
NAND2_X1 i_6562 (.ZN (n_6498), .A1 (n_6500), .A2 (n_6499));
NAND3_X1 i_6561 (.ZN (n_6497), .A1 (n_6829), .A2 (n_6828), .A3 (n_6823));
NAND2_X1 i_6560 (.ZN (n_6496), .A1 (n_6829), .A2 (n_6828));
NAND2_X1 i_6559 (.ZN (n_6495), .A1 (n_6496), .A2 (n_6824));
NAND2_X1 i_6558 (.ZN (n_6494), .A1 (n_6495), .A2 (n_6497));
NAND2_X1 i_6557 (.ZN (n_6493), .A1 (n_6498), .A2 (n_6494));
AOI21_X1 i_6556 (.ZN (n_6492), .A (n_6721), .B1 (n_6722), .B2 (n_6720));
NAND3_X1 i_6555 (.ZN (n_6491), .A1 (n_6722), .A2 (n_6721), .A3 (n_6720));
INV_X1 i_6554 (.ZN (n_6490), .A (n_6491));
AOI21_X1 i_6553 (.ZN (n_6489), .A (n_6738), .B1 (n_6739), .B2 (n_6736));
NAND3_X1 i_6552 (.ZN (n_6488), .A1 (n_6739), .A2 (n_6738), .A3 (n_6736));
INV_X1 i_6551 (.ZN (n_6487), .A (n_6488));
OAI22_X1 i_6550 (.ZN (n_6486), .A1 (n_6492), .A2 (n_6490), .B1 (n_6489), .B2 (n_6487));
NAND2_X1 i_6549 (.ZN (n_6485), .A1 (A_imm[27]), .A2 (B_imm[3]));
NAND2_X1 i_6548 (.ZN (n_6484), .A1 (B_imm[9]), .A2 (A_imm[20]));
OAI21_X1 i_6547 (.ZN (n_6483), .A (n_6484), .B1 (n_8948), .B2 (n_8293));
NAND2_X1 i_6546 (.ZN (n_6482), .A1 (B_imm[23]), .A2 (A_imm[6]));
INV_X1 i_6545 (.ZN (n_6481), .A (n_6482));
NAND4_X1 i_6544 (.ZN (n_6480), .A1 (B_imm[24]), .A2 (B_imm[9]), .A3 (A_imm[20]), .A4 (A_imm[5]));
INV_X1 i_6543 (.ZN (n_6479), .A (n_6480));
OAI21_X1 i_6542 (.ZN (n_6478), .A (n_6483), .B1 (n_6479), .B2 (n_6481));
NAND2_X1 i_6541 (.ZN (n_6477), .A1 (n_6478), .A2 (n_6485));
NAND2_X1 i_6540 (.ZN (n_6476), .A1 (B_imm[15]), .A2 (A_imm[14]));
OAI21_X1 i_6539 (.ZN (n_6475), .A (n_6476), .B1 (n_8974), .B2 (n_6678));
NAND2_X1 i_6538 (.ZN (n_6474), .A1 (B_imm[13]), .A2 (A_imm[16]));
INV_X1 i_6537 (.ZN (n_6473), .A (n_6474));
NAND4_X1 i_6536 (.ZN (n_6472), .A1 (B_imm[25]), .A2 (B_imm[15]), .A3 (A_imm[14]), .A4 (A_imm[4]));
INV_X1 i_6535 (.ZN (n_6471), .A (n_6472));
OAI21_X1 i_6534 (.ZN (n_6470), .A (n_6475), .B1 (n_6471), .B2 (n_6473));
NAND2_X1 i_6533 (.ZN (n_6469), .A1 (n_6480), .A2 (n_6482));
NAND4_X1 i_6532 (.ZN (n_6468), .A1 (n_6469), .A2 (B_imm[3]), .A3 (A_imm[27]), .A4 (n_6483));
NAND2_X1 i_6531 (.ZN (n_6467), .A1 (n_6468), .A2 (n_6470));
NAND2_X1 i_6530 (.ZN (n_6466), .A1 (n_6467), .A2 (n_6477));
INV_X1 i_6529 (.ZN (n_6465), .A (n_6466));
NOR2_X1 i_6528 (.ZN (n_6464), .A1 (n_6490), .A2 (n_6492));
NOR2_X1 i_6527 (.ZN (n_6463), .A1 (n_6489), .A2 (n_6487));
NAND2_X1 i_6526 (.ZN (n_6462), .A1 (n_6464), .A2 (n_6463));
NAND2_X1 i_6525 (.ZN (n_6461), .A1 (n_6465), .A2 (n_6462));
NAND2_X1 i_6524 (.ZN (n_6460), .A1 (n_6461), .A2 (n_6486));
NAND4_X1 i_6523 (.ZN (n_6459), .A1 (n_6500), .A2 (n_6495), .A3 (n_6499), .A4 (n_6497));
NAND2_X1 i_6522 (.ZN (n_6458), .A1 (n_6459), .A2 (n_6460));
NAND2_X1 i_6521 (.ZN (n_6457), .A1 (n_6458), .A2 (n_6493));
NAND3_X1 i_6520 (.ZN (n_6456), .A1 (n_6457), .A2 (n_6504), .A3 (n_6503));
INV_X1 i_6519 (.ZN (n_6455), .A (n_6456));
NAND2_X1 i_6518 (.ZN (n_6454), .A1 (n_6504), .A2 (n_6503));
INV_X1 i_6517 (.ZN (n_6453), .A (n_6457));
NAND2_X1 i_6516 (.ZN (n_6452), .A1 (B_imm[21]), .A2 (A_imm[8]));
OAI22_X1 i_6515 (.ZN (n_6451), .A1 (n_8859), .A2 (n_8573), .B1 (n_8909), .B2 (n_8926));
NAND2_X1 i_6514 (.ZN (n_6450), .A1 (A_imm[18]), .A2 (B_imm[10]));
NAND4_X1 i_6513 (.ZN (n_6449), .A1 (A_imm[21]), .A2 (B_imm[17]), .A3 (B_imm[7]), .A4 (A_imm[11]));
NAND2_X1 i_6512 (.ZN (n_6448), .A1 (n_6449), .A2 (n_6450));
NAND2_X1 i_6511 (.ZN (n_6447), .A1 (n_6448), .A2 (n_6451));
NAND2_X1 i_6510 (.ZN (n_6446), .A1 (n_6447), .A2 (n_6452));
NAND2_X1 i_6509 (.ZN (n_6445), .A1 (B_imm[22]), .A2 (A_imm[7]));
NAND4_X1 i_6508 (.ZN (n_6444), .A1 (n_6448), .A2 (n_6451), .A3 (B_imm[21]), .A4 (A_imm[8]));
NAND2_X1 i_6507 (.ZN (n_6443), .A1 (n_6444), .A2 (n_6445));
NAND2_X1 i_6506 (.ZN (n_6442), .A1 (n_6443), .A2 (n_6446));
OAI21_X1 i_6505 (.ZN (n_6441), .A (n_6442), .B1 (n_7913), .B2 (n_8858));
NAND2_X1 i_6504 (.ZN (n_6440), .A1 (A_imm[29]), .A2 (B_imm[1]));
NAND4_X1 i_6503 (.ZN (n_6439), .A1 (n_6443), .A2 (B_imm[14]), .A3 (A_imm[16]), .A4 (n_6446));
NAND2_X1 i_6502 (.ZN (n_6438), .A1 (n_6439), .A2 (n_6440));
NAND2_X1 i_6501 (.ZN (n_6437), .A1 (n_6438), .A2 (n_6441));
INV_X1 i_6500 (.ZN (n_6436), .A (n_6437));
INV_X1 i_6499 (.ZN (n_6435), .A (n_6810));
OAI21_X1 i_6498 (.ZN (n_6434), .A (n_6808), .B1 (n_6435), .B2 (n_6806));
NAND3_X1 i_6497 (.ZN (n_6433), .A1 (n_6810), .A2 (n_6809), .A3 (n_6807));
NAND2_X1 i_6496 (.ZN (n_6432), .A1 (n_6434), .A2 (n_6433));
NAND2_X1 i_6495 (.ZN (n_6431), .A1 (n_6436), .A2 (n_6432));
NAND3_X1 i_6494 (.ZN (n_6430), .A1 (n_6437), .A2 (n_6434), .A3 (n_6433));
NAND2_X1 i_6493 (.ZN (n_6429), .A1 (n_6536), .A2 (n_6534));
NAND2_X1 i_6492 (.ZN (n_6428), .A1 (n_6429), .A2 (n_6527));
NAND3_X1 i_6491 (.ZN (n_6427), .A1 (n_6536), .A2 (n_6535), .A3 (n_6534));
NAND2_X1 i_6490 (.ZN (n_6426), .A1 (n_6428), .A2 (n_6427));
NAND2_X1 i_6489 (.ZN (n_6425), .A1 (n_6430), .A2 (n_6426));
NAND2_X1 i_6488 (.ZN (n_6424), .A1 (n_6425), .A2 (n_6431));
NAND2_X1 i_6487 (.ZN (n_6423), .A1 (A_imm[30]), .A2 (B_imm[1]));
NAND2_X1 i_6486 (.ZN (n_6422), .A1 (n_6834), .A2 (n_6832));
NAND3_X1 i_6485 (.ZN (n_6421), .A1 (n_6422), .A2 (B_imm[28]), .A3 (A_imm[3]));
NAND3_X1 i_6484 (.ZN (n_6420), .A1 (n_6834), .A2 (n_6833), .A3 (n_6832));
NAND3_X1 i_6483 (.ZN (n_6419), .A1 (n_6423), .A2 (n_6421), .A3 (n_6420));
NAND2_X1 i_6482 (.ZN (n_6418), .A1 (n_6421), .A2 (n_6420));
NAND3_X1 i_6481 (.ZN (n_6417), .A1 (n_6418), .A2 (B_imm[1]), .A3 (A_imm[30]));
INV_X1 i_6480 (.ZN (n_6416), .A (n_6417));
NAND2_X1 i_6479 (.ZN (n_6415), .A1 (B_imm[20]), .A2 (A_imm[9]));
OAI21_X1 i_6478 (.ZN (n_6414), .A (n_6415), .B1 (n_9021), .B2 (n_6836));
NAND2_X1 i_6477 (.ZN (n_6413), .A1 (B_imm[26]), .A2 (A_imm[3]));
NAND4_X1 i_6476 (.ZN (n_6412), .A1 (B_imm[28]), .A2 (B_imm[20]), .A3 (A_imm[9]), .A4 (A_imm[1]));
NAND2_X1 i_6475 (.ZN (n_6411), .A1 (n_6412), .A2 (n_6413));
NAND4_X1 i_6474 (.ZN (n_6410), .A1 (n_6411), .A2 (B_imm[30]), .A3 (A_imm[0]), .A4 (n_6414));
AOI22_X1 i_6473 (.ZN (n_6409), .A1 (n_6411), .A2 (n_6414), .B1 (B_imm[30]), .B2 (A_imm[0]));
NAND2_X1 i_6472 (.ZN (n_6408), .A1 (n_6815), .A2 (n_6813));
XNOR2_X1 i_6471 (.ZN (n_6407), .A (n_6408), .B (n_6814));
OAI21_X1 i_6470 (.ZN (n_6406), .A (n_6410), .B1 (n_6409), .B2 (n_6407));
OAI21_X1 i_6469 (.ZN (n_6405), .A (n_6419), .B1 (n_6416), .B2 (n_6406));
INV_X1 i_6468 (.ZN (n_6404), .A (n_6405));
NAND2_X1 i_6467 (.ZN (n_6403), .A1 (n_6424), .A2 (n_6404));
NAND3_X1 i_6466 (.ZN (n_6402), .A1 (n_6425), .A2 (n_6405), .A3 (n_6431));
AOI21_X1 i_6465 (.ZN (n_6401), .A (n_6516), .B1 (n_6521), .B2 (n_6528));
NAND3_X1 i_6464 (.ZN (n_6400), .A1 (n_6521), .A2 (n_6528), .A3 (n_6516));
INV_X1 i_6463 (.ZN (n_6399), .A (n_6400));
NOR2_X1 i_6462 (.ZN (n_6398), .A1 (n_6401), .A2 (n_6399));
NAND2_X1 i_6461 (.ZN (n_6397), .A1 (n_6402), .A2 (n_6398));
AOI22_X1 i_6460 (.ZN (n_6396), .A1 (n_6454), .A2 (n_6453), .B1 (n_6397), .B2 (n_6403));
OAI21_X2 i_6459 (.ZN (n_6395), .A (n_6547), .B1 (n_6396), .B2 (n_6455));
INV_X1 i_6458 (.ZN (n_6394), .A (n_6547));
NAND2_X1 i_6457 (.ZN (n_6393), .A1 (n_6454), .A2 (n_6453));
NAND2_X1 i_6456 (.ZN (n_6392), .A1 (n_6397), .A2 (n_6403));
NAND2_X1 i_6455 (.ZN (n_6391), .A1 (n_6393), .A2 (n_6392));
NAND3_X1 i_6454 (.ZN (n_6390), .A1 (n_6391), .A2 (n_6394), .A3 (n_6456));
INV_X1 i_6453 (.ZN (n_6389), .A (n_6795));
INV_X1 i_6452 (.ZN (n_6388), .A (n_6800));
NAND3_X1 i_6451 (.ZN (n_6387), .A1 (n_6388), .A2 (n_6840), .A3 (n_6839));
NAND2_X1 i_6450 (.ZN (n_6386), .A1 (n_6387), .A2 (n_6799));
XNOR2_X2 i_6449 (.ZN (n_6385), .A (n_6386), .B (n_6389));
NAND2_X1 i_6448 (.ZN (n_6384), .A1 (n_6390), .A2 (n_6385));
NAND2_X1 i_6447 (.ZN (n_6383), .A1 (n_6384), .A2 (n_6395));
NAND2_X1 i_6446 (.ZN (n_6382), .A1 (n_6383), .A2 (n_6596));
NAND3_X2 i_6445 (.ZN (n_6381), .A1 (n_6384), .A2 (n_6597), .A3 (n_6395));
NAND2_X1 i_6444 (.ZN (n_6380), .A1 (n_6514), .A2 (n_6506));
NAND2_X1 i_6443 (.ZN (n_6379), .A1 (B_imm[19]), .A2 (A_imm[13]));
NAND2_X1 i_6442 (.ZN (n_6378), .A1 (B_imm[26]), .A2 (A_imm[6]));
NAND2_X1 i_6441 (.ZN (n_6377), .A1 (n_6379), .A2 (n_6378));
NAND2_X1 i_6440 (.ZN (n_6376), .A1 (B_imm[27]), .A2 (A_imm[5]));
NAND4_X1 i_6439 (.ZN (n_6375), .A1 (B_imm[19]), .A2 (B_imm[26]), .A3 (A_imm[13]), .A4 (A_imm[6]));
NAND2_X1 i_6438 (.ZN (n_6374), .A1 (n_6375), .A2 (n_6376));
NAND2_X1 i_6437 (.ZN (n_6373), .A1 (n_6374), .A2 (n_6377));
NAND2_X1 i_6436 (.ZN (n_6372), .A1 (B_imm[23]), .A2 (A_imm[9]));
NAND2_X1 i_6435 (.ZN (n_6371), .A1 (n_6671), .A2 (n_6668));
NAND2_X1 i_6434 (.ZN (n_6370), .A1 (n_6371), .A2 (n_6672));
NAND2_X1 i_6433 (.ZN (n_6369), .A1 (n_6370), .A2 (n_6372));
NAND2_X1 i_6432 (.ZN (n_6368), .A1 (B_imm[21]), .A2 (A_imm[11]));
NAND4_X1 i_6431 (.ZN (n_6367), .A1 (n_6371), .A2 (B_imm[23]), .A3 (A_imm[9]), .A4 (n_6672));
NAND2_X1 i_6430 (.ZN (n_6366), .A1 (n_6367), .A2 (n_6368));
NAND2_X1 i_6429 (.ZN (n_6365), .A1 (n_6366), .A2 (n_6369));
NAND2_X1 i_6428 (.ZN (n_6364), .A1 (n_6373), .A2 (n_6365));
NAND4_X1 i_6427 (.ZN (n_6363), .A1 (n_6374), .A2 (n_6366), .A3 (n_6377), .A4 (n_6369));
INV_X1 i_6426 (.ZN (n_6362), .A (n_6363));
NAND2_X1 i_6425 (.ZN (n_6361), .A1 (B_imm[14]), .A2 (A_imm[19]));
INV_X1 i_6424 (.ZN (n_6360), .A (n_6361));
OAI21_X1 i_6423 (.ZN (n_6359), .A (n_6364), .B1 (n_6362), .B2 (n_6360));
INV_X1 i_6422 (.ZN (n_6358), .A (n_6359));
NAND2_X1 i_6421 (.ZN (n_6357), .A1 (A_imm[30]), .A2 (B_imm[4]));
NAND2_X1 i_6420 (.ZN (n_6356), .A1 (B_imm[30]), .A2 (A_imm[3]));
NAND2_X1 i_6419 (.ZN (n_6355), .A1 (B_imm[20]), .A2 (A_imm[12]));
NAND2_X1 i_6418 (.ZN (n_6354), .A1 (B_imm[13]), .A2 (A_imm[19]));
NAND2_X1 i_6417 (.ZN (n_6353), .A1 (n_6355), .A2 (n_6354));
NAND2_X1 i_6416 (.ZN (n_6352), .A1 (B_imm[28]), .A2 (A_imm[4]));
INV_X1 i_6415 (.ZN (n_6351), .A (n_6352));
NAND4_X1 i_6414 (.ZN (n_6350), .A1 (B_imm[20]), .A2 (B_imm[13]), .A3 (A_imm[19]), .A4 (A_imm[12]));
INV_X1 i_6413 (.ZN (n_6349), .A (n_6350));
OAI21_X1 i_6412 (.ZN (n_6348), .A (n_6353), .B1 (n_6349), .B2 (n_6351));
NAND2_X1 i_6411 (.ZN (n_6347), .A1 (n_6348), .A2 (n_6356));
NAND2_X1 i_6410 (.ZN (n_6346), .A1 (n_6350), .A2 (n_6352));
NAND4_X1 i_6409 (.ZN (n_6345), .A1 (n_6346), .A2 (B_imm[30]), .A3 (A_imm[3]), .A4 (n_6353));
INV_X1 i_6408 (.ZN (n_6344), .A (n_6345));
NAND2_X1 i_6407 (.ZN (n_6343), .A1 (B_imm[31]), .A2 (A_imm[2]));
INV_X1 i_6406 (.ZN (n_6342), .A (n_6343));
OAI21_X1 i_6405 (.ZN (n_6341), .A (n_6347), .B1 (n_6344), .B2 (n_6342));
NAND2_X1 i_6404 (.ZN (n_6340), .A1 (n_6341), .A2 (n_6357));
OAI21_X1 i_6403 (.ZN (n_6339), .A (n_6343), .B1 (n_6348), .B2 (n_6356));
NAND4_X1 i_6402 (.ZN (n_6338), .A1 (n_6339), .A2 (B_imm[4]), .A3 (A_imm[30]), .A4 (n_6347));
NAND2_X1 i_6401 (.ZN (n_6337), .A1 (n_6338), .A2 (n_6340));
NAND2_X1 i_6400 (.ZN (n_6336), .A1 (n_6337), .A2 (n_6358));
NAND3_X1 i_6399 (.ZN (n_6335), .A1 (n_6340), .A2 (n_6338), .A3 (n_6359));
NAND4_X1 i_6398 (.ZN (n_6334), .A1 (n_6380), .A2 (n_6336), .A3 (n_6511), .A4 (n_6335));
NAND2_X1 i_6397 (.ZN (n_6333), .A1 (n_6380), .A2 (n_6511));
NAND2_X1 i_6396 (.ZN (n_6332), .A1 (n_6336), .A2 (n_6335));
NAND2_X1 i_6395 (.ZN (n_6331), .A1 (n_6333), .A2 (n_6332));
NAND2_X1 i_6394 (.ZN (n_6330), .A1 (n_7506), .A2 (n_7505));
INV_X1 i_6393 (.ZN (n_6329), .A (n_7501));
AOI21_X1 i_6392 (.ZN (n_6328), .A (n_6329), .B1 (n_6330), .B2 (n_7508));
NAND3_X1 i_6391 (.ZN (n_6327), .A1 (n_6330), .A2 (n_7508), .A3 (n_6329));
INV_X1 i_6390 (.ZN (n_6326), .A (n_6327));
NOR2_X2 i_6389 (.ZN (n_6325), .A1 (n_6326), .A2 (n_6328));
NAND3_X1 i_6388 (.ZN (n_6324), .A1 (n_6331), .A2 (n_6334), .A3 (n_6325));
NAND2_X1 i_6387 (.ZN (n_6323), .A1 (n_6331), .A2 (n_6334));
INV_X1 i_6386 (.ZN (n_6322), .A (n_6325));
NAND2_X1 i_6385 (.ZN (n_6321), .A1 (n_6323), .A2 (n_6322));
NAND2_X1 i_6384 (.ZN (n_6320), .A1 (n_6321), .A2 (n_6324));
INV_X1 i_6383 (.ZN (n_6319), .A (n_6320));
NAND2_X1 i_6382 (.ZN (n_6318), .A1 (B_imm[30]), .A2 (A_imm[1]));
NAND2_X1 i_6381 (.ZN (n_6317), .A1 (B_imm[13]), .A2 (A_imm[17]));
NAND2_X1 i_6380 (.ZN (n_6316), .A1 (B_imm[25]), .A2 (A_imm[5]));
NAND2_X1 i_6379 (.ZN (n_6315), .A1 (n_6316), .A2 (n_6317));
NAND2_X1 i_6378 (.ZN (n_6314), .A1 (B_imm[20]), .A2 (A_imm[10]));
NAND4_X1 i_6377 (.ZN (n_6313), .A1 (B_imm[25]), .A2 (B_imm[13]), .A3 (A_imm[17]), .A4 (A_imm[5]));
NAND2_X1 i_6376 (.ZN (n_6312), .A1 (n_6313), .A2 (n_6314));
NAND2_X1 i_6375 (.ZN (n_6311), .A1 (n_6312), .A2 (n_6315));
NAND2_X1 i_6374 (.ZN (n_6310), .A1 (n_6311), .A2 (n_6318));
NAND2_X1 i_6373 (.ZN (n_6309), .A1 (B_imm[31]), .A2 (A_imm[0]));
NAND4_X1 i_6372 (.ZN (n_6308), .A1 (n_6312), .A2 (B_imm[30]), .A3 (A_imm[1]), .A4 (n_6315));
NAND2_X1 i_6371 (.ZN (n_6307), .A1 (n_6308), .A2 (n_6309));
NAND2_X1 i_6370 (.ZN (n_6306), .A1 (A_imm[27]), .A2 (B_imm[4]));
NAND2_X1 i_6369 (.ZN (n_6305), .A1 (B_imm[22]), .A2 (A_imm[8]));
NAND2_X1 i_6368 (.ZN (n_6304), .A1 (B_imm[21]), .A2 (A_imm[9]));
NAND2_X1 i_6367 (.ZN (n_6303), .A1 (n_6305), .A2 (n_6304));
NAND2_X1 i_6366 (.ZN (n_6302), .A1 (B_imm[15]), .A2 (A_imm[15]));
INV_X1 i_6365 (.ZN (n_6301), .A (n_6302));
NAND4_X1 i_6364 (.ZN (n_6300), .A1 (B_imm[22]), .A2 (B_imm[21]), .A3 (A_imm[9]), .A4 (A_imm[8]));
INV_X1 i_6363 (.ZN (n_6299), .A (n_6300));
OAI21_X1 i_6362 (.ZN (n_6298), .A (n_6303), .B1 (n_6299), .B2 (n_6301));
NAND2_X1 i_6361 (.ZN (n_6297), .A1 (n_6298), .A2 (n_6306));
NAND2_X1 i_6360 (.ZN (n_6296), .A1 (B_imm[24]), .A2 (A_imm[6]));
OAI21_X1 i_6359 (.ZN (n_6295), .A (n_6296), .B1 (n_8821), .B2 (n_8644));
NAND2_X1 i_6358 (.ZN (n_6294), .A1 (A_imm[19]), .A2 (B_imm[10]));
OAI21_X1 i_6357 (.ZN (n_6293), .A (n_6294), .B1 (n_8908), .B2 (n_8927));
NAND2_X1 i_6356 (.ZN (n_6292), .A1 (A_imm[22]), .A2 (B_imm[7]));
INV_X1 i_6355 (.ZN (n_6291), .A (n_6292));
NAND4_X1 i_6354 (.ZN (n_6290), .A1 (B_imm[16]), .A2 (A_imm[19]), .A3 (B_imm[10]), .A4 (A_imm[13]));
INV_X1 i_6353 (.ZN (n_6289), .A (n_6290));
OAI21_X1 i_6352 (.ZN (n_6288), .A (n_6293), .B1 (n_6289), .B2 (n_6291));
NAND4_X1 i_6351 (.ZN (n_6287), .A1 (B_imm[23]), .A2 (B_imm[24]), .A3 (A_imm[7]), .A4 (A_imm[6]));
NAND2_X1 i_6350 (.ZN (n_6286), .A1 (n_6287), .A2 (n_6288));
NAND2_X1 i_6349 (.ZN (n_6285), .A1 (n_6286), .A2 (n_6295));
OAI21_X1 i_6348 (.ZN (n_6284), .A (n_6285), .B1 (n_6298), .B2 (n_6306));
NAND4_X1 i_6347 (.ZN (n_6283), .A1 (n_6307), .A2 (n_6284), .A3 (n_6310), .A4 (n_6297));
INV_X1 i_6346 (.ZN (n_6282), .A (n_6309));
INV_X1 i_6345 (.ZN (n_6281), .A (n_6308));
OAI21_X1 i_6344 (.ZN (n_6280), .A (n_6310), .B1 (n_6281), .B2 (n_6282));
INV_X1 i_6343 (.ZN (n_6279), .A (n_6285));
NAND2_X1 i_6342 (.ZN (n_6278), .A1 (n_6300), .A2 (n_6302));
NAND4_X1 i_6341 (.ZN (n_6277), .A1 (n_6278), .A2 (B_imm[4]), .A3 (A_imm[27]), .A4 (n_6303));
INV_X1 i_6340 (.ZN (n_6276), .A (n_6277));
OAI21_X1 i_6339 (.ZN (n_6275), .A (n_6297), .B1 (n_6276), .B2 (n_6279));
NAND2_X1 i_6338 (.ZN (n_6274), .A1 (n_6280), .A2 (n_6275));
AOI21_X1 i_6337 (.ZN (n_6273), .A (n_6368), .B1 (n_6367), .B2 (n_6369));
NAND3_X1 i_6336 (.ZN (n_6272), .A1 (n_6369), .A2 (n_6367), .A3 (n_6368));
INV_X1 i_6335 (.ZN (n_6271), .A (n_6272));
NOR2_X1 i_6334 (.ZN (n_6270), .A1 (n_6271), .A2 (n_6273));
INV_X1 i_6333 (.ZN (n_6269), .A (n_6270));
NAND2_X1 i_6332 (.ZN (n_6268), .A1 (n_6274), .A2 (n_6269));
NAND2_X1 i_6331 (.ZN (n_6267), .A1 (n_6353), .A2 (n_6350));
NAND2_X1 i_6330 (.ZN (n_6266), .A1 (n_6267), .A2 (n_6351));
NAND3_X1 i_6329 (.ZN (n_6265), .A1 (n_6353), .A2 (n_6350), .A3 (n_6352));
NAND2_X1 i_6328 (.ZN (n_6264), .A1 (n_6266), .A2 (n_6265));
INV_X1 i_6327 (.ZN (n_6263), .A (n_6376));
NAND2_X1 i_6326 (.ZN (n_6262), .A1 (n_6377), .A2 (n_6375));
NAND2_X1 i_6325 (.ZN (n_6261), .A1 (n_6262), .A2 (n_6263));
NAND3_X1 i_6324 (.ZN (n_6260), .A1 (n_6377), .A2 (n_6375), .A3 (n_6376));
NAND2_X1 i_6323 (.ZN (n_6259), .A1 (n_6261), .A2 (n_6260));
NAND2_X1 i_6322 (.ZN (n_6258), .A1 (n_6259), .A2 (n_6264));
NAND2_X1 i_6321 (.ZN (n_6257), .A1 (A_imm[30]), .A2 (B_imm[2]));
NAND4_X1 i_6320 (.ZN (n_6256), .A1 (n_6261), .A2 (n_6266), .A3 (n_6265), .A4 (n_6260));
INV_X1 i_6319 (.ZN (n_6255), .A (n_6256));
OAI21_X1 i_6318 (.ZN (n_6254), .A (n_6258), .B1 (n_6255), .B2 (n_6257));
INV_X1 i_6317 (.ZN (n_6253), .A (n_6254));
NAND3_X1 i_6316 (.ZN (n_6252), .A1 (n_6268), .A2 (n_6253), .A3 (n_6283));
INV_X1 i_6315 (.ZN (n_6251), .A (n_6283));
AOI21_X1 i_6314 (.ZN (n_6250), .A (n_6270), .B1 (n_6280), .B2 (n_6275));
OAI21_X1 i_6313 (.ZN (n_6249), .A (n_6254), .B1 (n_6250), .B2 (n_6251));
NAND2_X1 i_6312 (.ZN (n_6248), .A1 (n_8159), .A2 (n_8157));
NAND3_X1 i_6311 (.ZN (n_6247), .A1 (n_6248), .A2 (B_imm[10]), .A3 (A_imm[23]));
NAND3_X1 i_6310 (.ZN (n_6246), .A1 (n_8159), .A2 (n_8158), .A3 (n_8157));
NAND2_X1 i_6309 (.ZN (n_6245), .A1 (n_6247), .A2 (n_6246));
NAND3_X1 i_6308 (.ZN (n_6244), .A1 (n_6245), .A2 (B_imm[4]), .A3 (A_imm[29]));
OAI211_X1 i_6307 (.ZN (n_6243), .A (n_6247), .B (n_6246), .C1 (n_8994), .C2 (n_6577));
INV_X1 i_6306 (.ZN (n_6242), .A (n_8151));
OAI21_X1 i_6305 (.ZN (n_6241), .A (n_8149), .B1 (n_6242), .B2 (n_8147));
NAND3_X1 i_6304 (.ZN (n_6240), .A1 (n_8151), .A2 (n_8150), .A3 (n_8148));
NAND4_X1 i_6303 (.ZN (n_6239), .A1 (n_6243), .A2 (n_6244), .A3 (n_6241), .A4 (n_6240));
INV_X1 i_6302 (.ZN (n_6238), .A (n_6244));
INV_X1 i_6301 (.ZN (n_6237), .A (n_6243));
NAND2_X1 i_6300 (.ZN (n_6236), .A1 (n_6241), .A2 (n_6240));
OAI21_X1 i_6299 (.ZN (n_6235), .A (n_6236), .B1 (n_6237), .B2 (n_6238));
NAND2_X1 i_6298 (.ZN (n_6234), .A1 (n_6235), .A2 (n_6239));
NAND3_X1 i_6297 (.ZN (n_6233), .A1 (n_6252), .A2 (n_6249), .A3 (n_6234));
AOI21_X1 i_6296 (.ZN (n_6232), .A (n_6234), .B1 (n_6249), .B2 (n_6252));
INV_X1 i_6295 (.ZN (n_6231), .A (n_6232));
NAND2_X1 i_6294 (.ZN (n_6230), .A1 (A_imm[28]), .A2 (B_imm[3]));
NAND2_X1 i_6293 (.ZN (n_6229), .A1 (B_imm[12]), .A2 (A_imm[18]));
OAI21_X1 i_6292 (.ZN (n_6228), .A (n_6229), .B1 (n_8849), .B2 (n_8892));
NAND2_X1 i_6291 (.ZN (n_6227), .A1 (A_imm[25]), .A2 (B_imm[5]));
INV_X1 i_6290 (.ZN (n_6226), .A (n_6227));
NAND4_X1 i_6289 (.ZN (n_6225), .A1 (B_imm[11]), .A2 (B_imm[12]), .A3 (A_imm[19]), .A4 (A_imm[18]));
INV_X1 i_6288 (.ZN (n_6224), .A (n_6225));
OAI21_X1 i_6287 (.ZN (n_6223), .A (n_6228), .B1 (n_6224), .B2 (n_6226));
NAND2_X1 i_6286 (.ZN (n_6222), .A1 (n_6223), .A2 (n_6230));
NAND2_X1 i_6285 (.ZN (n_6221), .A1 (A_imm[26]), .A2 (B_imm[4]));
OAI21_X1 i_6284 (.ZN (n_6220), .A (n_6221), .B1 (n_8423), .B2 (n_8752));
NAND2_X1 i_6283 (.ZN (n_6219), .A1 (B_imm[9]), .A2 (A_imm[21]));
INV_X1 i_6282 (.ZN (n_6218), .A (n_6219));
NAND4_X1 i_6281 (.ZN (n_6217), .A1 (B_imm[18]), .A2 (A_imm[26]), .A3 (B_imm[4]), .A4 (A_imm[12]));
INV_X1 i_6280 (.ZN (n_6216), .A (n_6217));
OAI21_X1 i_6279 (.ZN (n_6215), .A (n_6220), .B1 (n_6216), .B2 (n_6218));
OAI21_X1 i_6278 (.ZN (n_6214), .A (n_6215), .B1 (n_6223), .B2 (n_6230));
NAND2_X1 i_6277 (.ZN (n_6213), .A1 (n_6214), .A2 (n_6222));
AOI21_X1 i_6276 (.ZN (n_6212), .A (n_7527), .B1 (n_7528), .B2 (n_7525));
INV_X1 i_6275 (.ZN (n_6211), .A (n_6212));
NAND3_X1 i_6274 (.ZN (n_6210), .A1 (n_7528), .A2 (n_7527), .A3 (n_7525));
NAND2_X1 i_6273 (.ZN (n_6209), .A1 (n_6211), .A2 (n_6210));
INV_X1 i_6272 (.ZN (n_6208), .A (n_6209));
NAND2_X1 i_6271 (.ZN (n_6207), .A1 (n_6213), .A2 (n_6208));
NAND3_X1 i_6270 (.ZN (n_6206), .A1 (n_6209), .A2 (n_6214), .A3 (n_6222));
NAND2_X1 i_6269 (.ZN (n_6205), .A1 (n_6207), .A2 (n_6206));
AOI21_X1 i_6268 (.ZN (n_6204), .A (n_7521), .B1 (n_7522), .B2 (n_7520));
NAND3_X1 i_6267 (.ZN (n_6203), .A1 (n_7522), .A2 (n_7521), .A3 (n_7520));
INV_X1 i_6266 (.ZN (n_6202), .A (n_6203));
NOR2_X2 i_6265 (.ZN (n_6201), .A1 (n_6204), .A2 (n_6202));
NAND2_X1 i_6264 (.ZN (n_6200), .A1 (n_6205), .A2 (n_6201));
INV_X1 i_6263 (.ZN (n_6199), .A (n_6201));
NAND3_X1 i_6262 (.ZN (n_6198), .A1 (n_6207), .A2 (n_6199), .A3 (n_6206));
AOI21_X1 i_6261 (.ZN (n_6197), .A (n_6269), .B1 (n_6283), .B2 (n_6274));
INV_X1 i_6260 (.ZN (n_6196), .A (n_6197));
NAND3_X1 i_6259 (.ZN (n_6195), .A1 (n_6274), .A2 (n_6283), .A3 (n_6269));
NAND4_X1 i_6258 (.ZN (n_6194), .A1 (n_6196), .A2 (n_6200), .A3 (n_6198), .A4 (n_6195));
INV_X1 i_6257 (.ZN (n_6193), .A (n_6194));
NAND2_X1 i_6256 (.ZN (n_6192), .A1 (n_6200), .A2 (n_6198));
NAND2_X1 i_6255 (.ZN (n_6191), .A1 (n_6196), .A2 (n_6195));
INV_X1 i_6254 (.ZN (n_6190), .A (n_6215));
NAND2_X1 i_6253 (.ZN (n_6189), .A1 (n_6225), .A2 (n_6227));
NAND4_X1 i_6252 (.ZN (n_6188), .A1 (n_6189), .A2 (B_imm[3]), .A3 (A_imm[28]), .A4 (n_6228));
NAND2_X1 i_6251 (.ZN (n_6187), .A1 (n_6222), .A2 (n_6188));
NAND2_X1 i_6250 (.ZN (n_6186), .A1 (n_6187), .A2 (n_6190));
NAND3_X1 i_6249 (.ZN (n_6185), .A1 (n_6222), .A2 (n_6188), .A3 (n_6215));
NAND2_X1 i_6248 (.ZN (n_6184), .A1 (n_6186), .A2 (n_6185));
NAND2_X1 i_6247 (.ZN (n_6183), .A1 (B_imm[19]), .A2 (A_imm[10]));
OAI21_X1 i_6246 (.ZN (n_6182), .A (n_6183), .B1 (n_9003), .B2 (n_6677));
NAND2_X1 i_6245 (.ZN (n_6181), .A1 (A_imm[12]), .A2 (B_imm[16]));
OAI21_X1 i_6244 (.ZN (n_6180), .A (n_6181), .B1 (n_8232), .B2 (n_8906));
NAND2_X1 i_6243 (.ZN (n_6179), .A1 (B_imm[8]), .A2 (A_imm[20]));
NAND4_X1 i_6242 (.ZN (n_6178), .A1 (B_imm[6]), .A2 (A_imm[12]), .A3 (B_imm[16]), .A4 (A_imm[22]));
NAND2_X1 i_6241 (.ZN (n_6177), .A1 (n_6178), .A2 (n_6179));
NAND2_X1 i_6240 (.ZN (n_6176), .A1 (n_6177), .A2 (n_6180));
NAND4_X1 i_6239 (.ZN (n_6175), .A1 (B_imm[27]), .A2 (B_imm[19]), .A3 (A_imm[10]), .A4 (A_imm[2]));
NAND2_X1 i_6238 (.ZN (n_6174), .A1 (n_6175), .A2 (n_6176));
AOI21_X1 i_6237 (.ZN (n_6173), .A (n_6540), .B1 (n_6541), .B2 (n_6539));
NAND3_X1 i_6236 (.ZN (n_6172), .A1 (n_6541), .A2 (n_6540), .A3 (n_6539));
INV_X1 i_6235 (.ZN (n_6171), .A (n_6172));
OAI211_X1 i_6234 (.ZN (n_6170), .A (n_6174), .B (n_6182), .C1 (n_6173), .C2 (n_6171));
INV_X1 i_6233 (.ZN (n_6169), .A (n_6176));
INV_X1 i_6232 (.ZN (n_6168), .A (n_6175));
OAI21_X1 i_6231 (.ZN (n_6167), .A (n_6182), .B1 (n_6168), .B2 (n_6169));
NOR2_X1 i_6230 (.ZN (n_6166), .A1 (n_6171), .A2 (n_6173));
NAND2_X1 i_6229 (.ZN (n_6165), .A1 (n_6167), .A2 (n_6166));
INV_X1 i_6228 (.ZN (n_6164), .A (n_6228));
OAI21_X1 i_6227 (.ZN (n_6163), .A (n_6226), .B1 (n_6164), .B2 (n_6224));
NAND3_X1 i_6226 (.ZN (n_6162), .A1 (n_6228), .A2 (n_6227), .A3 (n_6225));
NAND2_X1 i_6225 (.ZN (n_6161), .A1 (n_6163), .A2 (n_6162));
NAND2_X1 i_6224 (.ZN (n_6160), .A1 (n_6165), .A2 (n_6161));
NAND2_X1 i_6223 (.ZN (n_6159), .A1 (n_6160), .A2 (n_6170));
NAND2_X1 i_6222 (.ZN (n_6158), .A1 (n_6159), .A2 (n_6184));
AOI22_X1 i_6221 (.ZN (n_6157), .A1 (n_6278), .A2 (n_6303), .B1 (A_imm[27]), .B2 (B_imm[4]));
OAI21_X1 i_6220 (.ZN (n_6156), .A (n_6279), .B1 (n_6276), .B2 (n_6157));
OAI21_X1 i_6219 (.ZN (n_6155), .A (n_6156), .B1 (n_6157), .B2 (n_6284));
NAND4_X1 i_6218 (.ZN (n_6154), .A1 (n_6160), .A2 (n_6186), .A3 (n_6185), .A4 (n_6170));
NAND2_X1 i_6217 (.ZN (n_6153), .A1 (n_6154), .A2 (n_6155));
AOI22_X1 i_6216 (.ZN (n_6152), .A1 (n_6191), .A2 (n_6192), .B1 (n_6158), .B2 (n_6153));
OAI211_X1 i_6215 (.ZN (n_6151), .A (n_6233), .B (n_6231), .C1 (n_6152), .C2 (n_6193));
INV_X1 i_6214 (.ZN (n_6150), .A (n_6151));
INV_X1 i_6213 (.ZN (n_6149), .A (n_6233));
INV_X1 i_6212 (.ZN (n_6148), .A (n_6195));
OAI21_X1 i_6211 (.ZN (n_6147), .A (n_6192), .B1 (n_6148), .B2 (n_6197));
NAND2_X1 i_6210 (.ZN (n_6146), .A1 (n_6153), .A2 (n_6158));
NAND2_X1 i_6209 (.ZN (n_6145), .A1 (n_6147), .A2 (n_6146));
OAI211_X1 i_6208 (.ZN (n_6144), .A (n_6145), .B (n_6194), .C1 (n_6149), .C2 (n_6232));
AOI22_X1 i_6207 (.ZN (n_6143), .A1 (n_6346), .A2 (n_6353), .B1 (B_imm[30]), .B2 (A_imm[3]));
OAI21_X1 i_6206 (.ZN (n_6142), .A (n_6342), .B1 (n_6344), .B2 (n_6143));
NAND3_X1 i_6205 (.ZN (n_6141), .A1 (n_6347), .A2 (n_6345), .A3 (n_6343));
NAND2_X1 i_6204 (.ZN (n_6140), .A1 (n_6207), .A2 (n_6199));
NAND4_X1 i_6203 (.ZN (n_6139), .A1 (n_6140), .A2 (n_6206), .A3 (n_6142), .A4 (n_6141));
NAND2_X1 i_6202 (.ZN (n_6138), .A1 (n_6142), .A2 (n_6141));
NAND2_X1 i_6201 (.ZN (n_6137), .A1 (n_6140), .A2 (n_6206));
NAND2_X1 i_6200 (.ZN (n_6136), .A1 (n_6137), .A2 (n_6138));
NAND2_X1 i_6199 (.ZN (n_6135), .A1 (n_6136), .A2 (n_6139));
INV_X1 i_6198 (.ZN (n_6134), .A (n_6364));
OAI21_X1 i_6197 (.ZN (n_6133), .A (n_6360), .B1 (n_6134), .B2 (n_6362));
NAND3_X1 i_6196 (.ZN (n_6132), .A1 (n_6364), .A2 (n_6363), .A3 (n_6361));
NAND3_X1 i_6195 (.ZN (n_6131), .A1 (n_6135), .A2 (n_6133), .A3 (n_6132));
NAND2_X1 i_6194 (.ZN (n_6130), .A1 (n_6133), .A2 (n_6132));
NAND3_X1 i_6193 (.ZN (n_6129), .A1 (n_6136), .A2 (n_6139), .A3 (n_6130));
NAND2_X1 i_6192 (.ZN (n_6128), .A1 (n_6131), .A2 (n_6129));
INV_X1 i_6191 (.ZN (n_6127), .A (n_6128));
NAND2_X2 i_6190 (.ZN (n_6126), .A1 (n_6144), .A2 (n_6127));
INV_X1 i_6189 (.ZN (n_6125), .A (n_6126));
OAI21_X2 i_6188 (.ZN (n_6124), .A (n_6319), .B1 (n_6125), .B2 (n_6150));
NAND3_X1 i_6187 (.ZN (n_6123), .A1 (n_6126), .A2 (n_6320), .A3 (n_6151));
NAND2_X1 i_6186 (.ZN (n_6122), .A1 (n_6252), .A2 (n_6234));
NAND2_X1 i_6185 (.ZN (n_6121), .A1 (n_6139), .A2 (n_6130));
NAND4_X1 i_6184 (.ZN (n_6120), .A1 (n_6122), .A2 (n_6121), .A3 (n_6249), .A4 (n_6136));
NAND2_X1 i_6183 (.ZN (n_6119), .A1 (n_6122), .A2 (n_6249));
NAND2_X1 i_6182 (.ZN (n_6118), .A1 (n_6121), .A2 (n_6136));
NAND2_X1 i_6181 (.ZN (n_6117), .A1 (n_6119), .A2 (n_6118));
AOI21_X1 i_6180 (.ZN (n_6116), .A (n_8111), .B1 (n_8120), .B2 (n_8118));
NAND3_X1 i_6179 (.ZN (n_6115), .A1 (n_8120), .A2 (n_8118), .A3 (n_8111));
INV_X1 i_6178 (.ZN (n_6114), .A (n_6115));
INV_X1 i_6177 (.ZN (n_6113), .A (n_8146));
NAND2_X1 i_6176 (.ZN (n_6112), .A1 (n_8154), .A2 (n_8153));
NAND2_X1 i_6175 (.ZN (n_6111), .A1 (n_6112), .A2 (n_6113));
NAND3_X1 i_6174 (.ZN (n_6110), .A1 (n_8154), .A2 (n_8153), .A3 (n_8146));
NAND2_X1 i_6173 (.ZN (n_6109), .A1 (n_6111), .A2 (n_6110));
OAI21_X1 i_6172 (.ZN (n_6108), .A (n_6109), .B1 (n_6114), .B2 (n_6116));
INV_X1 i_6171 (.ZN (n_6107), .A (n_6116));
NAND4_X1 i_6170 (.ZN (n_6106), .A1 (n_6107), .A2 (n_6115), .A3 (n_6111), .A4 (n_6110));
NAND2_X1 i_6169 (.ZN (n_6105), .A1 (n_6106), .A2 (n_6108));
OAI21_X1 i_6168 (.ZN (n_6104), .A (n_6243), .B1 (n_6238), .B2 (n_6236));
INV_X1 i_6167 (.ZN (n_6103), .A (n_6104));
XNOR2_X2 i_6166 (.ZN (n_6102), .A (n_6105), .B (n_6103));
NAND3_X1 i_6165 (.ZN (n_6101), .A1 (n_6117), .A2 (n_6120), .A3 (n_6102));
NAND2_X1 i_6164 (.ZN (n_6100), .A1 (n_6117), .A2 (n_6120));
INV_X1 i_6163 (.ZN (n_6099), .A (n_6102));
NAND2_X1 i_6162 (.ZN (n_6098), .A1 (n_6100), .A2 (n_6099));
NAND2_X1 i_6161 (.ZN (n_6097), .A1 (n_6098), .A2 (n_6101));
INV_X1 i_6160 (.ZN (n_6096), .A (n_6097));
NAND2_X1 i_6159 (.ZN (n_6095), .A1 (n_6123), .A2 (n_6096));
NAND2_X2 i_6158 (.ZN (n_6094), .A1 (n_6095), .A2 (n_6124));
NAND2_X2 i_6157 (.ZN (n_6093), .A1 (n_6094), .A2 (n_6381));
NAND2_X2 i_6156 (.ZN (n_6092), .A1 (n_6093), .A2 (n_6382));
NAND2_X2 i_6155 (.ZN (n_6091), .A1 (n_6092), .A2 (n_6601));
AOI21_X2 i_6154 (.ZN (n_6090), .A (n_6766), .B1 (n_6091), .B2 (n_6602));
INV_X2 i_6153 (.ZN (n_6089), .A (n_6090));
NAND3_X2 i_6152 (.ZN (n_6088), .A1 (n_6091), .A2 (n_6766), .A3 (n_6602));
NAND3_X1 i_6151 (.ZN (n_6087), .A1 (n_8196), .A2 (n_8198), .A3 (n_8234));
OAI21_X1 i_6150 (.ZN (n_6086), .A (n_8209), .B1 (n_8197), .B2 (n_8235));
NAND2_X1 i_6149 (.ZN (n_6085), .A1 (n_6086), .A2 (n_6087));
INV_X1 i_6148 (.ZN (n_6084), .A (n_6085));
INV_X1 i_6147 (.ZN (n_6083), .A (n_6338));
OAI21_X1 i_6146 (.ZN (n_6082), .A (n_6340), .B1 (n_6083), .B2 (n_6358));
NAND2_X1 i_6145 (.ZN (n_6081), .A1 (n_8257), .A2 (n_8260));
NAND2_X1 i_6144 (.ZN (n_6080), .A1 (n_6081), .A2 (n_8250));
INV_X1 i_6143 (.ZN (n_6079), .A (n_8250));
NAND3_X1 i_6142 (.ZN (n_6078), .A1 (n_6079), .A2 (n_8260), .A3 (n_8257));
NAND2_X1 i_6141 (.ZN (n_6077), .A1 (n_6080), .A2 (n_6078));
NAND2_X1 i_6140 (.ZN (n_6076), .A1 (n_6082), .A2 (n_6077));
INV_X1 i_6139 (.ZN (n_6075), .A (n_6077));
OAI211_X1 i_6138 (.ZN (n_6074), .A (n_6075), .B (n_6340), .C1 (n_6083), .C2 (n_6358));
NAND2_X1 i_6137 (.ZN (n_6073), .A1 (n_6108), .A2 (n_6104));
NAND2_X1 i_6136 (.ZN (n_6072), .A1 (n_6073), .A2 (n_6106));
NAND2_X1 i_6135 (.ZN (n_6071), .A1 (n_6072), .A2 (n_6074));
INV_X1 i_6134 (.ZN (n_6070), .A (n_8211));
NAND2_X1 i_6133 (.ZN (n_6069), .A1 (n_8217), .A2 (n_8216));
NAND2_X1 i_6132 (.ZN (n_6068), .A1 (n_6069), .A2 (n_6070));
NAND3_X1 i_6131 (.ZN (n_6067), .A1 (n_8217), .A2 (n_8216), .A3 (n_8211));
NAND4_X1 i_6130 (.ZN (n_6066), .A1 (n_6071), .A2 (n_6076), .A3 (n_6068), .A4 (n_6067));
NAND2_X1 i_6129 (.ZN (n_6065), .A1 (n_6071), .A2 (n_6076));
NAND2_X1 i_6128 (.ZN (n_6064), .A1 (n_6068), .A2 (n_6067));
NAND2_X1 i_6127 (.ZN (n_6063), .A1 (n_6065), .A2 (n_6064));
OAI21_X2 i_6126 (.ZN (n_6062), .A (n_6702), .B1 (n_6704), .B2 (n_6696));
NAND2_X1 i_6125 (.ZN (n_6061), .A1 (n_6062), .A2 (n_6063));
NAND3_X1 i_6124 (.ZN (n_6060), .A1 (n_6061), .A2 (n_6084), .A3 (n_6066));
AOI21_X1 i_6123 (.ZN (n_6059), .A (n_6084), .B1 (n_6061), .B2 (n_6066));
INV_X1 i_6122 (.ZN (n_6058), .A (n_6059));
NAND3_X1 i_6121 (.ZN (n_6057), .A1 (n_8079), .A2 (n_8078), .A3 (n_8073));
INV_X1 i_6120 (.ZN (n_6056), .A (n_8073));
NAND2_X1 i_6119 (.ZN (n_6055), .A1 (n_8079), .A2 (n_8078));
NAND2_X1 i_6118 (.ZN (n_6054), .A1 (n_6055), .A2 (n_6056));
NAND2_X1 i_6117 (.ZN (n_6053), .A1 (n_6054), .A2 (n_6057));
NAND3_X1 i_6116 (.ZN (n_6052), .A1 (n_6058), .A2 (n_6060), .A3 (n_6053));
INV_X1 i_6115 (.ZN (n_6051), .A (n_6060));
INV_X1 i_6114 (.ZN (n_6050), .A (n_6053));
OAI21_X1 i_6113 (.ZN (n_6049), .A (n_6050), .B1 (n_6051), .B2 (n_6059));
NAND2_X1 i_6112 (.ZN (n_6048), .A1 (n_7555), .A2 (n_7558));
NAND3_X1 i_6111 (.ZN (n_6047), .A1 (n_6048), .A2 (n_7497), .A3 (n_7489));
NAND3_X1 i_6110 (.ZN (n_6046), .A1 (n_7488), .A2 (n_7558), .A3 (n_7555));
NAND2_X1 i_6109 (.ZN (n_6045), .A1 (n_6047), .A2 (n_6046));
NAND3_X2 i_6108 (.ZN (n_6044), .A1 (n_6049), .A2 (n_6052), .A3 (n_6045));
AOI21_X1 i_6107 (.ZN (n_6043), .A (n_6045), .B1 (n_6049), .B2 (n_6052));
INV_X2 i_6106 (.ZN (n_6042), .A (n_6043));
NAND3_X1 i_6105 (.ZN (n_6041), .A1 (n_6062), .A2 (n_6066), .A3 (n_6063));
INV_X1 i_6104 (.ZN (n_6040), .A (n_6062));
NAND2_X1 i_6103 (.ZN (n_6039), .A1 (n_6063), .A2 (n_6066));
NAND2_X1 i_6102 (.ZN (n_6038), .A1 (n_6039), .A2 (n_6040));
NAND3_X1 i_6101 (.ZN (n_6037), .A1 (n_6076), .A2 (n_6074), .A3 (n_6072));
INV_X1 i_6100 (.ZN (n_6036), .A (n_6072));
NAND2_X1 i_6099 (.ZN (n_6035), .A1 (n_6076), .A2 (n_6074));
NAND2_X1 i_6098 (.ZN (n_6034), .A1 (n_6035), .A2 (n_6036));
NAND2_X1 i_6097 (.ZN (n_6033), .A1 (n_6034), .A2 (n_6037));
NAND2_X1 i_6096 (.ZN (n_6032), .A1 (n_6334), .A2 (n_6325));
NAND2_X1 i_6095 (.ZN (n_6031), .A1 (n_6032), .A2 (n_6331));
NAND2_X1 i_6094 (.ZN (n_6030), .A1 (n_6031), .A2 (n_6033));
NAND4_X1 i_6093 (.ZN (n_6029), .A1 (n_6032), .A2 (n_6331), .A3 (n_6037), .A4 (n_6034));
NAND2_X1 i_6092 (.ZN (n_6028), .A1 (n_6120), .A2 (n_6102));
NAND2_X1 i_6091 (.ZN (n_6027), .A1 (n_6028), .A2 (n_6117));
NAND2_X1 i_6090 (.ZN (n_6026), .A1 (n_6027), .A2 (n_6029));
NAND2_X1 i_6089 (.ZN (n_6025), .A1 (n_6026), .A2 (n_6030));
NAND3_X1 i_6088 (.ZN (n_6024), .A1 (n_6025), .A2 (n_6041), .A3 (n_6038));
NAND2_X1 i_6087 (.ZN (n_6023), .A1 (n_6038), .A2 (n_6041));
NAND3_X2 i_6086 (.ZN (n_6022), .A1 (n_6023), .A2 (n_6030), .A3 (n_6026));
NAND3_X1 i_6085 (.ZN (n_6021), .A1 (n_6861), .A2 (n_6859), .A3 (n_6854));
INV_X1 i_6084 (.ZN (n_6020), .A (n_6854));
NAND2_X1 i_6083 (.ZN (n_6019), .A1 (n_6861), .A2 (n_6859));
NAND2_X1 i_6082 (.ZN (n_6018), .A1 (n_6019), .A2 (n_6020));
NAND3_X1 i_6081 (.ZN (n_6017), .A1 (n_6022), .A2 (n_6018), .A3 (n_6021));
NAND2_X1 i_6080 (.ZN (n_6016), .A1 (n_6017), .A2 (n_6024));
NAND3_X1 i_6079 (.ZN (n_6015), .A1 (n_6042), .A2 (n_6044), .A3 (n_6016));
INV_X1 i_6078 (.ZN (n_6014), .A (n_6044));
INV_X1 i_6077 (.ZN (n_6013), .A (n_6016));
OAI21_X1 i_6076 (.ZN (n_6012), .A (n_6013), .B1 (n_6014), .B2 (n_6043));
NAND2_X1 i_6075 (.ZN (n_6011), .A1 (n_6012), .A2 (n_6015));
NAND3_X1 i_6074 (.ZN (n_6010), .A1 (n_6089), .A2 (n_6088), .A3 (n_6011));
AOI21_X1 i_6073 (.ZN (n_6009), .A (n_6011), .B1 (n_6089), .B2 (n_6088));
INV_X1 i_6072 (.ZN (n_6008), .A (n_6009));
NAND2_X1 i_6071 (.ZN (n_6007), .A1 (n_6018), .A2 (n_6021));
NAND3_X1 i_6070 (.ZN (n_6006), .A1 (n_6007), .A2 (n_6024), .A3 (n_6022));
NAND2_X1 i_6069 (.ZN (n_6005), .A1 (n_6024), .A2 (n_6022));
NAND3_X1 i_6068 (.ZN (n_6004), .A1 (n_6005), .A2 (n_6021), .A3 (n_6018));
NAND2_X1 i_6067 (.ZN (n_6003), .A1 (n_6004), .A2 (n_6006));
NAND3_X1 i_6066 (.ZN (n_6002), .A1 (n_6610), .A2 (n_6613), .A3 (n_6606));
NAND2_X1 i_6065 (.ZN (n_6001), .A1 (n_6613), .A2 (n_6610));
NAND2_X1 i_6064 (.ZN (n_6000), .A1 (n_6001), .A2 (n_6605));
NAND3_X1 i_6063 (.ZN (n_5999), .A1 (n_6030), .A2 (n_6027), .A3 (n_6029));
NAND2_X1 i_6062 (.ZN (n_5998), .A1 (n_6030), .A2 (n_6029));
NAND3_X1 i_6061 (.ZN (n_5997), .A1 (n_5998), .A2 (n_6117), .A3 (n_6028));
NAND2_X1 i_6060 (.ZN (n_5996), .A1 (n_5997), .A2 (n_5999));
AOI21_X1 i_6059 (.ZN (n_5995), .A (n_5996), .B1 (n_6000), .B2 (n_6002));
NAND3_X1 i_6058 (.ZN (n_5994), .A1 (n_6000), .A2 (n_6002), .A3 (n_5996));
NAND3_X1 i_6057 (.ZN (n_5993), .A1 (n_6612), .A2 (n_6623), .A3 (n_6616));
INV_X1 i_6056 (.ZN (n_5992), .A (n_5993));
AOI21_X1 i_6055 (.ZN (n_5991), .A (n_6616), .B1 (n_6623), .B2 (n_6612));
NOR2_X1 i_6054 (.ZN (n_5990), .A1 (n_5992), .A2 (n_5991));
NAND3_X1 i_6053 (.ZN (n_5989), .A1 (n_6633), .A2 (n_6631), .A3 (n_6626));
INV_X1 i_6052 (.ZN (n_5988), .A (n_5989));
AOI21_X1 i_6051 (.ZN (n_5987), .A (n_6626), .B1 (n_6633), .B2 (n_6631));
NOR2_X1 i_6050 (.ZN (n_5986), .A1 (n_5988), .A2 (n_5987));
NAND2_X1 i_6049 (.ZN (n_5985), .A1 (A_imm[24]), .A2 (B_imm[4]));
OAI21_X1 i_6048 (.ZN (n_5984), .A (n_5985), .B1 (n_8907), .B2 (n_8429));
NAND2_X1 i_6047 (.ZN (n_5983), .A1 (B_imm[12]), .A2 (A_imm[16]));
NAND4_X1 i_6046 (.ZN (n_5982), .A1 (A_imm[23]), .A2 (A_imm[24]), .A3 (B_imm[5]), .A4 (B_imm[4]));
NAND2_X1 i_6045 (.ZN (n_5981), .A1 (n_5982), .A2 (n_5983));
AOI22_X1 i_6044 (.ZN (n_5980), .A1 (n_5981), .A2 (n_5984), .B1 (B_imm[29]), .B2 (A_imm[0]));
INV_X1 i_6043 (.ZN (n_5979), .A (n_5980));
NAND2_X1 i_6042 (.ZN (n_5978), .A1 (A_imm[28]), .A2 (B_imm[1]));
NAND4_X1 i_6041 (.ZN (n_5977), .A1 (n_5981), .A2 (B_imm[29]), .A3 (A_imm[0]), .A4 (n_5984));
NAND2_X1 i_6040 (.ZN (n_5976), .A1 (n_5977), .A2 (n_5978));
AOI21_X1 i_6039 (.ZN (n_5975), .A (n_6219), .B1 (n_6220), .B2 (n_6217));
NAND3_X1 i_6038 (.ZN (n_5974), .A1 (n_6220), .A2 (n_6219), .A3 (n_6217));
INV_X1 i_6037 (.ZN (n_5973), .A (n_5974));
NOR2_X1 i_6036 (.ZN (n_5972), .A1 (n_5973), .A2 (n_5975));
INV_X1 i_6035 (.ZN (n_5971), .A (n_5972));
NAND3_X1 i_6034 (.ZN (n_5970), .A1 (n_5971), .A2 (n_5976), .A3 (n_5979));
AOI21_X1 i_6033 (.ZN (n_5969), .A (n_6288), .B1 (n_6295), .B2 (n_6287));
NAND3_X1 i_6032 (.ZN (n_5968), .A1 (n_6295), .A2 (n_6288), .A3 (n_6287));
INV_X1 i_6031 (.ZN (n_5967), .A (n_5968));
NOR2_X1 i_6030 (.ZN (n_5966), .A1 (n_5967), .A2 (n_5969));
INV_X1 i_6029 (.ZN (n_5965), .A (n_5966));
NAND2_X1 i_6028 (.ZN (n_5964), .A1 (n_5976), .A2 (n_5979));
NAND2_X1 i_6027 (.ZN (n_5963), .A1 (n_5964), .A2 (n_5972));
NAND2_X1 i_6026 (.ZN (n_5962), .A1 (n_5963), .A2 (n_5965));
AOI22_X1 i_6025 (.ZN (n_5961), .A1 (n_6312), .A2 (n_6315), .B1 (B_imm[30]), .B2 (A_imm[1]));
OAI21_X1 i_6024 (.ZN (n_5960), .A (n_6282), .B1 (n_6281), .B2 (n_5961));
NAND3_X1 i_6023 (.ZN (n_5959), .A1 (n_6310), .A2 (n_6308), .A3 (n_6309));
NAND4_X1 i_6022 (.ZN (n_5958), .A1 (n_5962), .A2 (n_5970), .A3 (n_5960), .A4 (n_5959));
INV_X1 i_6021 (.ZN (n_5957), .A (n_5970));
AOI21_X1 i_6020 (.ZN (n_5956), .A (n_5966), .B1 (n_5964), .B2 (n_5972));
NAND2_X1 i_6019 (.ZN (n_5955), .A1 (n_5960), .A2 (n_5959));
OAI21_X1 i_6018 (.ZN (n_5954), .A (n_5955), .B1 (n_5957), .B2 (n_5956));
AOI21_X1 i_6017 (.ZN (n_5953), .A (n_6314), .B1 (n_6315), .B2 (n_6313));
INV_X1 i_6016 (.ZN (n_5952), .A (n_5953));
NAND3_X1 i_6015 (.ZN (n_5951), .A1 (n_6315), .A2 (n_6313), .A3 (n_6314));
NAND2_X1 i_6014 (.ZN (n_5950), .A1 (n_5952), .A2 (n_5951));
INV_X1 i_6013 (.ZN (n_5949), .A (n_5950));
OAI21_X1 i_6012 (.ZN (n_5948), .A (n_5949), .B1 (n_9005), .B2 (n_6740));
NAND2_X1 i_6011 (.ZN (n_5947), .A1 (A_imm[27]), .A2 (B_imm[2]));
NAND2_X1 i_6010 (.ZN (n_5946), .A1 (B_imm[13]), .A2 (A_imm[15]));
OAI21_X1 i_6009 (.ZN (n_5945), .A (n_5946), .B1 (n_8860), .B2 (n_8511));
NAND2_X1 i_6008 (.ZN (n_5944), .A1 (B_imm[28]), .A2 (A_imm[0]));
INV_X1 i_6007 (.ZN (n_5943), .A (n_5944));
NAND4_X1 i_6006 (.ZN (n_5942), .A1 (B_imm[20]), .A2 (B_imm[13]), .A3 (A_imm[15]), .A4 (A_imm[8]));
INV_X1 i_6005 (.ZN (n_5941), .A (n_5942));
OAI21_X2 i_6004 (.ZN (n_5940), .A (n_5945), .B1 (n_5941), .B2 (n_5943));
NAND2_X1 i_6003 (.ZN (n_5939), .A1 (n_5940), .A2 (n_5947));
OAI22_X1 i_6002 (.ZN (n_5938), .A1 (n_8880), .A2 (n_8955), .B1 (n_8751), .B2 (n_8909));
NAND2_X1 i_6001 (.ZN (n_5937), .A1 (B_imm[16]), .A2 (A_imm[11]));
NAND4_X1 i_6000 (.ZN (n_5936), .A1 (A_imm[17]), .A2 (A_imm[10]), .A3 (B_imm[17]), .A4 (B_imm[10]));
NAND2_X1 i_5999 (.ZN (n_5935), .A1 (n_5936), .A2 (n_5937));
NAND2_X1 i_5998 (.ZN (n_5934), .A1 (n_5935), .A2 (n_5938));
OAI21_X1 i_5997 (.ZN (n_5933), .A (n_5934), .B1 (n_8821), .B2 (n_8293));
NAND2_X1 i_5996 (.ZN (n_5932), .A1 (B_imm[21]), .A2 (A_imm[7]));
INV_X1 i_5995 (.ZN (n_5931), .A (n_5932));
NAND4_X1 i_5994 (.ZN (n_5930), .A1 (n_5935), .A2 (n_5938), .A3 (B_imm[23]), .A4 (A_imm[5]));
INV_X1 i_5993 (.ZN (n_5929), .A (n_5930));
OAI21_X1 i_5992 (.ZN (n_5928), .A (n_5933), .B1 (n_5929), .B2 (n_5931));
OAI21_X1 i_5991 (.ZN (n_5927), .A (n_5928), .B1 (n_5940), .B2 (n_5947));
NAND2_X1 i_5990 (.ZN (n_5926), .A1 (n_5927), .A2 (n_5939));
NAND3_X1 i_5989 (.ZN (n_5925), .A1 (n_5950), .A2 (B_imm[0]), .A3 (A_imm[30]));
NAND2_X1 i_5988 (.ZN (n_5924), .A1 (n_5925), .A2 (n_5926));
NAND2_X1 i_5987 (.ZN (n_5923), .A1 (n_5924), .A2 (n_5948));
NAND2_X1 i_5986 (.ZN (n_5922), .A1 (n_5954), .A2 (n_5923));
NAND2_X1 i_5985 (.ZN (n_5921), .A1 (n_6258), .A2 (n_6256));
NAND3_X1 i_5984 (.ZN (n_5920), .A1 (n_5921), .A2 (B_imm[2]), .A3 (A_imm[30]));
NAND3_X1 i_5983 (.ZN (n_5919), .A1 (n_6258), .A2 (n_6257), .A3 (n_6256));
NAND2_X1 i_5982 (.ZN (n_5918), .A1 (n_5920), .A2 (n_5919));
NAND3_X1 i_5981 (.ZN (n_5917), .A1 (n_5922), .A2 (n_5918), .A3 (n_5958));
INV_X1 i_5980 (.ZN (n_5916), .A (n_5917));
AOI21_X1 i_5979 (.ZN (n_5915), .A (n_5918), .B1 (n_5922), .B2 (n_5958));
INV_X1 i_5978 (.ZN (n_5914), .A (n_5915));
INV_X1 i_5977 (.ZN (n_5913), .A (n_6665));
OAI21_X1 i_5976 (.ZN (n_5912), .A (n_6664), .B1 (n_5913), .B2 (n_6663));
INV_X1 i_5975 (.ZN (n_5911), .A (n_6663));
NAND4_X1 i_5974 (.ZN (n_5910), .A1 (n_5911), .A2 (B_imm[14]), .A3 (A_imm[17]), .A4 (n_6665));
NAND2_X1 i_5973 (.ZN (n_5909), .A1 (n_5910), .A2 (n_5912));
INV_X1 i_5972 (.ZN (n_5908), .A (n_5909));
NAND2_X1 i_5971 (.ZN (n_5907), .A1 (B_imm[18]), .A2 (A_imm[10]));
OAI21_X1 i_5970 (.ZN (n_5906), .A (n_5907), .B1 (n_8347), .B2 (n_8892));
NAND2_X1 i_5969 (.ZN (n_5905), .A1 (B_imm[24]), .A2 (A_imm[4]));
NAND4_X1 i_5968 (.ZN (n_5904), .A1 (B_imm[9]), .A2 (B_imm[18]), .A3 (A_imm[19]), .A4 (A_imm[10]));
NAND2_X1 i_5967 (.ZN (n_5903), .A1 (n_5904), .A2 (n_5905));
NAND2_X1 i_5966 (.ZN (n_5902), .A1 (n_5903), .A2 (n_5906));
NAND2_X1 i_5965 (.ZN (n_5901), .A1 (B_imm[11]), .A2 (A_imm[17]));
OAI21_X1 i_5964 (.ZN (n_5900), .A (n_5901), .B1 (n_8794), .B2 (n_6817));
NAND2_X1 i_5963 (.ZN (n_5899), .A1 (A_imm[26]), .A2 (B_imm[2]));
NAND4_X1 i_5962 (.ZN (n_5898), .A1 (A_imm[25]), .A2 (B_imm[11]), .A3 (B_imm[3]), .A4 (A_imm[17]));
NAND2_X1 i_5961 (.ZN (n_5897), .A1 (n_5898), .A2 (n_5899));
NAND2_X1 i_5960 (.ZN (n_5896), .A1 (n_5897), .A2 (n_5900));
NAND2_X1 i_5959 (.ZN (n_5895), .A1 (n_5902), .A2 (n_5896));
NAND2_X1 i_5958 (.ZN (n_5894), .A1 (B_imm[22]), .A2 (A_imm[6]));
OAI21_X1 i_5957 (.ZN (n_5893), .A (n_5894), .B1 (n_8829), .B2 (n_8927));
NAND2_X1 i_5956 (.ZN (n_5892), .A1 (B_imm[25]), .A2 (A_imm[3]));
INV_X1 i_5955 (.ZN (n_5891), .A (n_5892));
NAND4_X1 i_5954 (.ZN (n_5890), .A1 (B_imm[15]), .A2 (B_imm[22]), .A3 (A_imm[13]), .A4 (A_imm[6]));
INV_X1 i_5953 (.ZN (n_5889), .A (n_5890));
OAI21_X1 i_5952 (.ZN (n_5888), .A (n_5893), .B1 (n_5889), .B2 (n_5891));
NAND4_X1 i_5951 (.ZN (n_5887), .A1 (n_5903), .A2 (n_5897), .A3 (n_5906), .A4 (n_5900));
NAND2_X1 i_5950 (.ZN (n_5886), .A1 (n_5887), .A2 (n_5888));
NAND2_X1 i_5949 (.ZN (n_5885), .A1 (n_6303), .A2 (n_6300));
NAND2_X1 i_5948 (.ZN (n_5884), .A1 (n_5885), .A2 (n_6301));
NAND3_X1 i_5947 (.ZN (n_5883), .A1 (n_6303), .A2 (n_6300), .A3 (n_6302));
NAND2_X1 i_5946 (.ZN (n_5882), .A1 (n_5884), .A2 (n_5883));
NAND3_X2 i_5945 (.ZN (n_5881), .A1 (n_5886), .A2 (n_5882), .A3 (n_5895));
NAND2_X1 i_5944 (.ZN (n_5880), .A1 (n_5886), .A2 (n_5895));
INV_X1 i_5943 (.ZN (n_5879), .A (n_5882));
NAND2_X1 i_5942 (.ZN (n_5878), .A1 (n_5880), .A2 (n_5879));
NAND2_X1 i_5941 (.ZN (n_5877), .A1 (n_6676), .A2 (n_6674));
NAND3_X1 i_5940 (.ZN (n_5876), .A1 (n_5877), .A2 (B_imm[19]), .A3 (A_imm[11]));
NAND3_X1 i_5939 (.ZN (n_5875), .A1 (n_6676), .A2 (n_6675), .A3 (n_6674));
NAND2_X1 i_5938 (.ZN (n_5874), .A1 (n_5876), .A2 (n_5875));
NAND2_X1 i_5937 (.ZN (n_5873), .A1 (n_5878), .A2 (n_5874));
NAND2_X1 i_5936 (.ZN (n_5872), .A1 (n_5873), .A2 (n_5881));
NAND2_X1 i_5935 (.ZN (n_5871), .A1 (n_5872), .A2 (n_5908));
NAND3_X1 i_5934 (.ZN (n_5870), .A1 (n_5909), .A2 (n_5873), .A3 (n_5881));
INV_X1 i_5933 (.ZN (n_5869), .A (n_6646));
OAI21_X1 i_5932 (.ZN (n_5868), .A (n_6637), .B1 (n_6643), .B2 (n_5869));
OAI211_X1 i_5931 (.ZN (n_5867), .A (n_6644), .B (n_6646), .C1 (n_6640), .C2 (n_6638));
NAND2_X1 i_5930 (.ZN (n_5866), .A1 (n_5868), .A2 (n_5867));
INV_X1 i_5929 (.ZN (n_5865), .A (n_5866));
NAND2_X1 i_5928 (.ZN (n_5864), .A1 (n_5870), .A2 (n_5865));
NAND2_X1 i_5927 (.ZN (n_5863), .A1 (n_5864), .A2 (n_5871));
NAND2_X1 i_5926 (.ZN (n_5862), .A1 (n_5914), .A2 (n_5863));
INV_X1 i_5925 (.ZN (n_5861), .A (n_5862));
OAI21_X2 i_5924 (.ZN (n_5860), .A (n_5986), .B1 (n_5916), .B2 (n_5861));
OAI211_X1 i_5923 (.ZN (n_5859), .A (n_5917), .B (n_5862), .C1 (n_5988), .C2 (n_5987));
INV_X1 i_5922 (.ZN (n_5858), .A (n_6636));
NAND2_X1 i_5921 (.ZN (n_5857), .A1 (n_6658), .A2 (n_6661));
NAND2_X1 i_5920 (.ZN (n_5856), .A1 (n_5857), .A2 (n_5858));
NAND3_X1 i_5919 (.ZN (n_5855), .A1 (n_6636), .A2 (n_6658), .A3 (n_6661));
NAND2_X1 i_5918 (.ZN (n_5854), .A1 (n_5856), .A2 (n_5855));
INV_X1 i_5917 (.ZN (n_5853), .A (n_5854));
INV_X1 i_5916 (.ZN (n_5852), .A (n_6563));
OAI21_X1 i_5915 (.ZN (n_5851), .A (n_6560), .B1 (n_5852), .B2 (n_6562));
NAND2_X1 i_5914 (.ZN (n_5850), .A1 (n_6569), .A2 (n_6578));
NAND3_X1 i_5913 (.ZN (n_5849), .A1 (n_5850), .A2 (n_6566), .A3 (n_6565));
INV_X1 i_5912 (.ZN (n_5848), .A (n_6560));
NAND3_X1 i_5911 (.ZN (n_5847), .A1 (n_5849), .A2 (n_6563), .A3 (n_5848));
INV_X1 i_5910 (.ZN (n_5846), .A (n_6649));
INV_X1 i_5909 (.ZN (n_5845), .A (n_6648));
OAI21_X1 i_5908 (.ZN (n_5844), .A (n_5846), .B1 (n_5845), .B2 (n_6651));
NAND3_X1 i_5907 (.ZN (n_5843), .A1 (n_6650), .A2 (n_6649), .A3 (n_6648));
NAND2_X1 i_5906 (.ZN (n_5842), .A1 (B_imm[14]), .A2 (A_imm[15]));
INV_X1 i_5905 (.ZN (n_5841), .A (n_6293));
OAI21_X1 i_5904 (.ZN (n_5840), .A (n_6291), .B1 (n_5841), .B2 (n_6289));
NAND3_X1 i_5903 (.ZN (n_5839), .A1 (n_6293), .A2 (n_6292), .A3 (n_6290));
NAND3_X1 i_5902 (.ZN (n_5838), .A1 (n_5842), .A2 (n_5840), .A3 (n_5839));
NAND2_X1 i_5901 (.ZN (n_5837), .A1 (n_5840), .A2 (n_5839));
NAND3_X1 i_5900 (.ZN (n_5836), .A1 (n_5837), .A2 (B_imm[14]), .A3 (A_imm[15]));
AOI21_X1 i_5899 (.ZN (n_5835), .A (n_6654), .B1 (n_6655), .B2 (n_6653));
NAND3_X1 i_5898 (.ZN (n_5834), .A1 (n_6655), .A2 (n_6654), .A3 (n_6653));
INV_X1 i_5897 (.ZN (n_5833), .A (n_5834));
NOR2_X1 i_5896 (.ZN (n_5832), .A1 (n_5835), .A2 (n_5833));
NAND2_X1 i_5895 (.ZN (n_5831), .A1 (n_5836), .A2 (n_5832));
NAND2_X1 i_5894 (.ZN (n_5830), .A1 (n_5831), .A2 (n_5838));
NAND3_X1 i_5893 (.ZN (n_5829), .A1 (n_5830), .A2 (n_5844), .A3 (n_5843));
AOI21_X1 i_5892 (.ZN (n_5828), .A (n_6571), .B1 (n_6570), .B2 (n_6578));
NAND3_X1 i_5891 (.ZN (n_5827), .A1 (n_6578), .A2 (n_6570), .A3 (n_6571));
INV_X1 i_5890 (.ZN (n_5826), .A (n_5827));
NOR2_X1 i_5889 (.ZN (n_5825), .A1 (n_5826), .A2 (n_5828));
NAND2_X1 i_5888 (.ZN (n_5824), .A1 (n_5843), .A2 (n_5844));
NAND3_X1 i_5887 (.ZN (n_5823), .A1 (n_5824), .A2 (n_5838), .A3 (n_5831));
NAND2_X1 i_5886 (.ZN (n_5822), .A1 (n_5825), .A2 (n_5823));
NAND4_X2 i_5885 (.ZN (n_5821), .A1 (n_5822), .A2 (n_5851), .A3 (n_5847), .A4 (n_5829));
NAND2_X1 i_5884 (.ZN (n_5820), .A1 (n_5851), .A2 (n_5847));
NAND2_X1 i_5883 (.ZN (n_5819), .A1 (n_5822), .A2 (n_5829));
NAND2_X1 i_5882 (.ZN (n_5818), .A1 (n_5820), .A2 (n_5819));
INV_X1 i_5881 (.ZN (n_5817), .A (n_6470));
NAND2_X1 i_5880 (.ZN (n_5816), .A1 (n_6477), .A2 (n_6468));
NAND2_X1 i_5879 (.ZN (n_5815), .A1 (n_5816), .A2 (n_5817));
NAND3_X1 i_5878 (.ZN (n_5814), .A1 (n_6477), .A2 (n_6468), .A3 (n_6470));
NAND2_X1 i_5877 (.ZN (n_5813), .A1 (n_5815), .A2 (n_5814));
OAI22_X1 i_5876 (.ZN (n_5812), .A1 (n_8232), .A2 (n_8859), .B1 (n_8906), .B2 (n_8429));
NAND2_X1 i_5875 (.ZN (n_5811), .A1 (A_imm[20]), .A2 (B_imm[7]));
NAND4_X1 i_5874 (.ZN (n_5810), .A1 (B_imm[6]), .A2 (A_imm[21]), .A3 (A_imm[22]), .A4 (B_imm[5]));
NAND2_X1 i_5873 (.ZN (n_5809), .A1 (n_5810), .A2 (n_5811));
NAND2_X1 i_5872 (.ZN (n_5808), .A1 (n_5809), .A2 (n_5812));
OAI21_X1 i_5871 (.ZN (n_5807), .A (n_5808), .B1 (n_8993), .B2 (n_6677));
NAND2_X1 i_5870 (.ZN (n_5806), .A1 (B_imm[19]), .A2 (A_imm[9]));
NAND4_X2 i_5869 (.ZN (n_5805), .A1 (n_5809), .A2 (B_imm[26]), .A3 (A_imm[2]), .A4 (n_5812));
NAND2_X1 i_5868 (.ZN (n_5804), .A1 (n_5805), .A2 (n_5806));
NAND4_X1 i_5867 (.ZN (n_5803), .A1 (n_5804), .A2 (B_imm[0]), .A3 (A_imm[29]), .A4 (n_5807));
NAND2_X1 i_5866 (.ZN (n_5802), .A1 (A_imm[29]), .A2 (B_imm[0]));
INV_X1 i_5865 (.ZN (n_5801), .A (n_5806));
INV_X1 i_5864 (.ZN (n_5800), .A (n_5805));
OAI21_X1 i_5863 (.ZN (n_5799), .A (n_5807), .B1 (n_5800), .B2 (n_5801));
NAND2_X1 i_5862 (.ZN (n_5798), .A1 (n_5799), .A2 (n_5802));
NAND2_X1 i_5861 (.ZN (n_5797), .A1 (n_6576), .A2 (n_6573));
NAND2_X1 i_5860 (.ZN (n_5796), .A1 (n_5797), .A2 (n_6574));
NAND3_X1 i_5859 (.ZN (n_5795), .A1 (n_6576), .A2 (n_6575), .A3 (n_6573));
NAND2_X1 i_5858 (.ZN (n_5794), .A1 (n_5796), .A2 (n_5795));
NAND2_X1 i_5857 (.ZN (n_5793), .A1 (n_5798), .A2 (n_5794));
NAND2_X1 i_5856 (.ZN (n_5792), .A1 (n_5793), .A2 (n_5803));
NAND2_X1 i_5855 (.ZN (n_5791), .A1 (n_5792), .A2 (n_5813));
NAND4_X1 i_5854 (.ZN (n_5790), .A1 (n_5793), .A2 (n_5815), .A3 (n_5814), .A4 (n_5803));
OAI22_X1 i_5853 (.ZN (n_5789), .A1 (n_6577), .A2 (n_8907), .B1 (n_8947), .B2 (n_8892));
NAND2_X1 i_5852 (.ZN (n_5788), .A1 (A_imm[24]), .A2 (B_imm[3]));
NAND4_X1 i_5851 (.ZN (n_5787), .A1 (A_imm[23]), .A2 (B_imm[8]), .A3 (B_imm[4]), .A4 (A_imm[19]));
NAND2_X1 i_5850 (.ZN (n_5786), .A1 (n_5787), .A2 (n_5788));
NAND2_X1 i_5849 (.ZN (n_5785), .A1 (n_5786), .A2 (n_5789));
OAI21_X1 i_5848 (.ZN (n_5784), .A (n_5785), .B1 (n_9003), .B2 (n_6836));
OAI22_X1 i_5847 (.ZN (n_5783), .A1 (n_8849), .A2 (n_8858), .B1 (n_8795), .B2 (n_8946));
NAND2_X1 i_5846 (.ZN (n_5782), .A1 (A_imm[25]), .A2 (B_imm[2]));
INV_X1 i_5845 (.ZN (n_5781), .A (n_5782));
NAND4_X1 i_5844 (.ZN (n_5780), .A1 (B_imm[11]), .A2 (B_imm[12]), .A3 (A_imm[16]), .A4 (A_imm[15]));
INV_X1 i_5843 (.ZN (n_5779), .A (n_5780));
OAI21_X1 i_5842 (.ZN (n_5778), .A (n_5783), .B1 (n_5779), .B2 (n_5781));
NAND4_X1 i_5841 (.ZN (n_5777), .A1 (n_5786), .A2 (n_5789), .A3 (B_imm[27]), .A4 (A_imm[1]));
NAND2_X1 i_5840 (.ZN (n_5776), .A1 (n_5777), .A2 (n_5778));
AOI21_X1 i_5839 (.ZN (n_5775), .A (n_6582), .B1 (n_6583), .B2 (n_6581));
INV_X1 i_5838 (.ZN (n_5774), .A (n_5775));
NAND3_X1 i_5837 (.ZN (n_5773), .A1 (n_6583), .A2 (n_6582), .A3 (n_6581));
NAND2_X1 i_5836 (.ZN (n_5772), .A1 (n_5774), .A2 (n_5773));
NAND3_X1 i_5835 (.ZN (n_5771), .A1 (n_5776), .A2 (n_5784), .A3 (n_5772));
NAND2_X1 i_5834 (.ZN (n_5770), .A1 (n_5776), .A2 (n_5784));
INV_X1 i_5833 (.ZN (n_5769), .A (n_5772));
NAND2_X1 i_5832 (.ZN (n_5768), .A1 (n_5770), .A2 (n_5769));
INV_X1 i_5831 (.ZN (n_5767), .A (n_6483));
OAI21_X1 i_5830 (.ZN (n_5766), .A (n_6481), .B1 (n_5767), .B2 (n_6479));
NAND3_X1 i_5829 (.ZN (n_5765), .A1 (n_6483), .A2 (n_6482), .A3 (n_6480));
NAND2_X1 i_5828 (.ZN (n_5764), .A1 (n_5766), .A2 (n_5765));
NAND2_X1 i_5827 (.ZN (n_5763), .A1 (n_5768), .A2 (n_5764));
NAND2_X1 i_5826 (.ZN (n_5762), .A1 (n_5763), .A2 (n_5771));
NAND2_X1 i_5825 (.ZN (n_5761), .A1 (n_5762), .A2 (n_5790));
NAND2_X1 i_5824 (.ZN (n_5760), .A1 (n_5761), .A2 (n_5791));
NAND2_X1 i_5823 (.ZN (n_5759), .A1 (n_5818), .A2 (n_5760));
NAND2_X1 i_5822 (.ZN (n_5758), .A1 (n_5759), .A2 (n_5821));
NAND2_X1 i_5821 (.ZN (n_5757), .A1 (n_5758), .A2 (n_5853));
NAND3_X1 i_5820 (.ZN (n_5756), .A1 (n_5759), .A2 (n_5854), .A3 (n_5821));
INV_X1 i_5819 (.ZN (n_5755), .A (n_5756));
NAND2_X1 i_5818 (.ZN (n_5754), .A1 (n_6586), .A2 (n_6585));
XNOR2_X1 i_5817 (.ZN (n_5753), .A (n_5754), .B (n_6559));
INV_X1 i_5816 (.ZN (n_5752), .A (n_5753));
OAI21_X1 i_5815 (.ZN (n_5751), .A (n_5757), .B1 (n_5752), .B2 (n_5755));
NAND2_X1 i_5814 (.ZN (n_5750), .A1 (n_5859), .A2 (n_5751));
NAND2_X1 i_5813 (.ZN (n_5749), .A1 (n_5750), .A2 (n_5860));
NAND2_X1 i_5812 (.ZN (n_5748), .A1 (n_5749), .A2 (n_5990));
OAI211_X2 i_5811 (.ZN (n_5747), .A (n_5750), .B (n_5860), .C1 (n_5992), .C2 (n_5991));
INV_X2 i_5810 (.ZN (n_5746), .A (n_5747));
INV_X1 i_5809 (.ZN (n_5745), .A (n_6385));
NAND2_X1 i_5808 (.ZN (n_5744), .A1 (n_6395), .A2 (n_6390));
NAND2_X1 i_5807 (.ZN (n_5743), .A1 (n_5744), .A2 (n_5745));
NAND3_X1 i_5806 (.ZN (n_5742), .A1 (n_6395), .A2 (n_6390), .A3 (n_6385));
NAND2_X1 i_5805 (.ZN (n_5741), .A1 (n_5743), .A2 (n_5742));
OAI21_X2 i_5804 (.ZN (n_5740), .A (n_5748), .B1 (n_5746), .B2 (n_5741));
NAND2_X1 i_5803 (.ZN (n_5739), .A1 (n_5740), .A2 (n_5994));
INV_X1 i_5802 (.ZN (n_5738), .A (n_5739));
OAI21_X2 i_5801 (.ZN (n_5737), .A (n_6003), .B1 (n_5738), .B2 (n_5995));
INV_X1 i_5800 (.ZN (n_5736), .A (n_6003));
NAND2_X1 i_5799 (.ZN (n_5735), .A1 (n_6000), .A2 (n_6002));
INV_X1 i_5798 (.ZN (n_5734), .A (n_5996));
NAND2_X1 i_5797 (.ZN (n_5733), .A1 (n_5735), .A2 (n_5734));
NAND3_X1 i_5796 (.ZN (n_5732), .A1 (n_5739), .A2 (n_5736), .A3 (n_5733));
INV_X1 i_5795 (.ZN (n_5731), .A (n_5732));
NAND3_X1 i_5794 (.ZN (n_5730), .A1 (n_6092), .A2 (n_6602), .A3 (n_6601));
NAND2_X1 i_5793 (.ZN (n_5729), .A1 (n_6602), .A2 (n_6601));
NAND3_X1 i_5792 (.ZN (n_5728), .A1 (n_5729), .A2 (n_6382), .A3 (n_6093));
NAND2_X1 i_5791 (.ZN (n_5727), .A1 (n_5728), .A2 (n_5730));
OAI21_X1 i_5790 (.ZN (n_5726), .A (n_5737), .B1 (n_5727), .B2 (n_5731));
INV_X1 i_5789 (.ZN (n_5725), .A (n_5726));
NAND3_X1 i_5788 (.ZN (n_5724), .A1 (n_5725), .A2 (n_6008), .A3 (n_6010));
NAND2_X1 i_5787 (.ZN (n_5723), .A1 (n_6770), .A2 (n_6852));
NAND2_X1 i_5786 (.ZN (n_5722), .A1 (n_5723), .A2 (n_6849));
NAND3_X1 i_5785 (.ZN (n_5721), .A1 (n_7583), .A2 (n_7582), .A3 (n_7576));
AOI21_X1 i_5784 (.ZN (n_5720), .A (n_7717), .B1 (n_7585), .B2 (n_7643));
INV_X1 i_5783 (.ZN (n_5719), .A (n_7576));
OAI21_X2 i_5782 (.ZN (n_5718), .A (n_5719), .B1 (n_7581), .B2 (n_5720));
NAND2_X1 i_5781 (.ZN (n_5717), .A1 (n_5718), .A2 (n_5721));
NAND2_X1 i_5780 (.ZN (n_5716), .A1 (n_6060), .A2 (n_6050));
NAND2_X1 i_5779 (.ZN (n_5715), .A1 (n_5716), .A2 (n_6058));
NAND2_X1 i_5778 (.ZN (n_5714), .A1 (n_5717), .A2 (n_5715));
NAND4_X1 i_5777 (.ZN (n_5713), .A1 (n_5718), .A2 (n_5721), .A3 (n_6058), .A4 (n_5716));
NAND3_X1 i_5776 (.ZN (n_5712), .A1 (n_5714), .A2 (n_5722), .A3 (n_5713));
INV_X1 i_5775 (.ZN (n_5711), .A (n_6849));
AOI21_X1 i_5774 (.ZN (n_5710), .A (n_5711), .B1 (n_6852), .B2 (n_6770));
NAND2_X1 i_5773 (.ZN (n_5709), .A1 (n_5714), .A2 (n_5713));
NAND2_X1 i_5772 (.ZN (n_5708), .A1 (n_5709), .A2 (n_5710));
NAND2_X1 i_5771 (.ZN (n_5707), .A1 (n_5708), .A2 (n_5712));
NAND2_X1 i_5770 (.ZN (n_5706), .A1 (n_7481), .A2 (n_7483));
NAND3_X1 i_5769 (.ZN (n_5705), .A1 (n_7485), .A2 (n_5706), .A3 (n_7484));
INV_X1 i_5768 (.ZN (n_5704), .A (n_5706));
NAND2_X1 i_5767 (.ZN (n_5703), .A1 (n_7485), .A2 (n_7484));
NAND2_X1 i_5766 (.ZN (n_5702), .A1 (n_5703), .A2 (n_5704));
NAND2_X1 i_5765 (.ZN (n_5701), .A1 (n_5702), .A2 (n_5705));
NAND2_X2 i_5764 (.ZN (n_5700), .A1 (n_6016), .A2 (n_6044));
NAND2_X1 i_5763 (.ZN (n_5699), .A1 (n_5700), .A2 (n_6042));
NAND2_X1 i_5762 (.ZN (n_5698), .A1 (n_5699), .A2 (n_5701));
INV_X1 i_5761 (.ZN (n_5697), .A (n_5701));
NAND3_X1 i_5760 (.ZN (n_5696), .A1 (n_5700), .A2 (n_5697), .A3 (n_6042));
NAND3_X1 i_5759 (.ZN (n_5695), .A1 (n_5707), .A2 (n_5698), .A3 (n_5696));
INV_X1 i_5758 (.ZN (n_5694), .A (n_5707));
NAND2_X1 i_5757 (.ZN (n_5693), .A1 (n_5698), .A2 (n_5696));
NAND2_X1 i_5756 (.ZN (n_5692), .A1 (n_5693), .A2 (n_5694));
INV_X1 i_5755 (.ZN (n_5691), .A (n_6011));
NAND2_X2 i_5754 (.ZN (n_5690), .A1 (n_6088), .A2 (n_5691));
NAND4_X4 i_5753 (.ZN (n_5689), .A1 (n_5692), .A2 (n_6089), .A3 (n_5695), .A4 (n_5690));
NAND3_X1 i_5752 (.ZN (n_5688), .A1 (n_7469), .A2 (n_7476), .A3 (n_7475));
INV_X1 i_5751 (.ZN (n_5687), .A (n_5688));
AOI22_X1 i_5750 (.ZN (n_5686), .A1 (n_7476), .A2 (n_7475), .B1 (n_7472), .B2 (n_7471));
NAND3_X1 i_5749 (.ZN (n_5685), .A1 (n_7920), .A2 (n_8068), .A3 (n_8066));
INV_X1 i_5748 (.ZN (n_5684), .A (n_7920));
NAND2_X1 i_5747 (.ZN (n_5683), .A1 (n_8068), .A2 (n_8066));
NAND2_X1 i_5746 (.ZN (n_5682), .A1 (n_5683), .A2 (n_5684));
NAND2_X1 i_5745 (.ZN (n_5681), .A1 (n_5682), .A2 (n_5685));
INV_X1 i_5744 (.ZN (n_5680), .A (n_5713));
OAI21_X1 i_5743 (.ZN (n_5679), .A (n_5714), .B1 (n_5680), .B2 (n_5710));
NAND2_X1 i_5742 (.ZN (n_5678), .A1 (n_5679), .A2 (n_5681));
INV_X1 i_5741 (.ZN (n_5677), .A (n_5681));
NAND2_X1 i_5740 (.ZN (n_5676), .A1 (n_5722), .A2 (n_5713));
NAND3_X2 i_5739 (.ZN (n_5675), .A1 (n_5677), .A2 (n_5676), .A3 (n_5714));
INV_X1 i_5738 (.ZN (n_5674), .A (n_5675));
NAND3_X1 i_5737 (.ZN (n_5673), .A1 (n_7571), .A2 (n_7479), .A3 (n_7574));
INV_X1 i_5736 (.ZN (n_5672), .A (n_7479));
NAND2_X1 i_5735 (.ZN (n_5671), .A1 (n_7571), .A2 (n_7574));
NAND2_X1 i_5734 (.ZN (n_5670), .A1 (n_5671), .A2 (n_5672));
NAND2_X1 i_5733 (.ZN (n_5669), .A1 (n_5670), .A2 (n_5673));
OAI21_X1 i_5732 (.ZN (n_5668), .A (n_5678), .B1 (n_5674), .B2 (n_5669));
INV_X1 i_5731 (.ZN (n_5667), .A (n_5668));
OAI21_X2 i_5730 (.ZN (n_5666), .A (n_5667), .B1 (n_5687), .B2 (n_5686));
NAND3_X1 i_5729 (.ZN (n_5665), .A1 (n_5678), .A2 (n_5675), .A3 (n_5669));
INV_X1 i_5728 (.ZN (n_5664), .A (n_5669));
NAND2_X1 i_5727 (.ZN (n_5663), .A1 (n_5678), .A2 (n_5675));
NAND2_X1 i_5726 (.ZN (n_5662), .A1 (n_5663), .A2 (n_5664));
NAND3_X1 i_5725 (.ZN (n_5661), .A1 (n_5696), .A2 (n_5712), .A3 (n_5708));
NAND2_X1 i_5724 (.ZN (n_5660), .A1 (n_5661), .A2 (n_5698));
INV_X1 i_5723 (.ZN (n_5659), .A (n_5660));
NAND3_X2 i_5722 (.ZN (n_5658), .A1 (n_5659), .A2 (n_5662), .A3 (n_5665));
NAND3_X2 i_5721 (.ZN (n_5657), .A1 (n_5689), .A2 (n_5666), .A3 (n_5658));
NAND2_X1 i_5719 (.ZN (n_5655), .A1 (n_6998), .A2 (n_7199));
NAND2_X1 i_5718 (.ZN (n_5654), .A1 (A_imm[29]), .A2 (B_imm[16]));
INV_X1 i_5717 (.ZN (n_5653), .A (n_7183));
INV_X1 i_5716 (.ZN (n_5652), .A (n_7181));
OAI21_X1 i_5715 (.ZN (n_5651), .A (n_7182), .B1 (n_5653), .B2 (n_5652));
OAI21_X1 i_5714 (.ZN (n_5650), .A (n_5651), .B1 (n_7913), .B2 (n_9037));
INV_X1 i_5713 (.ZN (n_5649), .A (n_5651));
NAND3_X1 i_5712 (.ZN (n_5648), .A1 (n_5649), .A2 (B_imm[14]), .A3 (opt_ipoPP_0));
NAND2_X1 i_5711 (.ZN (n_5647), .A1 (n_5648), .A2 (n_5650));
XNOR2_X1 i_5710 (.ZN (n_5646), .A (n_5647), .B (n_5654));
NAND2_X1 i_5709 (.ZN (n_5645), .A1 (B_imm[31]), .A2 (A_imm[14]));
INV_X1 i_5708 (.ZN (n_5644), .A (n_5645));
INV_X1 i_5707 (.ZN (n_5643), .A (n_7193));
OAI21_X1 i_5706 (.ZN (n_5642), .A (n_7194), .B1 (n_7195), .B2 (n_5643));
OAI21_X1 i_5705 (.ZN (n_5641), .A (n_5642), .B1 (n_9004), .B2 (n_8946));
INV_X1 i_5704 (.ZN (n_5640), .A (n_5642));
NAND3_X1 i_5703 (.ZN (n_5639), .A1 (n_5640), .A2 (B_imm[30]), .A3 (A_imm[15]));
NAND2_X1 i_5702 (.ZN (n_5638), .A1 (n_5639), .A2 (n_5641));
XNOR2_X1 i_5701 (.ZN (n_5637), .A (n_5638), .B (n_5644));
NAND2_X1 i_5700 (.ZN (n_5636), .A1 (A_imm[27]), .A2 (B_imm[18]));
INV_X1 i_5699 (.ZN (n_5635), .A (n_5636));
INV_X1 i_5698 (.ZN (n_5634), .A (n_7177));
INV_X1 i_5697 (.ZN (n_5633), .A (n_7175));
OAI21_X1 i_5696 (.ZN (n_5632), .A (n_7176), .B1 (n_5634), .B2 (n_5633));
INV_X1 i_5695 (.ZN (n_5631), .A (n_7410));
INV_X1 i_5694 (.ZN (n_5630), .A (n_7408));
OAI21_X1 i_5693 (.ZN (n_5629), .A (n_7409), .B1 (n_5631), .B2 (n_5630));
NAND2_X1 i_5692 (.ZN (n_5628), .A1 (n_5632), .A2 (n_5629));
INV_X1 i_5691 (.ZN (n_5627), .A (n_5632));
INV_X1 i_5690 (.ZN (n_5626), .A (n_5629));
NAND2_X1 i_5689 (.ZN (n_5625), .A1 (n_5627), .A2 (n_5626));
NAND2_X1 i_5688 (.ZN (n_5624), .A1 (n_5625), .A2 (n_5628));
XNOR2_X1 i_5687 (.ZN (n_5623), .A (n_5624), .B (n_5635));
NAND2_X1 i_5686 (.ZN (n_5622), .A1 (n_5637), .A2 (n_5623));
INV_X1 i_5685 (.ZN (n_5621), .A (n_5622));
INV_X1 i_5684 (.ZN (n_5620), .A (n_5637));
INV_X1 i_5683 (.ZN (n_5619), .A (n_5623));
NAND2_X1 i_5682 (.ZN (n_5618), .A1 (n_5620), .A2 (n_5619));
INV_X1 i_5681 (.ZN (n_5617), .A (n_5618));
OAI21_X1 i_5680 (.ZN (n_5616), .A (n_5646), .B1 (n_5617), .B2 (n_5621));
INV_X1 i_5679 (.ZN (n_5615), .A (n_5646));
NAND3_X1 i_5678 (.ZN (n_5614), .A1 (n_5618), .A2 (n_5615), .A3 (n_5622));
NAND2_X1 i_5677 (.ZN (n_5613), .A1 (n_7157), .A2 (n_7161));
NAND2_X1 i_5676 (.ZN (n_5612), .A1 (n_5613), .A2 (n_7162));
NAND3_X1 i_5675 (.ZN (n_5611), .A1 (n_5612), .A2 (n_5616), .A3 (n_5614));
NAND2_X1 i_5674 (.ZN (n_5610), .A1 (n_5616), .A2 (n_5614));
NAND3_X1 i_5673 (.ZN (n_5609), .A1 (n_5610), .A2 (n_5613), .A3 (n_7162));
NAND2_X1 i_5672 (.ZN (n_5608), .A1 (A_imm[30]), .A2 (B_imm[15]));
NAND2_X1 i_5671 (.ZN (n_5607), .A1 (n_7104), .A2 (n_7109));
NAND2_X1 i_5670 (.ZN (n_5606), .A1 (B_imm[19]), .A2 (A_imm[26]));
OAI22_X1 i_5669 (.ZN (n_5605), .A1 (n_9021), .A2 (n_8955), .B1 (n_8993), .B2 (n_8892));
NAND4_X1 i_5668 (.ZN (n_5604), .A1 (B_imm[28]), .A2 (B_imm[26]), .A3 (A_imm[19]), .A4 (A_imm[17]));
NAND2_X1 i_5667 (.ZN (n_5603), .A1 (n_5605), .A2 (n_5604));
XNOR2_X1 i_5666 (.ZN (n_5602), .A (n_5603), .B (n_5606));
INV_X1 i_5665 (.ZN (n_5601), .A (n_5602));
NAND3_X1 i_5664 (.ZN (n_5600), .A1 (n_5601), .A2 (n_7106), .A3 (n_5607));
NAND2_X1 i_5663 (.ZN (n_5599), .A1 (n_5607), .A2 (n_7106));
NAND2_X1 i_5662 (.ZN (n_5598), .A1 (n_5599), .A2 (n_5602));
NAND2_X1 i_5661 (.ZN (n_5597), .A1 (n_5600), .A2 (n_5598));
XNOR2_X1 i_5660 (.ZN (n_5596), .A (n_5597), .B (n_5608));
INV_X1 i_5659 (.ZN (n_5595), .A (n_5596));
NAND2_X1 i_5658 (.ZN (n_5594), .A1 (B_imm[20]), .A2 (A_imm[25]));
OAI22_X1 i_5657 (.ZN (n_5593), .A1 (n_8974), .A2 (n_8893), .B1 (n_8958), .B2 (n_8907));
NAND4_X1 i_5656 (.ZN (n_5592), .A1 (B_imm[25]), .A2 (B_imm[22]), .A3 (A_imm[23]), .A4 (A_imm[20]));
NAND2_X1 i_5655 (.ZN (n_5591), .A1 (n_5593), .A2 (n_5592));
XNOR2_X1 i_5654 (.ZN (n_5590), .A (n_5591), .B (n_5594));
NAND2_X1 i_5653 (.ZN (n_5589), .A1 (n_7100), .A2 (n_7097));
NAND2_X1 i_5652 (.ZN (n_5588), .A1 (n_5589), .A2 (n_7098));
NAND2_X1 i_5651 (.ZN (n_5587), .A1 (B_imm[21]), .A2 (A_imm[24]));
OAI22_X1 i_5650 (.ZN (n_5586), .A1 (n_8821), .A2 (n_8906), .B1 (n_8948), .B2 (n_8859));
NAND4_X1 i_5649 (.ZN (n_5585), .A1 (B_imm[23]), .A2 (B_imm[24]), .A3 (A_imm[22]), .A4 (A_imm[21]));
NAND2_X1 i_5648 (.ZN (n_5584), .A1 (n_5586), .A2 (n_5585));
XNOR2_X1 i_5647 (.ZN (n_5583), .A (n_5584), .B (n_5587));
OR2_X1 i_5646 (.ZN (n_5582), .A1 (n_5583), .A2 (n_5588));
NAND2_X1 i_5645 (.ZN (n_5581), .A1 (n_5583), .A2 (n_5588));
NAND3_X1 i_5644 (.ZN (n_5580), .A1 (n_5582), .A2 (n_5581), .A3 (n_5590));
INV_X1 i_5643 (.ZN (n_5579), .A (n_5590));
INV_X1 i_5642 (.ZN (n_5578), .A (n_5582));
INV_X1 i_5641 (.ZN (n_5577), .A (n_5581));
OAI21_X1 i_5640 (.ZN (n_5576), .A (n_5579), .B1 (n_5578), .B2 (n_5577));
NAND2_X1 i_5639 (.ZN (n_5575), .A1 (n_5576), .A2 (n_5580));
NAND2_X1 i_5638 (.ZN (n_5574), .A1 (n_7115), .A2 (n_7153));
NAND2_X1 i_5637 (.ZN (n_5573), .A1 (n_5574), .A2 (n_7118));
NAND2_X1 i_5636 (.ZN (n_5572), .A1 (n_5573), .A2 (n_5575));
NAND4_X1 i_5635 (.ZN (n_5571), .A1 (n_5574), .A2 (n_7118), .A3 (n_5580), .A4 (n_5576));
NAND3_X1 i_5634 (.ZN (n_5570), .A1 (n_5572), .A2 (n_5595), .A3 (n_5571));
NAND2_X1 i_5633 (.ZN (n_5569), .A1 (n_5572), .A2 (n_5571));
NAND2_X1 i_5632 (.ZN (n_5568), .A1 (n_5569), .A2 (n_5596));
NAND2_X1 i_5631 (.ZN (n_5567), .A1 (n_5568), .A2 (n_5570));
NAND3_X1 i_5630 (.ZN (n_5566), .A1 (n_5611), .A2 (n_5567), .A3 (n_5609));
NAND2_X1 i_5629 (.ZN (n_5565), .A1 (n_5611), .A2 (n_5609));
INV_X1 i_5628 (.ZN (n_5564), .A (n_5567));
NAND2_X1 i_5627 (.ZN (n_5563), .A1 (n_5565), .A2 (n_5564));
NAND2_X1 i_5626 (.ZN (n_5562), .A1 (n_5563), .A2 (n_5566));
AOI21_X1 i_5625 (.ZN (n_5561), .A (n_7047), .B1 (n_7006), .B2 (n_7022));
OAI21_X1 i_5624 (.ZN (n_5560), .A (n_5562), .B1 (n_5561), .B2 (n_7003));
INV_X1 i_5623 (.ZN (n_5559), .A (n_5562));
NAND2_X1 i_5622 (.ZN (n_5558), .A1 (n_7005), .A2 (n_7046));
NAND3_X1 i_5621 (.ZN (n_5557), .A1 (n_5558), .A2 (n_5559), .A3 (n_7048));
NAND2_X1 i_5620 (.ZN (n_5556), .A1 (n_7089), .A2 (n_7087));
NAND2_X1 i_5619 (.ZN (n_5555), .A1 (n_5556), .A2 (n_7091));
OAI21_X1 i_5618 (.ZN (n_5554), .A (n_7171), .B1 (n_7165), .B2 (n_7179));
NAND2_X1 i_5617 (.ZN (n_5553), .A1 (n_7188), .A2 (n_7198));
NAND3_X1 i_5616 (.ZN (n_5552), .A1 (n_5554), .A2 (n_7189), .A3 (n_5553));
NAND2_X1 i_5615 (.ZN (n_5551), .A1 (n_5553), .A2 (n_7189));
OAI211_X1 i_5614 (.ZN (n_5550), .A (n_5551), .B (n_7171), .C1 (n_7179), .C2 (n_7165));
NAND3_X1 i_5613 (.ZN (n_5549), .A1 (n_5550), .A2 (n_5555), .A3 (n_5552));
NAND2_X1 i_5612 (.ZN (n_5548), .A1 (n_5550), .A2 (n_5552));
NAND3_X1 i_5611 (.ZN (n_5547), .A1 (n_5548), .A2 (n_7091), .A3 (n_5556));
NAND2_X1 i_5610 (.ZN (n_5546), .A1 (n_5547), .A2 (n_5549));
OAI21_X1 i_5609 (.ZN (n_5545), .A (n_7398), .B1 (n_7393), .B2 (n_7406));
INV_X1 i_5608 (.ZN (n_5544), .A (n_7148));
OAI21_X1 i_5607 (.ZN (n_5543), .A (n_7149), .B1 (n_7150), .B2 (n_5544));
NAND2_X1 i_5606 (.ZN (n_5542), .A1 (A_imm[28]), .A2 (B_imm[17]));
OAI22_X1 i_5605 (.ZN (n_5541), .A1 (n_9006), .A2 (n_8858), .B1 (CLOCK_opt_ipo_n433), .B2 (n_8956));
NAND4_X1 i_5604 (.ZN (n_5540), .A1 (B_imm[29]), .A2 (B_imm[27]), .A3 (A_imm[18]), .A4 (A_imm[16]));
NAND2_X1 i_5603 (.ZN (n_5539), .A1 (n_5541), .A2 (n_5540));
XNOR2_X1 i_5602 (.ZN (n_5538), .A (n_5539), .B (n_5542));
OR2_X1 i_5601 (.ZN (n_5537), .A1 (n_5538), .A2 (n_5543));
NAND2_X1 i_5600 (.ZN (n_5536), .A1 (n_5538), .A2 (n_5543));
NAND3_X1 i_5599 (.ZN (n_5535), .A1 (n_5537), .A2 (n_5545), .A3 (n_5536));
INV_X1 i_5598 (.ZN (n_5534), .A (n_5545));
NAND2_X1 i_5597 (.ZN (n_5533), .A1 (n_5537), .A2 (n_5536));
NAND2_X1 i_5596 (.ZN (n_5532), .A1 (n_5533), .A2 (n_5534));
NAND2_X1 i_5595 (.ZN (n_5531), .A1 (n_5532), .A2 (n_5535));
INV_X1 i_5594 (.ZN (n_5530), .A (n_5531));
NAND2_X1 i_5593 (.ZN (n_5529), .A1 (n_7370), .A2 (n_7411));
NAND2_X1 i_5592 (.ZN (n_5528), .A1 (n_5529), .A2 (n_7371));
NAND2_X1 i_5591 (.ZN (n_5527), .A1 (n_5528), .A2 (n_5530));
NAND3_X1 i_5590 (.ZN (n_5526), .A1 (n_5531), .A2 (n_5529), .A3 (n_7371));
NAND3_X1 i_5589 (.ZN (n_5525), .A1 (n_5546), .A2 (n_5527), .A3 (n_5526));
INV_X1 i_5588 (.ZN (n_5524), .A (n_5546));
NAND2_X1 i_5587 (.ZN (n_5523), .A1 (n_5527), .A2 (n_5526));
NAND2_X1 i_5586 (.ZN (n_5522), .A1 (n_5523), .A2 (n_5524));
NAND2_X1 i_5585 (.ZN (n_5521), .A1 (n_5522), .A2 (n_5525));
NAND2_X1 i_5584 (.ZN (n_5520), .A1 (n_7080), .A2 (n_7053));
NAND2_X1 i_5583 (.ZN (n_5519), .A1 (n_5520), .A2 (n_7083));
NAND2_X1 i_5582 (.ZN (n_5518), .A1 (n_5521), .A2 (n_5519));
NAND4_X1 i_5581 (.ZN (n_5517), .A1 (n_5522), .A2 (n_5525), .A3 (n_7083), .A4 (n_5520));
NAND2_X1 i_5580 (.ZN (n_5516), .A1 (n_7233), .A2 (n_7301));
NAND2_X1 i_5579 (.ZN (n_5515), .A1 (n_5516), .A2 (n_7303));
NAND3_X1 i_5578 (.ZN (n_5514), .A1 (n_5515), .A2 (n_5518), .A3 (n_5517));
NAND2_X1 i_5577 (.ZN (n_5513), .A1 (n_5518), .A2 (n_5517));
INV_X1 i_5576 (.ZN (n_5512), .A (n_5515));
NAND2_X1 i_5575 (.ZN (n_5511), .A1 (n_5513), .A2 (n_5512));
NAND2_X1 i_5574 (.ZN (n_5510), .A1 (n_5511), .A2 (n_5514));
NAND3_X1 i_5573 (.ZN (n_5509), .A1 (n_5560), .A2 (n_5510), .A3 (n_5557));
NAND2_X1 i_5572 (.ZN (n_5508), .A1 (n_5560), .A2 (n_5557));
INV_X1 i_5571 (.ZN (n_5507), .A (n_5510));
NAND2_X1 i_5570 (.ZN (n_5506), .A1 (n_5508), .A2 (n_5507));
NAND4_X2 i_5569 (.ZN (n_5505), .A1 (n_5506), .A2 (n_7200), .A3 (n_5655), .A4 (n_5509));
NAND2_X1 i_5568 (.ZN (n_5504), .A1 (B_imm[26]), .A2 (A_imm[20]));
OAI22_X1 i_5567 (.ZN (n_5503), .A1 (n_9021), .A2 (n_8956), .B1 (n_8860), .B2 (n_8972));
NAND4_X1 i_5566 (.ZN (n_5502), .A1 (B_imm[28]), .A2 (B_imm[20]), .A3 (A_imm[26]), .A4 (A_imm[18]));
NAND2_X1 i_5565 (.ZN (n_5501), .A1 (n_5503), .A2 (n_5502));
XNOR2_X1 i_5564 (.ZN (n_5500), .A (n_5501), .B (n_5504));
INV_X1 i_5563 (.ZN (n_5499), .A (n_5500));
NAND2_X1 i_5562 (.ZN (n_5498), .A1 (B_imm[25]), .A2 (A_imm[21]));
OAI22_X1 i_5561 (.ZN (n_5497), .A1 (n_8829), .A2 (n_9037), .B1 (n_8958), .B2 (n_8767));
NAND4_X1 i_5560 (.ZN (n_5496), .A1 (B_imm[15]), .A2 (B_imm[22]), .A3 (opt_ipoPP_0), .A4 (A_imm[24]));
NAND2_X1 i_5559 (.ZN (n_5495), .A1 (n_5497), .A2 (n_5496));
XNOR2_X1 i_5558 (.ZN (n_5494), .A (n_5495), .B (n_5498));
INV_X1 i_5557 (.ZN (n_5493), .A (n_5494));
NAND2_X1 i_5556 (.ZN (n_5492), .A1 (n_5499), .A2 (n_5493));
INV_X1 i_5555 (.ZN (n_5491), .A (n_5625));
OAI21_X1 i_5554 (.ZN (n_5490), .A (n_5628), .B1 (n_5491), .B2 (n_5635));
INV_X1 i_5553 (.ZN (n_5489), .A (n_5490));
NAND2_X1 i_5552 (.ZN (n_5488), .A1 (n_5500), .A2 (n_5494));
NAND2_X1 i_5551 (.ZN (n_5487), .A1 (n_5488), .A2 (n_5489));
NAND2_X1 i_5550 (.ZN (n_5486), .A1 (A_imm[29]), .A2 (B_imm[18]));
INV_X1 i_5549 (.ZN (n_5485), .A (n_5486));
INV_X1 i_5548 (.ZN (n_5484), .A (n_5504));
INV_X1 i_5547 (.ZN (n_5483), .A (n_5502));
OAI21_X1 i_5546 (.ZN (n_5482), .A (n_5503), .B1 (n_5484), .B2 (n_5483));
OAI21_X1 i_5545 (.ZN (n_5481), .A (n_5482), .B1 (n_9038), .B2 (n_8858));
INV_X1 i_5544 (.ZN (n_5480), .A (n_5482));
NAND3_X1 i_5543 (.ZN (n_5479), .A1 (n_5480), .A2 (B_imm[31]), .A3 (A_imm[16]));
NAND2_X1 i_5542 (.ZN (n_5478), .A1 (n_5479), .A2 (n_5481));
NAND2_X1 i_5541 (.ZN (n_5477), .A1 (n_5478), .A2 (n_5485));
NAND3_X1 i_5540 (.ZN (n_5476), .A1 (n_5479), .A2 (n_5486), .A3 (n_5481));
NAND2_X1 i_5539 (.ZN (n_5475), .A1 (n_5477), .A2 (n_5476));
INV_X1 i_5538 (.ZN (n_5474), .A (n_5542));
INV_X1 i_5537 (.ZN (n_5473), .A (n_5540));
OAI21_X1 i_5536 (.ZN (n_5472), .A (n_5541), .B1 (n_5474), .B2 (n_5473));
INV_X1 i_5535 (.ZN (n_5471), .A (n_5472));
NAND3_X1 i_5534 (.ZN (n_5470), .A1 (n_5471), .A2 (B_imm[17]), .A3 (A_imm[29]));
INV_X1 i_5533 (.ZN (n_5469), .A (n_5470));
OAI21_X1 i_5532 (.ZN (n_5468), .A (n_5472), .B1 (n_8909), .B2 (n_8994));
INV_X1 i_5531 (.ZN (n_5467), .A (n_5468));
NAND2_X1 i_5530 (.ZN (n_5466), .A1 (B_imm[21]), .A2 (A_imm[25]));
OAI22_X1 i_5529 (.ZN (n_5465), .A1 (n_8821), .A2 (n_8907), .B1 (n_8948), .B2 (n_8906));
NAND4_X1 i_5528 (.ZN (n_5464), .A1 (B_imm[23]), .A2 (B_imm[24]), .A3 (A_imm[23]), .A4 (A_imm[22]));
NAND2_X1 i_5527 (.ZN (n_5463), .A1 (n_5465), .A2 (n_5464));
XNOR2_X1 i_5526 (.ZN (n_5462), .A (n_5463), .B (n_5466));
NOR2_X1 i_5525 (.ZN (n_5461), .A1 (n_5467), .A2 (n_5462));
OAI21_X1 i_5524 (.ZN (n_5460), .A (n_5475), .B1 (n_5469), .B2 (n_5461));
NOR2_X1 i_5523 (.ZN (n_5459), .A1 (n_5461), .A2 (n_5469));
NAND3_X1 i_5522 (.ZN (n_5458), .A1 (n_5459), .A2 (n_5477), .A3 (n_5476));
NAND4_X1 i_5521 (.ZN (n_5457), .A1 (n_5458), .A2 (n_5460), .A3 (n_5492), .A4 (n_5487));
NAND2_X1 i_5520 (.ZN (n_5456), .A1 (n_5487), .A2 (n_5492));
NAND2_X1 i_5519 (.ZN (n_5455), .A1 (n_5458), .A2 (n_5460));
NAND2_X1 i_5518 (.ZN (n_5454), .A1 (n_5455), .A2 (n_5456));
INV_X1 i_5517 (.ZN (n_5453), .A (n_5654));
INV_X1 i_5516 (.ZN (n_5452), .A (n_5648));
OAI21_X1 i_5515 (.ZN (n_5451), .A (n_5650), .B1 (n_5452), .B2 (n_5453));
INV_X1 i_5514 (.ZN (n_5450), .A (n_5451));
INV_X1 i_5513 (.ZN (n_5449), .A (n_5639));
OAI21_X1 i_5512 (.ZN (n_5448), .A (n_5641), .B1 (n_5449), .B2 (n_5644));
INV_X1 i_5511 (.ZN (n_5447), .A (n_5448));
NAND3_X1 i_5510 (.ZN (n_5446), .A1 (n_5447), .A2 (B_imm[16]), .A3 (A_imm[30]));
OAI21_X1 i_5509 (.ZN (n_5445), .A (n_5448), .B1 (n_8908), .B2 (n_9005));
NAND2_X1 i_5508 (.ZN (n_5444), .A1 (n_5446), .A2 (n_5445));
NAND2_X1 i_5507 (.ZN (n_5443), .A1 (n_5444), .A2 (n_5450));
INV_X1 i_5506 (.ZN (n_5442), .A (n_5444));
NAND2_X1 i_5505 (.ZN (n_5441), .A1 (n_5442), .A2 (n_5451));
NAND2_X1 i_5504 (.ZN (n_5440), .A1 (n_5441), .A2 (n_5443));
NAND2_X1 i_5503 (.ZN (n_5439), .A1 (n_5545), .A2 (n_5536));
NAND2_X1 i_5502 (.ZN (n_5438), .A1 (n_5537), .A2 (n_5439));
NAND2_X1 i_5501 (.ZN (n_5437), .A1 (n_5440), .A2 (n_5438));
OAI21_X1 i_5500 (.ZN (n_5436), .A (n_5622), .B1 (n_5617), .B2 (n_5646));
NAND4_X1 i_5499 (.ZN (n_5435), .A1 (n_5441), .A2 (n_5443), .A3 (n_5537), .A4 (n_5439));
NAND2_X1 i_5498 (.ZN (n_5434), .A1 (n_5436), .A2 (n_5435));
AOI22_X1 i_5497 (.ZN (n_5433), .A1 (n_5434), .A2 (n_5437), .B1 (n_5457), .B2 (n_5454));
INV_X1 i_5496 (.ZN (n_5432), .A (n_5433));
NAND2_X1 i_5495 (.ZN (n_5431), .A1 (n_5454), .A2 (n_5457));
INV_X1 i_5494 (.ZN (n_5430), .A (n_5431));
NAND3_X1 i_5493 (.ZN (n_5429), .A1 (n_5434), .A2 (n_5430), .A3 (n_5437));
INV_X1 i_5492 (.ZN (n_5428), .A (n_5446));
INV_X1 i_5491 (.ZN (n_5427), .A (n_5594));
INV_X1 i_5490 (.ZN (n_5426), .A (n_5592));
OAI21_X1 i_5489 (.ZN (n_5425), .A (n_5593), .B1 (n_5427), .B2 (n_5426));
INV_X1 i_5488 (.ZN (n_5424), .A (n_5425));
INV_X1 i_5487 (.ZN (n_5423), .A (n_5587));
INV_X1 i_5486 (.ZN (n_5422), .A (n_5585));
OAI21_X1 i_5485 (.ZN (n_5421), .A (n_5586), .B1 (n_5423), .B2 (n_5422));
OAI21_X1 i_5484 (.ZN (n_5420), .A (n_5421), .B1 (n_8525), .B2 (n_7912));
INV_X1 i_5483 (.ZN (n_5419), .A (n_5421));
NAND3_X1 i_5482 (.ZN (n_5418), .A1 (n_5419), .A2 (B_imm[19]), .A3 (A_imm[27]));
NAND2_X1 i_5481 (.ZN (n_5417), .A1 (n_5418), .A2 (n_5420));
NAND2_X1 i_5480 (.ZN (n_5416), .A1 (n_5417), .A2 (n_5424));
NAND3_X1 i_5479 (.ZN (n_5415), .A1 (n_5418), .A2 (n_5425), .A3 (n_5420));
NAND2_X1 i_5478 (.ZN (n_5414), .A1 (n_5416), .A2 (n_5415));
NAND2_X1 i_5477 (.ZN (n_5413), .A1 (A_imm[28]), .A2 (B_imm[18]));
OAI22_X1 i_5476 (.ZN (n_5412), .A1 (n_9006), .A2 (n_8955), .B1 (CLOCK_opt_ipo_n433), .B2 (n_8892));
NAND4_X1 i_5475 (.ZN (n_5411), .A1 (B_imm[29]), .A2 (B_imm[27]), .A3 (A_imm[19]), .A4 (A_imm[17]));
NAND2_X1 i_5474 (.ZN (n_5410), .A1 (n_5412), .A2 (n_5411));
XNOR2_X1 i_5473 (.ZN (n_5409), .A (n_5410), .B (n_5413));
INV_X1 i_5472 (.ZN (n_5408), .A (n_5409));
NAND2_X1 i_5471 (.ZN (n_5407), .A1 (n_5414), .A2 (n_5408));
NAND2_X1 i_5470 (.ZN (n_5406), .A1 (n_5604), .A2 (n_5606));
NAND2_X1 i_5469 (.ZN (n_5405), .A1 (n_5406), .A2 (n_5605));
INV_X1 i_5468 (.ZN (n_5404), .A (n_5405));
OAI22_X1 i_5467 (.ZN (n_5403), .A1 (n_9038), .A2 (n_8946), .B1 (n_9004), .B2 (n_8858));
NAND4_X1 i_5466 (.ZN (n_5402), .A1 (B_imm[31]), .A2 (B_imm[30]), .A3 (A_imm[16]), .A4 (A_imm[15]));
NAND2_X1 i_5465 (.ZN (n_5401), .A1 (n_5403), .A2 (n_5402));
XNOR2_X1 i_5464 (.ZN (n_5400), .A (n_5401), .B (n_5404));
NAND3_X1 i_5463 (.ZN (n_5399), .A1 (n_5416), .A2 (n_5409), .A3 (n_5415));
NAND2_X1 i_5462 (.ZN (n_5398), .A1 (n_5400), .A2 (n_5399));
NAND2_X1 i_5461 (.ZN (n_5397), .A1 (n_5398), .A2 (n_5407));
OAI211_X1 i_5460 (.ZN (n_5396), .A (n_5397), .B (n_5445), .C1 (n_5450), .C2 (n_5428));
OAI21_X1 i_5459 (.ZN (n_5395), .A (n_5445), .B1 (n_5428), .B2 (n_5450));
NAND3_X1 i_5458 (.ZN (n_5394), .A1 (n_5395), .A2 (n_5407), .A3 (n_5398));
NAND2_X1 i_5457 (.ZN (n_5393), .A1 (n_5394), .A2 (n_5396));
INV_X1 i_5456 (.ZN (n_5392), .A (n_5393));
NAND2_X1 i_5455 (.ZN (n_5391), .A1 (n_5411), .A2 (n_5413));
NAND2_X1 i_5454 (.ZN (n_5390), .A1 (n_5391), .A2 (n_5412));
INV_X1 i_5453 (.ZN (n_5389), .A (n_5390));
NAND2_X1 i_5452 (.ZN (n_5388), .A1 (B_imm[25]), .A2 (A_imm[22]));
INV_X1 i_5451 (.ZN (n_5387), .A (n_5388));
OAI22_X1 i_5450 (.ZN (n_5386), .A1 (n_8958), .A2 (n_8794), .B1 (n_8957), .B2 (n_8972));
NAND4_X1 i_5449 (.ZN (n_5385), .A1 (B_imm[22]), .A2 (B_imm[21]), .A3 (A_imm[26]), .A4 (A_imm[25]));
NAND2_X1 i_5448 (.ZN (n_5384), .A1 (n_5386), .A2 (n_5385));
XNOR2_X1 i_5447 (.ZN (n_5383), .A (n_5384), .B (n_5387));
NAND2_X1 i_5446 (.ZN (n_5382), .A1 (n_5383), .A2 (n_5389));
OR2_X1 i_5445 (.ZN (n_5381), .A1 (n_5383), .A2 (n_5389));
NAND2_X1 i_5444 (.ZN (n_5380), .A1 (n_5381), .A2 (n_5382));
NAND2_X1 i_5443 (.ZN (n_5379), .A1 (B_imm[23]), .A2 (A_imm[24]));
OAI22_X1 i_5442 (.ZN (n_5378), .A1 (n_8948), .A2 (n_8907), .B1 (n_9037), .B2 (n_8908));
NAND4_X1 i_5441 (.ZN (n_5377), .A1 (B_imm[24]), .A2 (A_imm[31]), .A3 (B_imm[16]), .A4 (A_imm[23]));
NAND2_X1 i_5440 (.ZN (n_5376), .A1 (n_5378), .A2 (n_5377));
XNOR2_X1 i_5439 (.ZN (n_5375), .A (n_5376), .B (n_5379));
XNOR2_X1 i_5438 (.ZN (n_5374), .A (n_5380), .B (n_5375));
NAND2_X1 i_5437 (.ZN (n_5373), .A1 (n_5392), .A2 (n_5374));
INV_X1 i_5436 (.ZN (n_5372), .A (n_5374));
NAND2_X1 i_5435 (.ZN (n_5371), .A1 (n_5393), .A2 (n_5372));
NAND2_X1 i_5434 (.ZN (n_5370), .A1 (n_5373), .A2 (n_5371));
NAND2_X1 i_5433 (.ZN (n_5369), .A1 (n_5370), .A2 (n_5429));
NAND2_X1 i_5432 (.ZN (n_5368), .A1 (n_5369), .A2 (n_5432));
INV_X1 i_5431 (.ZN (n_5367), .A (n_5498));
INV_X1 i_5430 (.ZN (n_5366), .A (n_5496));
OAI21_X1 i_5429 (.ZN (n_5365), .A (n_5497), .B1 (n_5367), .B2 (n_5366));
OAI21_X1 i_5428 (.ZN (n_5364), .A (n_5365), .B1 (n_8860), .B2 (n_7912));
NAND2_X1 i_5427 (.ZN (n_5363), .A1 (B_imm[30]), .A2 (A_imm[17]));
INV_X1 i_5426 (.ZN (n_5362), .A (n_5363));
INV_X1 i_5425 (.ZN (n_5361), .A (n_5365));
NAND3_X1 i_5424 (.ZN (n_5360), .A1 (n_5361), .A2 (B_imm[20]), .A3 (A_imm[27]));
INV_X1 i_5423 (.ZN (n_5359), .A (n_5360));
OAI21_X1 i_5422 (.ZN (n_5358), .A (n_5364), .B1 (n_5359), .B2 (n_5362));
OAI22_X1 i_5421 (.ZN (n_5357), .A1 (n_9020), .A2 (n_8525), .B1 (n_9006), .B2 (n_8956));
NAND2_X1 i_5420 (.ZN (n_5356), .A1 (n_5464), .A2 (n_5466));
NAND2_X1 i_5419 (.ZN (n_5355), .A1 (n_5356), .A2 (n_5465));
INV_X1 i_5418 (.ZN (n_5354), .A (n_5355));
NAND4_X1 i_5417 (.ZN (n_5353), .A1 (A_imm[28]), .A2 (B_imm[29]), .A3 (B_imm[19]), .A4 (A_imm[18]));
INV_X1 i_5416 (.ZN (n_5352), .A (n_5353));
OAI21_X1 i_5415 (.ZN (n_5351), .A (n_5357), .B1 (n_5354), .B2 (n_5352));
NAND2_X1 i_5414 (.ZN (n_5350), .A1 (B_imm[28]), .A2 (A_imm[20]));
OAI22_X1 i_5413 (.ZN (n_5349), .A1 (n_8974), .A2 (n_8907), .B1 (n_8958), .B2 (n_8972));
NAND4_X1 i_5412 (.ZN (n_5348), .A1 (B_imm[25]), .A2 (B_imm[22]), .A3 (A_imm[26]), .A4 (A_imm[23]));
NAND2_X1 i_5411 (.ZN (n_5347), .A1 (n_5349), .A2 (n_5348));
XNOR2_X1 i_5410 (.ZN (n_5346), .A (n_5347), .B (n_5350));
NAND2_X1 i_5409 (.ZN (n_5345), .A1 (n_5346), .A2 (n_5351));
OR2_X1 i_5408 (.ZN (n_5344), .A1 (n_5346), .A2 (n_5351));
NAND2_X1 i_5407 (.ZN (n_5343), .A1 (n_5344), .A2 (n_5345));
NAND2_X1 i_5406 (.ZN (n_5342), .A1 (n_5343), .A2 (n_5358));
OR2_X1 i_5405 (.ZN (n_5341), .A1 (n_5343), .A2 (n_5358));
NAND2_X1 i_5404 (.ZN (n_5340), .A1 (n_5458), .A2 (n_5456));
NAND2_X1 i_5403 (.ZN (n_5339), .A1 (n_5340), .A2 (n_5460));
NAND3_X1 i_5402 (.ZN (n_5338), .A1 (n_5339), .A2 (n_5342), .A3 (n_5341));
NAND2_X1 i_5401 (.ZN (n_5337), .A1 (n_5341), .A2 (n_5342));
INV_X1 i_5400 (.ZN (n_5336), .A (n_5339));
NAND2_X1 i_5399 (.ZN (n_5335), .A1 (n_5337), .A2 (n_5336));
INV_X1 i_5398 (.ZN (n_5334), .A (n_5479));
OAI21_X1 i_5397 (.ZN (n_5333), .A (n_5481), .B1 (n_5334), .B2 (n_5485));
NAND2_X1 i_5396 (.ZN (n_5332), .A1 (A_imm[30]), .A2 (B_imm[18]));
INV_X1 i_5395 (.ZN (n_5331), .A (n_5332));
NAND2_X1 i_5394 (.ZN (n_5330), .A1 (B_imm[29]), .A2 (A_imm[19]));
INV_X1 i_5393 (.ZN (n_5329), .A (n_5330));
OAI22_X1 i_5392 (.ZN (n_5328), .A1 (CLOCK_opt_ipo_n433), .A2 (n_8859), .B1 (n_8993), .B2 (n_8906));
NAND4_X1 i_5391 (.ZN (n_5327), .A1 (B_imm[27]), .A2 (B_imm[26]), .A3 (A_imm[22]), .A4 (A_imm[21]));
NAND2_X1 i_5390 (.ZN (n_5326), .A1 (n_5328), .A2 (n_5327));
XNOR2_X1 i_5389 (.ZN (n_5325), .A (n_5326), .B (n_5329));
OR2_X1 i_5388 (.ZN (n_5324), .A1 (n_5325), .A2 (n_5331));
NAND2_X1 i_5387 (.ZN (n_5323), .A1 (n_5325), .A2 (n_5331));
NAND2_X1 i_5386 (.ZN (n_5322), .A1 (n_5324), .A2 (n_5323));
XNOR2_X1 i_5385 (.ZN (n_5321), .A (n_5322), .B (n_5333));
NAND3_X1 i_5384 (.ZN (n_5320), .A1 (n_5335), .A2 (n_5338), .A3 (n_5321));
INV_X1 i_5383 (.ZN (n_5319), .A (n_5320));
AOI21_X1 i_5382 (.ZN (n_5318), .A (n_5321), .B1 (n_5335), .B2 (n_5338));
NAND2_X1 i_5381 (.ZN (n_5317), .A1 (n_5418), .A2 (n_5425));
NAND2_X1 i_5380 (.ZN (n_5316), .A1 (n_5317), .A2 (n_5420));
INV_X1 i_5379 (.ZN (n_5315), .A (n_5316));
NAND2_X1 i_5378 (.ZN (n_5314), .A1 (B_imm[27]), .A2 (A_imm[20]));
OAI22_X1 i_5377 (.ZN (n_5313), .A1 (n_9021), .A2 (n_8892), .B1 (n_8993), .B2 (n_8859));
NAND4_X1 i_5376 (.ZN (n_5312), .A1 (B_imm[28]), .A2 (B_imm[26]), .A3 (A_imm[21]), .A4 (A_imm[19]));
NAND2_X1 i_5375 (.ZN (n_5311), .A1 (n_5313), .A2 (n_5312));
XNOR2_X1 i_5374 (.ZN (n_5310), .A (n_5311), .B (n_5314));
INV_X1 i_5373 (.ZN (n_5309), .A (n_5310));
NAND2_X1 i_5372 (.ZN (n_5308), .A1 (n_5315), .A2 (n_5309));
INV_X1 i_5371 (.ZN (n_5307), .A (n_5308));
NAND2_X1 i_5370 (.ZN (n_5306), .A1 (n_5316), .A2 (n_5310));
INV_X1 i_5369 (.ZN (n_5305), .A (n_5306));
OAI211_X1 i_5368 (.ZN (n_5304), .A (B_imm[17]), .B (A_imm[30]), .C1 (n_5307), .C2 (n_5305));
NAND2_X1 i_5367 (.ZN (n_5303), .A1 (A_imm[30]), .A2 (B_imm[17]));
NAND3_X1 i_5366 (.ZN (n_5302), .A1 (n_5308), .A2 (n_5303), .A3 (n_5306));
NAND2_X1 i_5365 (.ZN (n_5301), .A1 (n_5304), .A2 (n_5302));
INV_X1 i_5364 (.ZN (n_5300), .A (n_5608));
NAND2_X1 i_5363 (.ZN (n_5299), .A1 (n_5598), .A2 (n_5300));
NAND2_X1 i_5362 (.ZN (n_5298), .A1 (n_5299), .A2 (n_5600));
NAND2_X1 i_5361 (.ZN (n_5297), .A1 (n_5581), .A2 (n_5579));
NAND2_X1 i_5360 (.ZN (n_5296), .A1 (n_5582), .A2 (n_5297));
NAND2_X1 i_5359 (.ZN (n_5295), .A1 (n_5298), .A2 (n_5296));
NAND4_X1 i_5358 (.ZN (n_5294), .A1 (n_5299), .A2 (n_5600), .A3 (n_5582), .A4 (n_5297));
NAND2_X1 i_5357 (.ZN (n_5293), .A1 (n_5470), .A2 (n_5468));
XNOR2_X1 i_5356 (.ZN (n_5292), .A (n_5293), .B (n_5462));
INV_X1 i_5355 (.ZN (n_5291), .A (n_5292));
NAND2_X1 i_5354 (.ZN (n_5290), .A1 (n_5294), .A2 (n_5291));
NAND2_X1 i_5353 (.ZN (n_5289), .A1 (n_5290), .A2 (n_5295));
NAND2_X1 i_5352 (.ZN (n_5288), .A1 (n_5289), .A2 (n_5301));
NAND4_X1 i_5351 (.ZN (n_5287), .A1 (n_5290), .A2 (n_5304), .A3 (n_5302), .A4 (n_5295));
NAND2_X1 i_5350 (.ZN (n_5286), .A1 (n_5360), .A2 (n_5364));
XNOR2_X1 i_5349 (.ZN (n_5285), .A (n_5286), .B (n_5362));
INV_X1 i_5348 (.ZN (n_5284), .A (n_5402));
OAI21_X1 i_5347 (.ZN (n_5283), .A (n_5403), .B1 (n_5404), .B2 (n_5284));
INV_X1 i_5346 (.ZN (n_5282), .A (n_5283));
NAND2_X1 i_5345 (.ZN (n_5281), .A1 (n_5357), .A2 (n_5353));
XNOR2_X1 i_5344 (.ZN (n_5280), .A (n_5281), .B (n_5354));
NAND2_X1 i_5343 (.ZN (n_5279), .A1 (n_5280), .A2 (n_5282));
OR2_X1 i_5342 (.ZN (n_5278), .A1 (n_5280), .A2 (n_5282));
NAND2_X1 i_5341 (.ZN (n_5277), .A1 (n_5278), .A2 (n_5279));
XNOR2_X1 i_5340 (.ZN (n_5276), .A (n_5277), .B (n_5285));
NAND2_X1 i_5339 (.ZN (n_5275), .A1 (n_5276), .A2 (n_5287));
NAND2_X1 i_5338 (.ZN (n_5274), .A1 (n_5275), .A2 (n_5288));
OAI21_X1 i_5337 (.ZN (n_5273), .A (n_5274), .B1 (n_5319), .B2 (n_5318));
INV_X1 i_5336 (.ZN (n_5272), .A (n_5318));
NAND4_X1 i_5335 (.ZN (n_5271), .A1 (n_5272), .A2 (n_5320), .A3 (n_5288), .A4 (n_5275));
NAND3_X1 i_5334 (.ZN (n_5270), .A1 (n_5368), .A2 (n_5273), .A3 (n_5271));
NAND2_X1 i_5333 (.ZN (n_5269), .A1 (n_5273), .A2 (n_5271));
NAND3_X1 i_5332 (.ZN (n_5268), .A1 (n_5269), .A2 (n_5432), .A3 (n_5369));
NAND2_X1 i_5331 (.ZN (n_5267), .A1 (n_5268), .A2 (n_5270));
NAND2_X1 i_5330 (.ZN (n_5266), .A1 (n_5278), .A2 (n_5285));
NAND2_X1 i_5329 (.ZN (n_5265), .A1 (n_5266), .A2 (n_5279));
NAND2_X1 i_5328 (.ZN (n_5264), .A1 (B_imm[23]), .A2 (A_imm[25]));
INV_X1 i_5327 (.ZN (n_5263), .A (n_5264));
OAI22_X1 i_5326 (.ZN (n_5262), .A1 (n_8948), .A2 (n_8767), .B1 (n_9037), .B2 (n_8909));
NAND4_X1 i_5325 (.ZN (n_5261), .A1 (B_imm[24]), .A2 (A_imm[31]), .A3 (B_imm[17]), .A4 (A_imm[24]));
NAND2_X1 i_5324 (.ZN (n_5260), .A1 (n_5262), .A2 (n_5261));
XNOR2_X1 i_5323 (.ZN (n_5259), .A (n_5260), .B (n_5263));
INV_X1 i_5322 (.ZN (n_5258), .A (n_5314));
INV_X1 i_5321 (.ZN (n_5257), .A (n_5312));
OAI21_X1 i_5320 (.ZN (n_5256), .A (n_5313), .B1 (n_5258), .B2 (n_5257));
OAI21_X1 i_5319 (.ZN (n_5255), .A (n_5256), .B1 (n_8525), .B2 (n_8994));
INV_X1 i_5318 (.ZN (n_5254), .A (n_5256));
NAND3_X1 i_5317 (.ZN (n_5253), .A1 (n_5254), .A2 (B_imm[19]), .A3 (A_imm[29]));
NAND2_X1 i_5316 (.ZN (n_5252), .A1 (n_5253), .A2 (n_5255));
XNOR2_X1 i_5315 (.ZN (n_5251), .A (n_5252), .B (n_5259));
OAI21_X1 i_5314 (.ZN (n_5250), .A (n_5308), .B1 (n_5305), .B2 (n_5303));
NAND2_X1 i_5313 (.ZN (n_5249), .A1 (n_5250), .A2 (n_5251));
OR2_X1 i_5312 (.ZN (n_5248), .A1 (n_5251), .A2 (n_5250));
NAND2_X1 i_5311 (.ZN (n_5247), .A1 (n_5248), .A2 (n_5249));
XNOR2_X1 i_5310 (.ZN (n_5246), .A (n_5247), .B (n_5265));
INV_X1 i_5309 (.ZN (n_5245), .A (n_5375));
NAND2_X1 i_5308 (.ZN (n_5244), .A1 (n_5381), .A2 (n_5245));
NAND2_X1 i_5307 (.ZN (n_5243), .A1 (B_imm[31]), .A2 (A_imm[17]));
OAI22_X1 i_5306 (.ZN (n_5242), .A1 (n_9004), .A2 (n_8956), .B1 (n_7912), .B2 (n_8957));
NAND4_X1 i_5305 (.ZN (n_5241), .A1 (B_imm[30]), .A2 (A_imm[27]), .A3 (B_imm[21]), .A4 (A_imm[18]));
NAND2_X1 i_5304 (.ZN (n_5240), .A1 (n_5242), .A2 (n_5241));
XNOR2_X1 i_5303 (.ZN (n_5239), .A (n_5240), .B (n_5243));
INV_X1 i_5302 (.ZN (n_5238), .A (n_5239));
INV_X1 i_5301 (.ZN (n_5237), .A (n_5385));
OAI21_X1 i_5300 (.ZN (n_5236), .A (n_5386), .B1 (n_5387), .B2 (n_5237));
INV_X1 i_5299 (.ZN (n_5235), .A (n_5236));
INV_X1 i_5298 (.ZN (n_5234), .A (n_5379));
INV_X1 i_5297 (.ZN (n_5233), .A (n_5377));
OAI21_X1 i_5296 (.ZN (n_5232), .A (n_5378), .B1 (n_5234), .B2 (n_5233));
OAI21_X1 i_5295 (.ZN (n_5231), .A (n_5232), .B1 (n_8860), .B2 (n_9020));
INV_X1 i_5294 (.ZN (n_5230), .A (n_5232));
NAND3_X1 i_5293 (.ZN (n_5229), .A1 (n_5230), .A2 (B_imm[20]), .A3 (A_imm[28]));
NAND2_X1 i_5292 (.ZN (n_5228), .A1 (n_5229), .A2 (n_5231));
XNOR2_X1 i_5291 (.ZN (n_5227), .A (n_5228), .B (n_5235));
NAND2_X1 i_5290 (.ZN (n_5226), .A1 (n_5227), .A2 (n_5238));
OR2_X1 i_5289 (.ZN (n_5225), .A1 (n_5227), .A2 (n_5238));
NAND4_X1 i_5288 (.ZN (n_5224), .A1 (n_5225), .A2 (n_5382), .A3 (n_5244), .A4 (n_5226));
NAND2_X1 i_5287 (.ZN (n_5223), .A1 (n_5244), .A2 (n_5382));
NAND2_X1 i_5286 (.ZN (n_5222), .A1 (n_5225), .A2 (n_5226));
NAND2_X1 i_5285 (.ZN (n_5221), .A1 (n_5222), .A2 (n_5223));
NAND2_X1 i_5284 (.ZN (n_5220), .A1 (n_5221), .A2 (n_5224));
NAND2_X1 i_5283 (.ZN (n_5219), .A1 (n_5372), .A2 (n_5394));
NAND2_X1 i_5282 (.ZN (n_5218), .A1 (n_5219), .A2 (n_5396));
NAND2_X1 i_5281 (.ZN (n_5217), .A1 (n_5218), .A2 (n_5220));
NAND4_X1 i_5280 (.ZN (n_5216), .A1 (n_5219), .A2 (n_5396), .A3 (n_5224), .A4 (n_5221));
NAND3_X1 i_5279 (.ZN (n_5215), .A1 (n_5246), .A2 (n_5217), .A3 (n_5216));
INV_X1 i_5278 (.ZN (n_5214), .A (n_5246));
NAND2_X1 i_5277 (.ZN (n_5213), .A1 (n_5217), .A2 (n_5216));
NAND2_X1 i_5276 (.ZN (n_5212), .A1 (n_5213), .A2 (n_5214));
NAND3_X1 i_5275 (.ZN (n_5211), .A1 (n_5276), .A2 (n_5288), .A3 (n_5287));
INV_X1 i_5274 (.ZN (n_5210), .A (n_5276));
NAND2_X1 i_5273 (.ZN (n_5209), .A1 (n_5288), .A2 (n_5287));
NAND2_X1 i_5272 (.ZN (n_5208), .A1 (n_5209), .A2 (n_5210));
NAND2_X1 i_5271 (.ZN (n_5207), .A1 (n_5492), .A2 (n_5488));
XNOR2_X1 i_5270 (.ZN (n_5206), .A (n_5207), .B (n_5489));
NAND2_X1 i_5269 (.ZN (n_5205), .A1 (n_5550), .A2 (n_5555));
NAND2_X1 i_5268 (.ZN (n_5204), .A1 (n_5205), .A2 (n_5552));
NAND2_X1 i_5267 (.ZN (n_5203), .A1 (n_5204), .A2 (n_5206));
INV_X1 i_5266 (.ZN (n_5202), .A (n_5206));
NAND3_X1 i_5265 (.ZN (n_5201), .A1 (n_5205), .A2 (n_5202), .A3 (n_5552));
NAND3_X1 i_5264 (.ZN (n_5200), .A1 (n_5295), .A2 (n_5294), .A3 (n_5291));
NAND2_X1 i_5263 (.ZN (n_5199), .A1 (n_5295), .A2 (n_5294));
NAND2_X1 i_5262 (.ZN (n_5198), .A1 (n_5199), .A2 (n_5292));
NAND2_X1 i_5261 (.ZN (n_5197), .A1 (n_5198), .A2 (n_5200));
INV_X1 i_5260 (.ZN (n_5196), .A (n_5197));
NAND2_X1 i_5259 (.ZN (n_5195), .A1 (n_5196), .A2 (n_5201));
NAND2_X1 i_5258 (.ZN (n_5194), .A1 (n_5195), .A2 (n_5203));
NAND3_X1 i_5257 (.ZN (n_5193), .A1 (n_5194), .A2 (n_5211), .A3 (n_5208));
NAND2_X1 i_5256 (.ZN (n_5192), .A1 (n_5208), .A2 (n_5211));
NAND3_X1 i_5255 (.ZN (n_5191), .A1 (n_5192), .A2 (n_5203), .A3 (n_5195));
NAND2_X1 i_5254 (.ZN (n_5190), .A1 (n_5595), .A2 (n_5571));
INV_X1 i_5253 (.ZN (n_5189), .A (n_5400));
NAND3_X1 i_5252 (.ZN (n_5188), .A1 (n_5407), .A2 (n_5189), .A3 (n_5399));
INV_X1 i_5251 (.ZN (n_5187), .A (n_5188));
AOI21_X1 i_5250 (.ZN (n_5186), .A (n_5189), .B1 (n_5407), .B2 (n_5399));
NOR2_X1 i_5249 (.ZN (n_5185), .A1 (n_5187), .A2 (n_5186));
AOI21_X1 i_5248 (.ZN (n_5184), .A (n_5185), .B1 (n_5190), .B2 (n_5572));
INV_X1 i_5247 (.ZN (n_5183), .A (n_5184));
NAND3_X1 i_5246 (.ZN (n_5182), .A1 (n_5190), .A2 (n_5572), .A3 (n_5185));
NAND3_X1 i_5245 (.ZN (n_5181), .A1 (n_5547), .A2 (n_5526), .A3 (n_5549));
NAND2_X1 i_5244 (.ZN (n_5180), .A1 (n_5181), .A2 (n_5527));
NAND2_X1 i_5243 (.ZN (n_5179), .A1 (n_5180), .A2 (n_5182));
NAND2_X1 i_5242 (.ZN (n_5178), .A1 (n_5179), .A2 (n_5183));
NAND2_X1 i_5241 (.ZN (n_5177), .A1 (n_5178), .A2 (n_5191));
NAND2_X1 i_5240 (.ZN (n_5176), .A1 (n_5177), .A2 (n_5193));
NAND3_X1 i_5239 (.ZN (n_5175), .A1 (n_5176), .A2 (n_5215), .A3 (n_5212));
NAND2_X1 i_5238 (.ZN (n_5174), .A1 (n_5212), .A2 (n_5215));
NAND3_X1 i_5237 (.ZN (n_5173), .A1 (n_5174), .A2 (n_5177), .A3 (n_5193));
NAND3_X1 i_5236 (.ZN (n_5172), .A1 (n_5175), .A2 (n_5267), .A3 (n_5173));
INV_X1 i_5235 (.ZN (n_5171), .A (n_5267));
AOI21_X1 i_5234 (.ZN (n_5170), .A (n_5174), .B1 (n_5177), .B2 (n_5193));
INV_X1 i_5233 (.ZN (n_5169), .A (n_5173));
OAI21_X1 i_5232 (.ZN (n_5168), .A (n_5171), .B1 (n_5170), .B2 (n_5169));
NAND3_X1 i_5231 (.ZN (n_5167), .A1 (n_5432), .A2 (n_5370), .A3 (n_5429));
INV_X1 i_5230 (.ZN (n_5166), .A (n_5429));
INV_X1 i_5229 (.ZN (n_5165), .A (n_5370));
OAI21_X1 i_5228 (.ZN (n_5164), .A (n_5165), .B1 (n_5166), .B2 (n_5433));
NAND3_X1 i_5227 (.ZN (n_5163), .A1 (n_5203), .A2 (n_5197), .A3 (n_5201));
NAND2_X1 i_5226 (.ZN (n_5162), .A1 (n_5203), .A2 (n_5201));
NAND2_X1 i_5225 (.ZN (n_5161), .A1 (n_5162), .A2 (n_5196));
NAND2_X1 i_5224 (.ZN (n_5160), .A1 (n_5161), .A2 (n_5163));
AOI21_X1 i_5223 (.ZN (n_5159), .A (n_5436), .B1 (n_5437), .B2 (n_5435));
INV_X1 i_5222 (.ZN (n_5158), .A (n_5159));
NAND3_X1 i_5221 (.ZN (n_5157), .A1 (n_5437), .A2 (n_5436), .A3 (n_5435));
NAND3_X1 i_5220 (.ZN (n_5156), .A1 (n_5160), .A2 (n_5158), .A3 (n_5157));
NAND2_X1 i_5219 (.ZN (n_5155), .A1 (n_5158), .A2 (n_5157));
NAND3_X1 i_5218 (.ZN (n_5154), .A1 (n_5155), .A2 (n_5161), .A3 (n_5163));
NAND3_X1 i_5217 (.ZN (n_5153), .A1 (n_5180), .A2 (n_5183), .A3 (n_5182));
INV_X1 i_5216 (.ZN (n_5152), .A (n_5182));
OAI211_X1 i_5215 (.ZN (n_5151), .A (n_5527), .B (n_5181), .C1 (n_5152), .C2 (n_5184));
NAND3_X1 i_5214 (.ZN (n_5150), .A1 (n_5154), .A2 (n_5151), .A3 (n_5153));
NAND2_X1 i_5213 (.ZN (n_5149), .A1 (n_5150), .A2 (n_5156));
NAND3_X1 i_5212 (.ZN (n_5148), .A1 (n_5149), .A2 (n_5167), .A3 (n_5164));
NAND2_X1 i_5211 (.ZN (n_5147), .A1 (n_5167), .A2 (n_5164));
NAND3_X1 i_5210 (.ZN (n_5146), .A1 (n_5150), .A2 (n_5147), .A3 (n_5156));
NAND3_X1 i_5209 (.ZN (n_5145), .A1 (n_5178), .A2 (n_5191), .A3 (n_5193));
NAND2_X1 i_5208 (.ZN (n_5144), .A1 (n_5191), .A2 (n_5193));
NAND3_X1 i_5207 (.ZN (n_5143), .A1 (n_5144), .A2 (n_5183), .A3 (n_5179));
NAND2_X1 i_5206 (.ZN (n_5142), .A1 (n_5143), .A2 (n_5145));
INV_X1 i_5205 (.ZN (n_5141), .A (n_5142));
NAND2_X1 i_5204 (.ZN (n_5140), .A1 (n_5141), .A2 (n_5146));
NAND4_X2 i_5203 (.ZN (n_5139), .A1 (n_5168), .A2 (n_5172), .A3 (n_5148), .A4 (n_5140));
NAND3_X1 i_5202 (.ZN (n_5138), .A1 (n_5148), .A2 (n_5142), .A3 (n_5146));
AOI21_X1 i_5201 (.ZN (n_5137), .A (n_5147), .B1 (n_5150), .B2 (n_5156));
INV_X1 i_5200 (.ZN (n_5136), .A (n_5146));
OAI21_X1 i_5199 (.ZN (n_5135), .A (n_5141), .B1 (n_5137), .B2 (n_5136));
NAND2_X1 i_5198 (.ZN (n_5134), .A1 (n_5515), .A2 (n_5517));
NAND2_X1 i_5197 (.ZN (n_5133), .A1 (n_5134), .A2 (n_5518));
NAND2_X1 i_5196 (.ZN (n_5132), .A1 (n_5564), .A2 (n_5609));
NAND2_X1 i_5195 (.ZN (n_5131), .A1 (n_5132), .A2 (n_5611));
NAND2_X1 i_5194 (.ZN (n_5130), .A1 (n_5133), .A2 (n_5131));
NAND4_X1 i_5193 (.ZN (n_5129), .A1 (n_5134), .A2 (n_5611), .A3 (n_5518), .A4 (n_5132));
NAND2_X1 i_5192 (.ZN (n_5128), .A1 (n_5151), .A2 (n_5153));
NAND3_X1 i_5191 (.ZN (n_5127), .A1 (n_5156), .A2 (n_5128), .A3 (n_5154));
INV_X1 i_5190 (.ZN (n_5126), .A (n_5128));
NAND2_X1 i_5189 (.ZN (n_5125), .A1 (n_5156), .A2 (n_5154));
NAND2_X1 i_5188 (.ZN (n_5124), .A1 (n_5125), .A2 (n_5126));
NAND2_X1 i_5187 (.ZN (n_5123), .A1 (n_5124), .A2 (n_5127));
NAND2_X1 i_5186 (.ZN (n_5122), .A1 (n_5123), .A2 (n_5129));
NAND4_X2 i_5185 (.ZN (n_5121), .A1 (n_5135), .A2 (n_5138), .A3 (n_5122), .A4 (n_5130));
NAND3_X1 i_5184 (.ZN (n_5120), .A1 (n_5123), .A2 (n_5130), .A3 (n_5129));
INV_X1 i_5183 (.ZN (n_5119), .A (n_5123));
NAND2_X1 i_5182 (.ZN (n_5118), .A1 (n_5130), .A2 (n_5129));
NAND2_X1 i_5181 (.ZN (n_5117), .A1 (n_5118), .A2 (n_5119));
NAND2_X1 i_5180 (.ZN (n_5116), .A1 (n_5117), .A2 (n_5120));
INV_X1 i_5179 (.ZN (n_5115), .A (n_5557));
OAI21_X1 i_5178 (.ZN (n_5114), .A (n_5560), .B1 (n_5115), .B2 (n_5510));
INV_X1 i_5177 (.ZN (n_5113), .A (n_5114));
NAND2_X2 i_5176 (.ZN (n_5112), .A1 (n_5116), .A2 (n_5113));
NAND4_X2 i_5175 (.ZN (n_5111), .A1 (n_5112), .A2 (n_5505), .A3 (n_5139), .A4 (n_5121));
AOI21_X1 i_5171 (.ZN (n_5107), .A (n_6460), .B1 (n_6459), .B2 (n_6493));
INV_X1 i_5170 (.ZN (n_5106), .A (n_5107));
NAND3_X1 i_5169 (.ZN (n_5105), .A1 (n_6493), .A2 (n_6459), .A3 (n_6460));
NAND2_X1 i_5168 (.ZN (n_5104), .A1 (n_5106), .A2 (n_5105));
INV_X1 i_5167 (.ZN (n_5103), .A (n_5104));
INV_X1 i_5166 (.ZN (n_5102), .A (n_6406));
NAND3_X1 i_5165 (.ZN (n_5101), .A1 (n_6419), .A2 (n_6417), .A3 (n_5102));
NAND2_X1 i_5164 (.ZN (n_5100), .A1 (n_6419), .A2 (n_6417));
NAND2_X1 i_5163 (.ZN (n_5099), .A1 (n_5100), .A2 (n_6406));
NAND2_X1 i_5162 (.ZN (n_5098), .A1 (n_5099), .A2 (n_5101));
NAND2_X1 i_5161 (.ZN (n_5097), .A1 (n_6462), .A2 (n_6486));
NAND2_X1 i_5160 (.ZN (n_5096), .A1 (n_5097), .A2 (n_6465));
NAND3_X1 i_5159 (.ZN (n_5095), .A1 (n_6486), .A2 (n_6462), .A3 (n_6466));
NAND2_X1 i_5158 (.ZN (n_5094), .A1 (n_5096), .A2 (n_5095));
NAND2_X1 i_5157 (.ZN (n_5093), .A1 (n_5098), .A2 (n_5094));
NAND4_X1 i_5156 (.ZN (n_5092), .A1 (n_5099), .A2 (n_5095), .A3 (n_5101), .A4 (n_5096));
NAND2_X1 i_5155 (.ZN (n_5091), .A1 (A_imm[26]), .A2 (B_imm[1]));
OAI21_X1 i_5154 (.ZN (n_5090), .A (n_5091), .B1 (n_8423), .B2 (n_8645));
NAND2_X1 i_5153 (.ZN (n_5089), .A1 (B_imm[9]), .A2 (A_imm[18]));
NAND4_X1 i_5152 (.ZN (n_5088), .A1 (B_imm[18]), .A2 (A_imm[26]), .A3 (B_imm[1]), .A4 (A_imm[9]));
NAND2_X1 i_5151 (.ZN (n_5087), .A1 (n_5088), .A2 (n_5089));
AOI22_X1 i_5150 (.ZN (n_5086), .A1 (n_5087), .A2 (n_5090), .B1 (A_imm[28]), .B2 (B_imm[0]));
INV_X1 i_5149 (.ZN (n_5085), .A (n_5086));
NAND2_X1 i_5148 (.ZN (n_5084), .A1 (B_imm[21]), .A2 (A_imm[6]));
OAI21_X1 i_5147 (.ZN (n_5083), .A (n_5084), .B1 (n_8958), .B2 (n_8293));
NAND2_X1 i_5146 (.ZN (n_5082), .A1 (B_imm[15]), .A2 (A_imm[12]));
INV_X1 i_5145 (.ZN (n_5081), .A (n_5082));
NAND4_X1 i_5144 (.ZN (n_5080), .A1 (B_imm[22]), .A2 (B_imm[21]), .A3 (A_imm[6]), .A4 (A_imm[5]));
INV_X1 i_5143 (.ZN (n_5079), .A (n_5080));
OAI21_X1 i_5142 (.ZN (n_5078), .A (n_5083), .B1 (n_5079), .B2 (n_5081));
NAND4_X1 i_5141 (.ZN (n_5077), .A1 (n_5087), .A2 (B_imm[0]), .A3 (A_imm[28]), .A4 (n_5090));
NAND2_X1 i_5140 (.ZN (n_5076), .A1 (n_5077), .A2 (n_5078));
NAND2_X1 i_5139 (.ZN (n_5075), .A1 (n_6475), .A2 (n_6472));
NAND2_X1 i_5138 (.ZN (n_5074), .A1 (n_5075), .A2 (n_6473));
NAND3_X1 i_5137 (.ZN (n_5073), .A1 (n_6475), .A2 (n_6474), .A3 (n_6472));
NAND2_X1 i_5136 (.ZN (n_5072), .A1 (n_5074), .A2 (n_5073));
NAND3_X1 i_5135 (.ZN (n_5071), .A1 (n_5072), .A2 (n_5076), .A3 (n_5085));
AOI21_X1 i_5134 (.ZN (n_5070), .A (n_5086), .B1 (n_5078), .B2 (n_5077));
AOI21_X1 i_5133 (.ZN (n_5069), .A (n_6413), .B1 (n_6414), .B2 (n_6412));
INV_X1 i_5132 (.ZN (n_5068), .A (n_5069));
NAND3_X1 i_5131 (.ZN (n_5067), .A1 (n_6414), .A2 (n_6413), .A3 (n_6412));
NAND2_X1 i_5130 (.ZN (n_5066), .A1 (n_5068), .A2 (n_5067));
OAI21_X1 i_5129 (.ZN (n_5065), .A (n_5066), .B1 (n_5070), .B2 (n_5072));
NAND2_X1 i_5128 (.ZN (n_5064), .A1 (n_5065), .A2 (n_5071));
INV_X1 i_5127 (.ZN (n_5063), .A (n_6410));
OAI21_X1 i_5126 (.ZN (n_5062), .A (n_6407), .B1 (n_5063), .B2 (n_6409));
INV_X1 i_5125 (.ZN (n_5061), .A (n_6409));
INV_X1 i_5124 (.ZN (n_5060), .A (n_6407));
NAND3_X1 i_5123 (.ZN (n_5059), .A1 (n_5061), .A2 (n_6410), .A3 (n_5060));
NAND3_X1 i_5122 (.ZN (n_5058), .A1 (n_5064), .A2 (n_5062), .A3 (n_5059));
NAND2_X1 i_5121 (.ZN (n_5057), .A1 (n_5062), .A2 (n_5059));
NAND3_X1 i_5120 (.ZN (n_5056), .A1 (n_5057), .A2 (n_5065), .A3 (n_5071));
NAND2_X1 i_5119 (.ZN (n_5055), .A1 (n_6441), .A2 (n_6439));
NAND3_X1 i_5118 (.ZN (n_5054), .A1 (n_5055), .A2 (B_imm[1]), .A3 (A_imm[29]));
NAND3_X1 i_5117 (.ZN (n_5053), .A1 (n_6441), .A2 (n_6440), .A3 (n_6439));
NAND2_X1 i_5116 (.ZN (n_5052), .A1 (n_5054), .A2 (n_5053));
NAND2_X1 i_5115 (.ZN (n_5051), .A1 (n_5056), .A2 (n_5052));
NAND2_X1 i_5114 (.ZN (n_5050), .A1 (n_5058), .A2 (n_5051));
NAND2_X1 i_5113 (.ZN (n_5049), .A1 (n_5050), .A2 (n_5092));
NAND2_X1 i_5112 (.ZN (n_5048), .A1 (n_5049), .A2 (n_5093));
NAND2_X1 i_5111 (.ZN (n_5047), .A1 (n_5048), .A2 (n_5103));
NAND3_X2 i_5110 (.ZN (n_5046), .A1 (n_5104), .A2 (n_5093), .A3 (n_5049));
OAI211_X1 i_5109 (.ZN (n_5045), .A (n_6403), .B (n_6402), .C1 (n_6401), .C2 (n_6399));
NAND2_X1 i_5108 (.ZN (n_5044), .A1 (n_6403), .A2 (n_6402));
NAND2_X1 i_5107 (.ZN (n_5043), .A1 (n_5044), .A2 (n_6398));
NAND2_X1 i_5106 (.ZN (n_5042), .A1 (n_5043), .A2 (n_5045));
NAND2_X1 i_5105 (.ZN (n_5041), .A1 (n_5042), .A2 (n_5046));
INV_X1 i_5104 (.ZN (n_5040), .A (n_6548));
NAND3_X1 i_5103 (.ZN (n_5039), .A1 (n_6552), .A2 (n_6551), .A3 (n_5040));
NAND2_X1 i_5102 (.ZN (n_5038), .A1 (n_6551), .A2 (n_6552));
NAND2_X1 i_5101 (.ZN (n_5037), .A1 (n_5038), .A2 (n_6548));
NAND2_X1 i_5100 (.ZN (n_5036), .A1 (n_5037), .A2 (n_5039));
NAND3_X1 i_5099 (.ZN (n_5035), .A1 (n_5041), .A2 (n_5047), .A3 (n_5036));
NAND2_X1 i_5098 (.ZN (n_5034), .A1 (n_5041), .A2 (n_5047));
INV_X1 i_5097 (.ZN (n_5033), .A (n_5036));
NAND2_X1 i_5096 (.ZN (n_5032), .A1 (n_5034), .A2 (n_5033));
AOI21_X1 i_5095 (.ZN (n_5031), .A (n_6392), .B1 (n_6393), .B2 (n_6456));
NAND3_X1 i_5094 (.ZN (n_5030), .A1 (n_6393), .A2 (n_6392), .A3 (n_6456));
INV_X1 i_5093 (.ZN (n_5029), .A (n_5030));
NOR2_X1 i_5092 (.ZN (n_5028), .A1 (n_5029), .A2 (n_5031));
NAND3_X1 i_5091 (.ZN (n_5027), .A1 (n_5032), .A2 (n_5035), .A3 (n_5028));
INV_X1 i_5090 (.ZN (n_5026), .A (n_5027));
AOI21_X1 i_5089 (.ZN (n_5025), .A (n_5028), .B1 (n_5032), .B2 (n_5035));
INV_X1 i_5088 (.ZN (n_5024), .A (n_5751));
NAND2_X1 i_5087 (.ZN (n_5023), .A1 (n_5860), .A2 (n_5859));
NAND2_X1 i_5086 (.ZN (n_5022), .A1 (n_5023), .A2 (n_5024));
NAND3_X1 i_5085 (.ZN (n_5021), .A1 (n_5860), .A2 (n_5859), .A3 (n_5751));
NAND2_X1 i_5084 (.ZN (n_5020), .A1 (n_5022), .A2 (n_5021));
OAI21_X1 i_5083 (.ZN (n_5019), .A (n_5020), .B1 (n_5026), .B2 (n_5025));
NAND2_X1 i_5082 (.ZN (n_5018), .A1 (n_5032), .A2 (n_5035));
INV_X1 i_5081 (.ZN (n_5017), .A (n_5028));
NAND2_X1 i_5080 (.ZN (n_5016), .A1 (n_5018), .A2 (n_5017));
NAND4_X1 i_5079 (.ZN (n_5015), .A1 (n_5016), .A2 (n_5027), .A3 (n_5022), .A4 (n_5021));
NAND2_X1 i_5078 (.ZN (n_5014), .A1 (n_5015), .A2 (n_5019));
NAND3_X1 i_5077 (.ZN (n_5013), .A1 (n_5050), .A2 (n_5093), .A3 (n_5092));
NAND2_X1 i_5076 (.ZN (n_5012), .A1 (n_5093), .A2 (n_5092));
NAND3_X1 i_5075 (.ZN (n_5011), .A1 (n_5012), .A2 (n_5058), .A3 (n_5051));
NAND2_X1 i_5074 (.ZN (n_5010), .A1 (n_5011), .A2 (n_5013));
INV_X1 i_5073 (.ZN (n_5009), .A (n_5010));
INV_X1 i_5072 (.ZN (n_5008), .A (n_6161));
NAND2_X1 i_5071 (.ZN (n_5007), .A1 (n_6170), .A2 (n_6165));
NAND2_X1 i_5070 (.ZN (n_5006), .A1 (n_5007), .A2 (n_5008));
NAND3_X1 i_5069 (.ZN (n_5005), .A1 (n_6170), .A2 (n_6165), .A3 (n_6161));
NAND2_X1 i_5068 (.ZN (n_5004), .A1 (n_5006), .A2 (n_5005));
NAND2_X1 i_5067 (.ZN (n_5003), .A1 (n_6182), .A2 (n_6175));
NAND2_X1 i_5066 (.ZN (n_5002), .A1 (n_5003), .A2 (n_6169));
NAND3_X1 i_5065 (.ZN (n_5001), .A1 (n_6182), .A2 (n_6176), .A3 (n_6175));
NAND2_X1 i_5064 (.ZN (n_5000), .A1 (n_5002), .A2 (n_5001));
NAND2_X1 i_5063 (.ZN (n_4999), .A1 (A_imm[27]), .A2 (B_imm[1]));
NAND2_X1 i_5062 (.ZN (n_4998), .A1 (B_imm[13]), .A2 (A_imm[14]));
NAND2_X1 i_5061 (.ZN (n_4997), .A1 (B_imm[25]), .A2 (A_imm[2]));
NAND2_X1 i_5060 (.ZN (n_4996), .A1 (n_4997), .A2 (n_4998));
NAND2_X1 i_5059 (.ZN (n_4995), .A1 (B_imm[20]), .A2 (A_imm[7]));
NAND4_X1 i_5058 (.ZN (n_4994), .A1 (B_imm[25]), .A2 (B_imm[13]), .A3 (A_imm[14]), .A4 (A_imm[2]));
NAND2_X1 i_5057 (.ZN (n_4993), .A1 (n_4994), .A2 (n_4995));
NAND2_X1 i_5056 (.ZN (n_4992), .A1 (n_4993), .A2 (n_4996));
NAND2_X1 i_5055 (.ZN (n_4991), .A1 (n_4992), .A2 (n_4999));
NAND2_X1 i_5054 (.ZN (n_4990), .A1 (B_imm[24]), .A2 (A_imm[3]));
NAND2_X1 i_5053 (.ZN (n_4989), .A1 (A_imm[19]), .A2 (B_imm[7]));
NAND2_X1 i_5052 (.ZN (n_4988), .A1 (A_imm[9]), .A2 (B_imm[17]));
NAND2_X1 i_5051 (.ZN (n_4987), .A1 (n_4989), .A2 (n_4988));
NAND2_X1 i_5050 (.ZN (n_4986), .A1 (B_imm[16]), .A2 (A_imm[10]));
INV_X1 i_5049 (.ZN (n_4985), .A (n_4986));
NAND4_X1 i_5048 (.ZN (n_4984), .A1 (A_imm[19]), .A2 (B_imm[17]), .A3 (A_imm[9]), .A4 (B_imm[7]));
INV_X1 i_5047 (.ZN (n_4983), .A (n_4984));
OAI21_X1 i_5046 (.ZN (n_4982), .A (n_4987), .B1 (n_4983), .B2 (n_4985));
NAND2_X1 i_5045 (.ZN (n_4981), .A1 (n_4982), .A2 (n_4990));
NAND2_X1 i_5044 (.ZN (n_4980), .A1 (B_imm[23]), .A2 (A_imm[4]));
INV_X1 i_5043 (.ZN (n_4979), .A (n_4980));
NAND2_X1 i_5042 (.ZN (n_4978), .A1 (n_4984), .A2 (n_4986));
NAND4_X1 i_5041 (.ZN (n_4977), .A1 (n_4978), .A2 (B_imm[24]), .A3 (A_imm[3]), .A4 (n_4987));
INV_X1 i_5040 (.ZN (n_4976), .A (n_4977));
OAI21_X1 i_5039 (.ZN (n_4975), .A (n_4981), .B1 (n_4976), .B2 (n_4979));
NAND4_X1 i_5038 (.ZN (n_4974), .A1 (n_4993), .A2 (B_imm[1]), .A3 (A_imm[27]), .A4 (n_4996));
NAND2_X1 i_5037 (.ZN (n_4973), .A1 (n_4974), .A2 (n_4975));
NAND3_X1 i_5036 (.ZN (n_4972), .A1 (n_5000), .A2 (n_4973), .A3 (n_4991));
INV_X1 i_5035 (.ZN (n_4971), .A (n_5000));
INV_X1 i_5034 (.ZN (n_4970), .A (n_4975));
INV_X1 i_5033 (.ZN (n_4969), .A (n_4974));
OAI21_X1 i_5032 (.ZN (n_4968), .A (n_4991), .B1 (n_4969), .B2 (n_4970));
AOI21_X1 i_5031 (.ZN (n_4967), .A (n_6445), .B1 (n_6444), .B2 (n_6446));
NAND3_X1 i_5030 (.ZN (n_4966), .A1 (n_6446), .A2 (n_6445), .A3 (n_6444));
INV_X1 i_5029 (.ZN (n_4965), .A (n_4966));
NOR2_X1 i_5028 (.ZN (n_4964), .A1 (n_4965), .A2 (n_4967));
AOI21_X1 i_5027 (.ZN (n_4963), .A (n_4964), .B1 (n_4968), .B2 (n_4971));
INV_X1 i_5026 (.ZN (n_4962), .A (n_4963));
NAND3_X1 i_5025 (.ZN (n_4961), .A1 (n_4962), .A2 (n_5004), .A3 (n_4972));
INV_X1 i_5024 (.ZN (n_4960), .A (n_4972));
OAI211_X1 i_5023 (.ZN (n_4959), .A (n_5006), .B (n_5005), .C1 (n_4963), .C2 (n_4960));
NAND3_X1 i_5022 (.ZN (n_4958), .A1 (n_5963), .A2 (n_5970), .A3 (n_5966));
NAND2_X1 i_5021 (.ZN (n_4957), .A1 (n_5963), .A2 (n_5970));
NAND2_X1 i_5020 (.ZN (n_4956), .A1 (n_4957), .A2 (n_5965));
NAND2_X1 i_5019 (.ZN (n_4955), .A1 (n_4956), .A2 (n_4958));
NAND3_X1 i_5018 (.ZN (n_4954), .A1 (n_4959), .A2 (n_4961), .A3 (n_4955));
INV_X1 i_5017 (.ZN (n_4953), .A (n_4954));
AOI21_X1 i_5016 (.ZN (n_4952), .A (n_4955), .B1 (n_4959), .B2 (n_4961));
NOR2_X1 i_5015 (.ZN (n_4951), .A1 (n_4953), .A2 (n_4952));
NAND2_X1 i_5014 (.ZN (n_4950), .A1 (n_4968), .A2 (n_4971));
INV_X1 i_5013 (.ZN (n_4949), .A (n_4964));
AOI21_X1 i_5012 (.ZN (n_4948), .A (n_4949), .B1 (n_4950), .B2 (n_4972));
INV_X1 i_5011 (.ZN (n_4947), .A (n_4948));
NAND3_X1 i_5010 (.ZN (n_4946), .A1 (n_4950), .A2 (n_4972), .A3 (n_4949));
NAND2_X1 i_5009 (.ZN (n_4945), .A1 (n_5076), .A2 (n_5085));
INV_X1 i_5008 (.ZN (n_4944), .A (n_5072));
NAND2_X1 i_5007 (.ZN (n_4943), .A1 (n_4945), .A2 (n_4944));
AOI21_X1 i_5006 (.ZN (n_4942), .A (n_5066), .B1 (n_4943), .B2 (n_5071));
INV_X1 i_5005 (.ZN (n_4941), .A (n_4942));
NAND3_X1 i_5004 (.ZN (n_4940), .A1 (n_4943), .A2 (n_5071), .A3 (n_5066));
NAND4_X2 i_5003 (.ZN (n_4939), .A1 (n_4947), .A2 (n_4941), .A3 (n_4946), .A4 (n_4940));
INV_X1 i_5002 (.ZN (n_4938), .A (n_4946));
NOR2_X1 i_5001 (.ZN (n_4937), .A1 (n_4948), .A2 (n_4938));
INV_X1 i_5000 (.ZN (n_4936), .A (n_4940));
NOR2_X1 i_4999 (.ZN (n_4935), .A1 (n_4936), .A2 (n_4942));
NAND2_X1 i_4998 (.ZN (n_4934), .A1 (n_4991), .A2 (n_4974));
NAND2_X1 i_4997 (.ZN (n_4933), .A1 (n_4934), .A2 (n_4970));
NAND3_X1 i_4996 (.ZN (n_4932), .A1 (n_4991), .A2 (n_4974), .A3 (n_4975));
NAND2_X1 i_4995 (.ZN (n_4931), .A1 (n_4933), .A2 (n_4932));
NAND2_X1 i_4994 (.ZN (n_4930), .A1 (n_5083), .A2 (n_5080));
NAND2_X1 i_4993 (.ZN (n_4929), .A1 (n_4930), .A2 (n_5081));
NAND3_X1 i_4992 (.ZN (n_4928), .A1 (n_5083), .A2 (n_5080), .A3 (n_5082));
NAND2_X1 i_4991 (.ZN (n_4927), .A1 (n_4929), .A2 (n_4928));
INV_X1 i_4990 (.ZN (n_4926), .A (n_5089));
NAND2_X1 i_4989 (.ZN (n_4925), .A1 (n_5090), .A2 (n_5088));
NAND2_X1 i_4988 (.ZN (n_4924), .A1 (n_4925), .A2 (n_4926));
NAND3_X1 i_4987 (.ZN (n_4923), .A1 (n_5090), .A2 (n_5088), .A3 (n_5089));
NAND2_X1 i_4986 (.ZN (n_4922), .A1 (n_4924), .A2 (n_4923));
NAND2_X1 i_4985 (.ZN (n_4921), .A1 (n_4927), .A2 (n_4922));
OAI22_X1 i_4984 (.ZN (n_4920), .A1 (n_8971), .A2 (n_8880), .B1 (n_8909), .B2 (n_8644));
NAND2_X1 i_4983 (.ZN (n_4919), .A1 (A_imm[19]), .A2 (B_imm[5]));
NAND4_X1 i_4982 (.ZN (n_4918), .A1 (A_imm[14]), .A2 (B_imm[10]), .A3 (B_imm[17]), .A4 (A_imm[7]));
NAND2_X1 i_4981 (.ZN (n_4917), .A1 (n_4919), .A2 (n_4918));
NAND2_X1 i_4980 (.ZN (n_4916), .A1 (n_4917), .A2 (n_4920));
OAI21_X1 i_4979 (.ZN (n_4915), .A (n_4916), .B1 (n_8347), .B2 (n_8858));
NAND2_X1 i_4978 (.ZN (n_4914), .A1 (B_imm[24]), .A2 (A_imm[1]));
NAND4_X1 i_4977 (.ZN (n_4913), .A1 (n_4917), .A2 (B_imm[9]), .A3 (A_imm[16]), .A4 (n_4920));
NAND2_X1 i_4976 (.ZN (n_4912), .A1 (n_4913), .A2 (n_4914));
NAND2_X1 i_4975 (.ZN (n_4911), .A1 (n_4912), .A2 (n_4915));
NAND2_X1 i_4974 (.ZN (n_4910), .A1 (B_imm[11]), .A2 (A_imm[14]));
OAI21_X1 i_4973 (.ZN (n_4909), .A (n_4910), .B1 (n_8794), .B2 (n_6740));
NAND2_X1 i_4972 (.ZN (n_4908), .A1 (B_imm[18]), .A2 (A_imm[7]));
NAND4_X1 i_4971 (.ZN (n_4907), .A1 (A_imm[25]), .A2 (B_imm[11]), .A3 (B_imm[0]), .A4 (A_imm[14]));
NAND2_X1 i_4970 (.ZN (n_4906), .A1 (n_4907), .A2 (n_4908));
NAND2_X1 i_4969 (.ZN (n_4905), .A1 (n_4906), .A2 (n_4909));
NAND2_X1 i_4968 (.ZN (n_4904), .A1 (n_4911), .A2 (n_4905));
NAND2_X1 i_4967 (.ZN (n_4903), .A1 (B_imm[15]), .A2 (A_imm[10]));
NAND2_X1 i_4966 (.ZN (n_4902), .A1 (B_imm[22]), .A2 (A_imm[3]));
NAND2_X1 i_4965 (.ZN (n_4901), .A1 (n_4903), .A2 (n_4902));
NAND2_X1 i_4964 (.ZN (n_4900), .A1 (B_imm[25]), .A2 (A_imm[0]));
INV_X1 i_4963 (.ZN (n_4899), .A (n_4900));
NAND4_X1 i_4962 (.ZN (n_4898), .A1 (B_imm[15]), .A2 (B_imm[22]), .A3 (A_imm[10]), .A4 (A_imm[3]));
INV_X1 i_4961 (.ZN (n_4897), .A (n_4898));
OAI21_X1 i_4960 (.ZN (n_4896), .A (n_4901), .B1 (n_4897), .B2 (n_4899));
NAND4_X1 i_4959 (.ZN (n_4895), .A1 (n_4912), .A2 (n_4906), .A3 (n_4915), .A4 (n_4909));
NAND2_X1 i_4958 (.ZN (n_4894), .A1 (n_4895), .A2 (n_4896));
NAND4_X1 i_4957 (.ZN (n_4893), .A1 (n_4929), .A2 (n_4928), .A3 (n_4924), .A4 (n_4923));
NAND3_X1 i_4956 (.ZN (n_4892), .A1 (n_4893), .A2 (n_4904), .A3 (n_4894));
NAND2_X1 i_4955 (.ZN (n_4891), .A1 (n_4892), .A2 (n_4921));
NAND2_X1 i_4954 (.ZN (n_4890), .A1 (n_4891), .A2 (n_4931));
NAND4_X1 i_4953 (.ZN (n_4889), .A1 (n_4892), .A2 (n_4933), .A3 (n_4932), .A4 (n_4921));
INV_X1 i_4952 (.ZN (n_4888), .A (n_4889));
NAND2_X1 i_4951 (.ZN (n_4887), .A1 (B_imm[14]), .A2 (A_imm[14]));
INV_X1 i_4950 (.ZN (n_4886), .A (n_6450));
NAND2_X1 i_4949 (.ZN (n_4885), .A1 (n_6451), .A2 (n_6449));
NAND2_X1 i_4948 (.ZN (n_4884), .A1 (n_4885), .A2 (n_4886));
NAND3_X1 i_4947 (.ZN (n_4883), .A1 (n_6451), .A2 (n_6450), .A3 (n_6449));
NAND2_X1 i_4946 (.ZN (n_4882), .A1 (n_4884), .A2 (n_4883));
INV_X1 i_4945 (.ZN (n_4881), .A (n_4882));
NAND2_X1 i_4944 (.ZN (n_4880), .A1 (n_4887), .A2 (n_4881));
NAND3_X1 i_4943 (.ZN (n_4879), .A1 (n_4882), .A2 (B_imm[14]), .A3 (A_imm[14]));
NAND2_X1 i_4942 (.ZN (n_4878), .A1 (n_4880), .A2 (n_4879));
NAND2_X1 i_4941 (.ZN (n_4877), .A1 (n_6180), .A2 (n_6178));
NAND3_X1 i_4940 (.ZN (n_4876), .A1 (n_4877), .A2 (B_imm[8]), .A3 (A_imm[20]));
NAND3_X1 i_4939 (.ZN (n_4875), .A1 (n_6180), .A2 (n_6179), .A3 (n_6178));
NAND3_X1 i_4938 (.ZN (n_4874), .A1 (n_4878), .A2 (n_4876), .A3 (n_4875));
NAND2_X1 i_4937 (.ZN (n_4873), .A1 (n_4876), .A2 (n_4875));
NAND3_X1 i_4936 (.ZN (n_4872), .A1 (n_4880), .A2 (n_4879), .A3 (n_4873));
NAND2_X1 i_4935 (.ZN (n_4871), .A1 (n_4874), .A2 (n_4872));
OAI21_X1 i_4934 (.ZN (n_4870), .A (n_4890), .B1 (n_4888), .B2 (n_4871));
OAI21_X1 i_4933 (.ZN (n_4869), .A (n_4870), .B1 (n_4937), .B2 (n_4935));
NAND2_X1 i_4932 (.ZN (n_4868), .A1 (n_4869), .A2 (n_4939));
NAND2_X1 i_4931 (.ZN (n_4867), .A1 (n_4951), .A2 (n_4868));
OAI211_X2 i_4930 (.ZN (n_4866), .A (n_4869), .B (n_4939), .C1 (n_4953), .C2 (n_4952));
INV_X1 i_4929 (.ZN (n_4865), .A (n_5895));
NAND2_X1 i_4928 (.ZN (n_4864), .A1 (n_5887), .A2 (n_5895));
INV_X1 i_4927 (.ZN (n_4863), .A (n_4864));
OAI22_X1 i_4926 (.ZN (n_4862), .A1 (n_4863), .A2 (n_5888), .B1 (n_5886), .B2 (n_4865));
INV_X1 i_4925 (.ZN (n_4861), .A (n_4862));
INV_X1 i_4924 (.ZN (n_4860), .A (n_5978));
INV_X1 i_4923 (.ZN (n_4859), .A (n_5977));
OAI21_X1 i_4922 (.ZN (n_4858), .A (n_4860), .B1 (n_4859), .B2 (n_5980));
NAND3_X1 i_4921 (.ZN (n_4857), .A1 (n_5979), .A2 (n_5978), .A3 (n_5977));
NAND2_X1 i_4920 (.ZN (n_4856), .A1 (n_4880), .A2 (n_4873));
NAND4_X1 i_4919 (.ZN (n_4855), .A1 (n_4856), .A2 (n_4857), .A3 (n_4858), .A4 (n_4879));
NAND2_X1 i_4918 (.ZN (n_4854), .A1 (n_4857), .A2 (n_4858));
NAND2_X1 i_4917 (.ZN (n_4853), .A1 (n_4856), .A2 (n_4879));
NAND2_X1 i_4916 (.ZN (n_4852), .A1 (n_4853), .A2 (n_4854));
NAND3_X1 i_4915 (.ZN (n_4851), .A1 (n_4861), .A2 (n_4855), .A3 (n_4852));
NAND2_X1 i_4914 (.ZN (n_4850), .A1 (n_4855), .A2 (n_4852));
NAND2_X1 i_4913 (.ZN (n_4849), .A1 (n_4850), .A2 (n_4862));
NAND2_X1 i_4912 (.ZN (n_4848), .A1 (n_4849), .A2 (n_4851));
NAND2_X1 i_4911 (.ZN (n_4847), .A1 (n_4981), .A2 (n_4977));
NAND2_X1 i_4910 (.ZN (n_4846), .A1 (n_4847), .A2 (n_4979));
NAND3_X1 i_4909 (.ZN (n_4845), .A1 (n_4981), .A2 (n_4980), .A3 (n_4977));
NAND2_X1 i_4908 (.ZN (n_4844), .A1 (n_4846), .A2 (n_4845));
INV_X1 i_4907 (.ZN (n_4843), .A (n_4995));
NAND2_X1 i_4906 (.ZN (n_4842), .A1 (n_4996), .A2 (n_4994));
NAND2_X1 i_4905 (.ZN (n_4841), .A1 (n_4842), .A2 (n_4843));
NAND3_X1 i_4904 (.ZN (n_4840), .A1 (n_4996), .A2 (n_4994), .A3 (n_4995));
NAND2_X1 i_4903 (.ZN (n_4839), .A1 (n_4841), .A2 (n_4840));
NAND2_X1 i_4902 (.ZN (n_4838), .A1 (n_4844), .A2 (n_4839));
NAND4_X1 i_4901 (.ZN (n_4837), .A1 (n_4841), .A2 (n_4846), .A3 (n_4845), .A4 (n_4840));
NAND2_X1 i_4900 (.ZN (n_4836), .A1 (B_imm[19]), .A2 (A_imm[8]));
INV_X1 i_4899 (.ZN (n_4835), .A (n_4836));
NAND2_X1 i_4898 (.ZN (n_4834), .A1 (B_imm[26]), .A2 (A_imm[1]));
NAND2_X1 i_4897 (.ZN (n_4833), .A1 (A_imm[22]), .A2 (B_imm[4]));
OAI21_X1 i_4896 (.ZN (n_4832), .A (n_4833), .B1 (n_8859), .B2 (n_8429));
NAND2_X1 i_4895 (.ZN (n_4831), .A1 (A_imm[16]), .A2 (B_imm[10]));
NAND4_X1 i_4894 (.ZN (n_4830), .A1 (A_imm[21]), .A2 (A_imm[22]), .A3 (B_imm[5]), .A4 (B_imm[4]));
NAND2_X1 i_4893 (.ZN (n_4829), .A1 (n_4830), .A2 (n_4831));
NAND2_X1 i_4892 (.ZN (n_4828), .A1 (n_4829), .A2 (n_4832));
NAND2_X1 i_4891 (.ZN (n_4827), .A1 (n_4828), .A2 (n_4834));
NAND4_X1 i_4890 (.ZN (n_4826), .A1 (n_4829), .A2 (B_imm[26]), .A3 (A_imm[1]), .A4 (n_4832));
NAND2_X1 i_4889 (.ZN (n_4825), .A1 (n_4827), .A2 (n_4826));
NAND2_X1 i_4888 (.ZN (n_4824), .A1 (n_4825), .A2 (n_4835));
NAND3_X1 i_4887 (.ZN (n_4823), .A1 (n_4827), .A2 (n_4836), .A3 (n_4826));
NAND2_X1 i_4886 (.ZN (n_4822), .A1 (n_4824), .A2 (n_4823));
NAND2_X1 i_4885 (.ZN (n_4821), .A1 (n_4837), .A2 (n_4822));
NAND2_X1 i_4884 (.ZN (n_4820), .A1 (n_4821), .A2 (n_4838));
OAI22_X1 i_4883 (.ZN (n_4819), .A1 (n_8795), .A2 (n_8971), .B1 (n_8767), .B2 (n_6584));
NAND2_X1 i_4882 (.ZN (n_4818), .A1 (B_imm[11]), .A2 (A_imm[15]));
INV_X1 i_4881 (.ZN (n_4817), .A (n_4818));
NAND4_X1 i_4880 (.ZN (n_4816), .A1 (B_imm[12]), .A2 (A_imm[24]), .A3 (B_imm[2]), .A4 (A_imm[14]));
INV_X1 i_4879 (.ZN (n_4815), .A (n_4816));
OAI21_X1 i_4878 (.ZN (n_4814), .A (n_4819), .B1 (n_4815), .B2 (n_4817));
INV_X1 i_4877 (.ZN (n_4813), .A (n_4814));
OAI22_X1 i_4876 (.ZN (n_4812), .A1 (n_8947), .A2 (n_8956), .B1 (n_8893), .B2 (n_8232));
NAND2_X1 i_4875 (.ZN (n_4811), .A1 (A_imm[23]), .A2 (B_imm[3]));
NAND4_X1 i_4874 (.ZN (n_4810), .A1 (B_imm[8]), .A2 (A_imm[20]), .A3 (B_imm[6]), .A4 (A_imm[18]));
NAND2_X1 i_4873 (.ZN (n_4809), .A1 (n_4810), .A2 (n_4811));
AOI22_X1 i_4872 (.ZN (n_4808), .A1 (n_4809), .A2 (n_4812), .B1 (B_imm[27]), .B2 (A_imm[0]));
NAND2_X1 i_4871 (.ZN (n_4807), .A1 (B_imm[27]), .A2 (A_imm[0]));
INV_X1 i_4870 (.ZN (n_4806), .A (n_4807));
NAND3_X1 i_4869 (.ZN (n_4805), .A1 (n_4806), .A2 (n_4812), .A3 (n_4809));
INV_X1 i_4868 (.ZN (n_4804), .A (n_4805));
OAI21_X1 i_4867 (.ZN (n_4803), .A (n_4813), .B1 (n_4804), .B2 (n_4808));
INV_X1 i_4866 (.ZN (n_4802), .A (n_4808));
NAND3_X1 i_4865 (.ZN (n_4801), .A1 (n_4802), .A2 (n_4814), .A3 (n_4805));
NAND2_X1 i_4864 (.ZN (n_4800), .A1 (n_4803), .A2 (n_4801));
NAND2_X1 i_4863 (.ZN (n_4799), .A1 (B_imm[23]), .A2 (A_imm[2]));
NAND2_X1 i_4862 (.ZN (n_4798), .A1 (A_imm[17]), .A2 (B_imm[7]));
OAI21_X1 i_4861 (.ZN (n_4797), .A (n_4798), .B1 (n_8908), .B2 (n_8511));
NAND2_X1 i_4860 (.ZN (n_4796), .A1 (A_imm[22]), .A2 (B_imm[2]));
NAND4_X1 i_4859 (.ZN (n_4795), .A1 (B_imm[16]), .A2 (A_imm[17]), .A3 (B_imm[7]), .A4 (A_imm[8]));
NAND2_X1 i_4858 (.ZN (n_4794), .A1 (n_4795), .A2 (n_4796));
NAND2_X1 i_4857 (.ZN (n_4793), .A1 (n_4794), .A2 (n_4797));
NAND2_X1 i_4856 (.ZN (n_4792), .A1 (n_4793), .A2 (n_4799));
NAND2_X1 i_4855 (.ZN (n_4791), .A1 (B_imm[21]), .A2 (A_imm[4]));
OAI21_X1 i_4854 (.ZN (n_4790), .A (n_4791), .B1 (n_4793), .B2 (n_4799));
NAND2_X1 i_4853 (.ZN (n_4789), .A1 (n_4987), .A2 (n_4984));
NAND2_X1 i_4852 (.ZN (n_4788), .A1 (n_4789), .A2 (n_4985));
NAND3_X1 i_4851 (.ZN (n_4787), .A1 (n_4987), .A2 (n_4986), .A3 (n_4984));
NAND2_X1 i_4850 (.ZN (n_4786), .A1 (n_4788), .A2 (n_4787));
NAND3_X1 i_4849 (.ZN (n_4785), .A1 (n_4790), .A2 (n_4792), .A3 (n_4786));
AOI21_X1 i_4848 (.ZN (n_4784), .A (n_4786), .B1 (n_4792), .B2 (n_4790));
NAND2_X1 i_4847 (.ZN (n_4783), .A1 (n_4832), .A2 (n_4830));
XNOR2_X1 i_4846 (.ZN (n_4782), .A (n_4783), .B (n_4831));
OAI21_X1 i_4845 (.ZN (n_4781), .A (n_4785), .B1 (n_4784), .B2 (n_4782));
NAND2_X1 i_4844 (.ZN (n_4780), .A1 (n_4781), .A2 (n_4800));
OAI22_X1 i_4843 (.ZN (n_4779), .A1 (n_8860), .A2 (n_8293), .B1 (n_8973), .B2 (n_8752));
OAI22_X1 i_4842 (.ZN (n_4778), .A1 (n_8232), .A2 (n_8956), .B1 (n_8859), .B2 (n_6817));
NAND2_X1 i_4841 (.ZN (n_4777), .A1 (A_imm[20]), .A2 (B_imm[4]));
INV_X1 i_4840 (.ZN (n_4776), .A (n_4777));
NAND4_X1 i_4839 (.ZN (n_4775), .A1 (B_imm[6]), .A2 (A_imm[18]), .A3 (A_imm[21]), .A4 (B_imm[3]));
INV_X1 i_4838 (.ZN (n_4774), .A (n_4775));
OAI21_X1 i_4837 (.ZN (n_4773), .A (n_4778), .B1 (n_4774), .B2 (n_4776));
NAND4_X1 i_4836 (.ZN (n_4772), .A1 (B_imm[20]), .A2 (B_imm[13]), .A3 (A_imm[12]), .A4 (A_imm[5]));
NAND2_X1 i_4835 (.ZN (n_4771), .A1 (n_4773), .A2 (n_4772));
NAND4_X1 i_4834 (.ZN (n_4770), .A1 (n_4771), .A2 (n_4779), .A3 (B_imm[14]), .A4 (A_imm[12]));
NAND2_X1 i_4833 (.ZN (n_4769), .A1 (B_imm[14]), .A2 (A_imm[12]));
NAND2_X1 i_4832 (.ZN (n_4768), .A1 (n_4771), .A2 (n_4779));
NAND2_X1 i_4831 (.ZN (n_4767), .A1 (n_4768), .A2 (n_4769));
NAND2_X1 i_4830 (.ZN (n_4766), .A1 (n_4812), .A2 (n_4810));
NAND3_X1 i_4829 (.ZN (n_4765), .A1 (n_4766), .A2 (B_imm[3]), .A3 (A_imm[23]));
NAND3_X1 i_4828 (.ZN (n_4764), .A1 (n_4812), .A2 (n_4811), .A3 (n_4810));
NAND2_X1 i_4827 (.ZN (n_4763), .A1 (n_4765), .A2 (n_4764));
NAND2_X1 i_4826 (.ZN (n_4762), .A1 (n_4767), .A2 (n_4763));
NAND2_X1 i_4825 (.ZN (n_4761), .A1 (n_4762), .A2 (n_4770));
OAI21_X1 i_4824 (.ZN (n_4760), .A (n_4761), .B1 (n_4800), .B2 (n_4781));
NAND2_X1 i_4823 (.ZN (n_4759), .A1 (n_4760), .A2 (n_4780));
NAND2_X1 i_4822 (.ZN (n_4758), .A1 (n_4759), .A2 (n_4820));
INV_X1 i_4821 (.ZN (n_4757), .A (n_4820));
NAND3_X1 i_4820 (.ZN (n_4756), .A1 (n_4760), .A2 (n_4757), .A3 (n_4780));
INV_X1 i_4819 (.ZN (n_4755), .A (n_4826));
OAI21_X1 i_4818 (.ZN (n_4754), .A (n_4827), .B1 (n_4755), .B2 (n_4835));
AOI21_X1 i_4817 (.ZN (n_4753), .A (n_5983), .B1 (n_5984), .B2 (n_5982));
NAND3_X1 i_4816 (.ZN (n_4752), .A1 (n_5984), .A2 (n_5983), .A3 (n_5982));
INV_X1 i_4815 (.ZN (n_4751), .A (n_4752));
NOR2_X1 i_4814 (.ZN (n_4750), .A1 (n_4751), .A2 (n_4753));
NAND2_X1 i_4813 (.ZN (n_4749), .A1 (n_4750), .A2 (n_4754));
NAND2_X1 i_4812 (.ZN (n_4748), .A1 (n_4826), .A2 (n_4836));
INV_X1 i_4811 (.ZN (n_4747), .A (n_5983));
NAND2_X1 i_4810 (.ZN (n_4746), .A1 (n_5984), .A2 (n_5982));
NAND2_X1 i_4809 (.ZN (n_4745), .A1 (n_4746), .A2 (n_4747));
NAND2_X1 i_4808 (.ZN (n_4744), .A1 (n_4745), .A2 (n_4752));
NAND3_X1 i_4807 (.ZN (n_4743), .A1 (n_4744), .A2 (n_4827), .A3 (n_4748));
NAND2_X1 i_4806 (.ZN (n_4742), .A1 (n_4743), .A2 (n_4749));
INV_X1 i_4805 (.ZN (n_4741), .A (n_5899));
NAND2_X1 i_4804 (.ZN (n_4740), .A1 (n_5900), .A2 (n_5898));
NAND2_X1 i_4803 (.ZN (n_4739), .A1 (n_4740), .A2 (n_4741));
NAND3_X1 i_4802 (.ZN (n_4738), .A1 (n_5900), .A2 (n_5899), .A3 (n_5898));
NAND3_X1 i_4801 (.ZN (n_4737), .A1 (n_4742), .A2 (n_4739), .A3 (n_4738));
NAND2_X1 i_4800 (.ZN (n_4736), .A1 (n_4739), .A2 (n_4738));
NAND3_X1 i_4799 (.ZN (n_4735), .A1 (n_4743), .A2 (n_4749), .A3 (n_4736));
NAND2_X1 i_4798 (.ZN (n_4734), .A1 (n_4737), .A2 (n_4735));
INV_X1 i_4797 (.ZN (n_4733), .A (n_4734));
NAND2_X1 i_4796 (.ZN (n_4732), .A1 (n_4756), .A2 (n_4733));
NAND2_X1 i_4795 (.ZN (n_4731), .A1 (n_4732), .A2 (n_4758));
NAND2_X1 i_4794 (.ZN (n_4730), .A1 (n_4731), .A2 (n_4848));
INV_X1 i_4793 (.ZN (n_4729), .A (n_4848));
NAND3_X1 i_4792 (.ZN (n_4728), .A1 (n_4729), .A2 (n_4732), .A3 (n_4758));
INV_X1 i_4791 (.ZN (n_4727), .A (n_5940));
NAND3_X1 i_4790 (.ZN (n_4726), .A1 (n_4727), .A2 (B_imm[2]), .A3 (A_imm[27]));
NAND2_X1 i_4789 (.ZN (n_4725), .A1 (n_4726), .A2 (n_5939));
INV_X1 i_4788 (.ZN (n_4724), .A (n_4725));
INV_X1 i_4787 (.ZN (n_4723), .A (n_5927));
NAND2_X1 i_4786 (.ZN (n_4722), .A1 (n_4723), .A2 (n_5939));
OAI21_X1 i_4785 (.ZN (n_4721), .A (n_4722), .B1 (n_4724), .B2 (n_5928));
INV_X1 i_4784 (.ZN (n_4720), .A (n_4721));
AOI21_X1 i_4783 (.ZN (n_4719), .A (n_4808), .B1 (n_4814), .B2 (n_4805));
INV_X1 i_4782 (.ZN (n_4718), .A (n_5905));
NAND2_X1 i_4781 (.ZN (n_4717), .A1 (n_5906), .A2 (n_5904));
NAND2_X1 i_4780 (.ZN (n_4716), .A1 (n_4717), .A2 (n_4718));
NAND3_X1 i_4779 (.ZN (n_4715), .A1 (n_5906), .A2 (n_5905), .A3 (n_5904));
NAND2_X1 i_4778 (.ZN (n_4714), .A1 (n_4716), .A2 (n_4715));
NAND2_X1 i_4777 (.ZN (n_4713), .A1 (n_4719), .A2 (n_4714));
NAND2_X1 i_4776 (.ZN (n_4712), .A1 (B_imm[9]), .A2 (A_imm[17]));
OAI21_X1 i_4775 (.ZN (n_4711), .A (n_4712), .B1 (n_8948), .B2 (n_6677));
OAI22_X1 i_4774 (.ZN (n_4710), .A1 (n_8946), .A2 (n_8880), .B1 (n_8909), .B2 (n_8511));
NAND2_X1 i_4773 (.ZN (n_4709), .A1 (B_imm[16]), .A2 (A_imm[9]));
INV_X1 i_4772 (.ZN (n_4708), .A (n_4709));
NAND4_X1 i_4771 (.ZN (n_4707), .A1 (A_imm[15]), .A2 (B_imm[17]), .A3 (B_imm[10]), .A4 (A_imm[8]));
INV_X1 i_4770 (.ZN (n_4706), .A (n_4707));
OAI21_X1 i_4769 (.ZN (n_4705), .A (n_4710), .B1 (n_4708), .B2 (n_4706));
INV_X1 i_4768 (.ZN (n_4704), .A (n_4705));
NAND4_X1 i_4767 (.ZN (n_4703), .A1 (B_imm[24]), .A2 (B_imm[9]), .A3 (A_imm[17]), .A4 (A_imm[2]));
INV_X1 i_4766 (.ZN (n_4702), .A (n_4703));
OAI21_X1 i_4765 (.ZN (n_4701), .A (n_4711), .B1 (n_4702), .B2 (n_4704));
NAND2_X1 i_4764 (.ZN (n_4700), .A1 (A_imm[26]), .A2 (B_imm[0]));
NAND2_X1 i_4763 (.ZN (n_4699), .A1 (A_imm[25]), .A2 (B_imm[1]));
NAND2_X1 i_4762 (.ZN (n_4698), .A1 (n_4700), .A2 (n_4699));
NAND2_X1 i_4761 (.ZN (n_4697), .A1 (B_imm[18]), .A2 (A_imm[8]));
INV_X1 i_4760 (.ZN (n_4696), .A (n_4697));
NAND4_X1 i_4759 (.ZN (n_4695), .A1 (A_imm[26]), .A2 (A_imm[25]), .A3 (B_imm[1]), .A4 (B_imm[0]));
INV_X1 i_4758 (.ZN (n_4694), .A (n_4695));
OAI21_X1 i_4757 (.ZN (n_4693), .A (n_4698), .B1 (n_4694), .B2 (n_4696));
NAND2_X1 i_4756 (.ZN (n_4692), .A1 (n_4701), .A2 (n_4693));
NAND2_X1 i_4755 (.ZN (n_4691), .A1 (B_imm[22]), .A2 (A_imm[4]));
OAI21_X1 i_4754 (.ZN (n_4690), .A (n_4691), .B1 (n_8829), .B2 (n_8926));
NAND2_X1 i_4753 (.ZN (n_4689), .A1 (B_imm[25]), .A2 (A_imm[1]));
INV_X1 i_4752 (.ZN (n_4688), .A (n_4689));
NAND4_X1 i_4751 (.ZN (n_4687), .A1 (B_imm[15]), .A2 (B_imm[22]), .A3 (A_imm[11]), .A4 (A_imm[4]));
INV_X1 i_4750 (.ZN (n_4686), .A (n_4687));
OAI21_X1 i_4749 (.ZN (n_4685), .A (n_4690), .B1 (n_4686), .B2 (n_4688));
OAI21_X1 i_4748 (.ZN (n_4684), .A (n_4685), .B1 (n_4701), .B2 (n_4693));
OAI211_X1 i_4747 (.ZN (n_4683), .A (n_4684), .B (n_4692), .C1 (n_4719), .C2 (n_4714));
INV_X1 i_4746 (.ZN (n_4682), .A (n_4743));
AOI22_X1 i_4745 (.ZN (n_4681), .A1 (n_4754), .A2 (n_4750), .B1 (n_4739), .B2 (n_4738));
NOR2_X1 i_4744 (.ZN (n_4680), .A1 (n_4681), .A2 (n_4682));
NAND3_X1 i_4743 (.ZN (n_4679), .A1 (n_4680), .A2 (n_4713), .A3 (n_4683));
INV_X1 i_4742 (.ZN (n_4678), .A (n_4679));
NAND2_X1 i_4741 (.ZN (n_4677), .A1 (n_4749), .A2 (n_4736));
AOI22_X1 i_4740 (.ZN (n_4676), .A1 (n_4683), .A2 (n_4713), .B1 (n_4743), .B2 (n_4677));
OAI21_X1 i_4739 (.ZN (n_4675), .A (n_4720), .B1 (n_4678), .B2 (n_4676));
NAND2_X1 i_4738 (.ZN (n_4674), .A1 (n_4683), .A2 (n_4713));
INV_X1 i_4737 (.ZN (n_4673), .A (n_4680));
NAND2_X1 i_4736 (.ZN (n_4672), .A1 (n_4674), .A2 (n_4673));
NAND3_X1 i_4735 (.ZN (n_4671), .A1 (n_4672), .A2 (n_4721), .A3 (n_4679));
NAND2_X1 i_4734 (.ZN (n_4670), .A1 (n_4675), .A2 (n_4671));
INV_X1 i_4733 (.ZN (n_4669), .A (n_4670));
NAND2_X1 i_4732 (.ZN (n_4668), .A1 (n_4728), .A2 (n_4669));
NAND2_X2 i_4731 (.ZN (n_4667), .A1 (n_4668), .A2 (n_4730));
NAND2_X2 i_4730 (.ZN (n_4666), .A1 (n_4667), .A2 (n_4866));
NAND2_X1 i_4729 (.ZN (n_4665), .A1 (n_4666), .A2 (n_4867));
NAND2_X1 i_4728 (.ZN (n_4664), .A1 (n_4665), .A2 (n_5009));
NAND3_X2 i_4727 (.ZN (n_4663), .A1 (n_4666), .A2 (n_5010), .A3 (n_4867));
INV_X1 i_4726 (.ZN (n_4662), .A (n_6155));
NAND2_X1 i_4725 (.ZN (n_4661), .A1 (n_6158), .A2 (n_6154));
NAND2_X1 i_4724 (.ZN (n_4660), .A1 (n_4661), .A2 (n_4662));
NAND3_X1 i_4723 (.ZN (n_4659), .A1 (n_6158), .A2 (n_6154), .A3 (n_6155));
NAND2_X1 i_4722 (.ZN (n_4658), .A1 (n_4660), .A2 (n_4659));
AOI21_X1 i_4721 (.ZN (n_4657), .A (n_6426), .B1 (n_6431), .B2 (n_6430));
NAND3_X1 i_4720 (.ZN (n_4656), .A1 (n_6430), .A2 (n_6431), .A3 (n_6426));
INV_X1 i_4719 (.ZN (n_4655), .A (n_4656));
OAI21_X1 i_4718 (.ZN (n_4654), .A (n_4658), .B1 (n_4657), .B2 (n_4655));
INV_X1 i_4717 (.ZN (n_4653), .A (n_4657));
NAND4_X1 i_4716 (.ZN (n_4652), .A1 (n_4660), .A2 (n_4653), .A3 (n_4659), .A4 (n_4656));
INV_X1 i_4715 (.ZN (n_4651), .A (n_4961));
INV_X1 i_4714 (.ZN (n_4650), .A (n_4955));
OAI21_X1 i_4713 (.ZN (n_4649), .A (n_4959), .B1 (n_4651), .B2 (n_4650));
NAND3_X1 i_4712 (.ZN (n_4648), .A1 (n_4654), .A2 (n_4652), .A3 (n_4649));
NAND2_X1 i_4711 (.ZN (n_4647), .A1 (n_4654), .A2 (n_4652));
INV_X1 i_4710 (.ZN (n_4646), .A (n_4649));
NAND2_X1 i_4709 (.ZN (n_4645), .A1 (n_4647), .A2 (n_4646));
NAND2_X1 i_4708 (.ZN (n_4644), .A1 (n_4645), .A2 (n_4648));
INV_X1 i_4707 (.ZN (n_4643), .A (n_4644));
NAND2_X2 i_4706 (.ZN (n_4642), .A1 (n_4663), .A2 (n_4643));
NAND2_X1 i_4705 (.ZN (n_4641), .A1 (n_4642), .A2 (n_4664));
INV_X1 i_4704 (.ZN (n_4640), .A (n_5042));
NAND2_X1 i_4703 (.ZN (n_4639), .A1 (n_5047), .A2 (n_5046));
NAND2_X1 i_4702 (.ZN (n_4638), .A1 (n_4639), .A2 (n_4640));
NAND3_X1 i_4701 (.ZN (n_4637), .A1 (n_5042), .A2 (n_5047), .A3 (n_5046));
NAND2_X1 i_4700 (.ZN (n_4636), .A1 (n_4638), .A2 (n_4637));
INV_X1 i_4699 (.ZN (n_4635), .A (n_4636));
NAND2_X1 i_4698 (.ZN (n_4634), .A1 (n_4641), .A2 (n_4635));
NAND3_X1 i_4697 (.ZN (n_4633), .A1 (n_4642), .A2 (n_4664), .A3 (n_4636));
AOI21_X1 i_4696 (.ZN (n_4632), .A (n_6146), .B1 (n_6194), .B2 (n_6147));
NAND3_X1 i_4695 (.ZN (n_4631), .A1 (n_6194), .A2 (n_6147), .A3 (n_6146));
INV_X1 i_4694 (.ZN (n_4630), .A (n_4631));
NAND2_X1 i_4693 (.ZN (n_4629), .A1 (n_4654), .A2 (n_4649));
OAI211_X1 i_4692 (.ZN (n_4628), .A (n_4629), .B (n_4652), .C1 (n_4630), .C2 (n_4632));
NOR2_X1 i_4691 (.ZN (n_4627), .A1 (n_4630), .A2 (n_4632));
NAND2_X1 i_4690 (.ZN (n_4626), .A1 (n_4629), .A2 (n_4652));
NAND2_X1 i_4689 (.ZN (n_4625), .A1 (n_4626), .A2 (n_4627));
OAI211_X1 i_4688 (.ZN (n_4624), .A (n_5871), .B (n_5864), .C1 (n_5916), .C2 (n_5915));
NAND3_X1 i_4687 (.ZN (n_4623), .A1 (n_5914), .A2 (n_5863), .A3 (n_5917));
NAND2_X1 i_4686 (.ZN (n_4622), .A1 (n_4624), .A2 (n_4623));
NAND3_X1 i_4685 (.ZN (n_4621), .A1 (n_4625), .A2 (n_4628), .A3 (n_4622));
NAND2_X1 i_4684 (.ZN (n_4620), .A1 (n_4625), .A2 (n_4628));
INV_X1 i_4683 (.ZN (n_4619), .A (n_4622));
NAND2_X1 i_4682 (.ZN (n_4618), .A1 (n_4620), .A2 (n_4619));
NAND2_X1 i_4681 (.ZN (n_4617), .A1 (n_4618), .A2 (n_4621));
NAND2_X1 i_4680 (.ZN (n_4616), .A1 (n_4633), .A2 (n_4617));
NAND2_X2 i_4679 (.ZN (n_4615), .A1 (n_4616), .A2 (n_4634));
INV_X1 i_4678 (.ZN (n_4614), .A (n_4615));
NAND2_X1 i_4677 (.ZN (n_4613), .A1 (n_5014), .A2 (n_4614));
NAND3_X1 i_4676 (.ZN (n_4612), .A1 (n_4615), .A2 (n_5019), .A3 (n_5015));
NAND2_X1 i_4675 (.ZN (n_4611), .A1 (n_4613), .A2 (n_4612));
NAND3_X1 i_4674 (.ZN (n_4610), .A1 (n_6151), .A2 (n_6144), .A3 (n_6127));
INV_X1 i_4673 (.ZN (n_4609), .A (n_4610));
AOI21_X1 i_4672 (.ZN (n_4608), .A (n_6127), .B1 (n_6151), .B2 (n_6144));
NAND2_X1 i_4671 (.ZN (n_4607), .A1 (n_4628), .A2 (n_4619));
OAI211_X1 i_4670 (.ZN (n_4606), .A (n_4607), .B (n_4625), .C1 (n_4609), .C2 (n_4608));
NOR2_X1 i_4669 (.ZN (n_4605), .A1 (n_4608), .A2 (n_4609));
NAND2_X1 i_4668 (.ZN (n_4604), .A1 (n_4607), .A2 (n_4625));
NAND2_X1 i_4667 (.ZN (n_4603), .A1 (n_4604), .A2 (n_4605));
NAND2_X1 i_4666 (.ZN (n_4602), .A1 (n_4603), .A2 (n_4606));
NAND3_X1 i_4665 (.ZN (n_4601), .A1 (n_5757), .A2 (n_5756), .A3 (n_5753));
AOI21_X1 i_4664 (.ZN (n_4600), .A (n_5854), .B1 (n_5759), .B2 (n_5821));
OAI21_X1 i_4663 (.ZN (n_4599), .A (n_5752), .B1 (n_5755), .B2 (n_4600));
NAND3_X1 i_4662 (.ZN (n_4598), .A1 (n_5958), .A2 (n_5954), .A3 (n_5923));
INV_X1 i_4661 (.ZN (n_4597), .A (n_4598));
AOI21_X1 i_4660 (.ZN (n_4596), .A (n_5923), .B1 (n_5958), .B2 (n_5954));
AOI21_X1 i_4659 (.ZN (n_4595), .A (n_5874), .B1 (n_5878), .B2 (n_5881));
NAND3_X1 i_4658 (.ZN (n_4594), .A1 (n_5878), .A2 (n_5881), .A3 (n_5874));
INV_X1 i_4657 (.ZN (n_4593), .A (n_4594));
NOR2_X1 i_4656 (.ZN (n_4592), .A1 (n_4595), .A2 (n_4593));
NAND2_X1 i_4655 (.ZN (n_4591), .A1 (n_4862), .A2 (n_4855));
NAND2_X1 i_4654 (.ZN (n_4590), .A1 (n_4591), .A2 (n_4852));
NAND2_X1 i_4653 (.ZN (n_4589), .A1 (n_4592), .A2 (n_4590));
OAI211_X2 i_4652 (.ZN (n_4588), .A (n_4852), .B (n_4591), .C1 (n_4595), .C2 (n_4593));
NAND2_X1 i_4651 (.ZN (n_4587), .A1 (n_4679), .A2 (n_4721));
NAND2_X1 i_4650 (.ZN (n_4586), .A1 (n_4587), .A2 (n_4672));
NAND2_X1 i_4649 (.ZN (n_4585), .A1 (n_4588), .A2 (n_4586));
NAND2_X1 i_4648 (.ZN (n_4584), .A1 (n_4585), .A2 (n_4589));
OAI21_X1 i_4647 (.ZN (n_4583), .A (n_4584), .B1 (n_4597), .B2 (n_4596));
NOR2_X1 i_4646 (.ZN (n_4582), .A1 (n_4597), .A2 (n_4596));
NAND3_X1 i_4645 (.ZN (n_4581), .A1 (n_4582), .A2 (n_4589), .A3 (n_4585));
NAND3_X1 i_4644 (.ZN (n_4580), .A1 (n_5871), .A2 (n_5870), .A3 (n_5865));
INV_X1 i_4643 (.ZN (n_4579), .A (n_4580));
AOI21_X1 i_4642 (.ZN (n_4578), .A (n_5865), .B1 (n_5871), .B2 (n_5870));
NOR2_X1 i_4641 (.ZN (n_4577), .A1 (n_4579), .A2 (n_4578));
NAND2_X1 i_4640 (.ZN (n_4576), .A1 (n_4581), .A2 (n_4577));
NAND2_X2 i_4639 (.ZN (n_4575), .A1 (n_4576), .A2 (n_4583));
NAND3_X1 i_4638 (.ZN (n_4574), .A1 (n_4575), .A2 (n_4601), .A3 (n_4599));
NAND2_X1 i_4637 (.ZN (n_4573), .A1 (n_4599), .A2 (n_4601));
INV_X1 i_4636 (.ZN (n_4572), .A (n_4575));
NAND2_X1 i_4635 (.ZN (n_4571), .A1 (n_4573), .A2 (n_4572));
INV_X1 i_4634 (.ZN (n_4570), .A (n_5760));
NAND2_X1 i_4633 (.ZN (n_4569), .A1 (n_5818), .A2 (n_5821));
NAND2_X1 i_4632 (.ZN (n_4568), .A1 (n_4569), .A2 (n_4570));
NAND3_X1 i_4631 (.ZN (n_4567), .A1 (n_5760), .A2 (n_5818), .A3 (n_5821));
NAND3_X1 i_4630 (.ZN (n_4566), .A1 (n_5948), .A2 (n_5926), .A3 (n_5925));
NAND2_X1 i_4629 (.ZN (n_4565), .A1 (n_5948), .A2 (n_5925));
NAND3_X1 i_4628 (.ZN (n_4564), .A1 (n_4565), .A2 (n_5939), .A3 (n_5927));
NAND2_X1 i_4627 (.ZN (n_4563), .A1 (n_4564), .A2 (n_4566));
INV_X1 i_4626 (.ZN (n_4562), .A (n_5893));
OAI21_X1 i_4625 (.ZN (n_4561), .A (n_5891), .B1 (n_4562), .B2 (n_5889));
NAND3_X1 i_4624 (.ZN (n_4560), .A1 (n_5893), .A2 (n_5892), .A3 (n_5890));
NAND2_X1 i_4623 (.ZN (n_4559), .A1 (n_4561), .A2 (n_4560));
AOI22_X1 i_4622 (.ZN (n_4558), .A1 (n_5938), .A2 (n_5935), .B1 (B_imm[23]), .B2 (A_imm[5]));
OAI21_X1 i_4621 (.ZN (n_4557), .A (n_5931), .B1 (n_5929), .B2 (n_4558));
NAND3_X1 i_4620 (.ZN (n_4556), .A1 (n_5933), .A2 (n_5932), .A3 (n_5930));
NAND2_X1 i_4619 (.ZN (n_4555), .A1 (n_4556), .A2 (n_4557));
NAND2_X1 i_4618 (.ZN (n_4554), .A1 (n_4559), .A2 (n_4555));
NAND4_X1 i_4617 (.ZN (n_4553), .A1 (n_4561), .A2 (n_4557), .A3 (n_4556), .A4 (n_4560));
INV_X1 i_4616 (.ZN (n_4552), .A (n_4553));
NAND2_X1 i_4615 (.ZN (n_4551), .A1 (n_5945), .A2 (n_5942));
NAND2_X1 i_4614 (.ZN (n_4550), .A1 (n_4551), .A2 (n_5943));
INV_X1 i_4613 (.ZN (n_4549), .A (n_4551));
NAND2_X1 i_4612 (.ZN (n_4548), .A1 (n_4549), .A2 (n_5944));
NAND2_X1 i_4611 (.ZN (n_4547), .A1 (n_4548), .A2 (n_4550));
INV_X1 i_4610 (.ZN (n_4546), .A (n_4547));
OAI21_X1 i_4609 (.ZN (n_4545), .A (n_4554), .B1 (n_4552), .B2 (n_4546));
NAND3_X1 i_4608 (.ZN (n_4544), .A1 (n_5838), .A2 (n_5836), .A3 (n_5832));
INV_X1 i_4607 (.ZN (n_4543), .A (n_5832));
NAND2_X1 i_4606 (.ZN (n_4542), .A1 (n_5838), .A2 (n_5836));
NAND2_X1 i_4605 (.ZN (n_4541), .A1 (n_4542), .A2 (n_4543));
NAND2_X1 i_4604 (.ZN (n_4540), .A1 (n_4541), .A2 (n_4544));
NAND2_X1 i_4603 (.ZN (n_4539), .A1 (n_4545), .A2 (n_4540));
NAND2_X1 i_4602 (.ZN (n_4538), .A1 (n_4553), .A2 (n_4547));
NAND4_X1 i_4601 (.ZN (n_4537), .A1 (n_4538), .A2 (n_4554), .A3 (n_4544), .A4 (n_4541));
AOI21_X1 i_4600 (.ZN (n_4536), .A (n_5794), .B1 (n_5803), .B2 (n_5798));
NAND3_X1 i_4599 (.ZN (n_4535), .A1 (n_5798), .A2 (n_5803), .A3 (n_5794));
INV_X1 i_4598 (.ZN (n_4534), .A (n_4535));
NOR2_X2 i_4597 (.ZN (n_4533), .A1 (n_4534), .A2 (n_4536));
NAND2_X1 i_4596 (.ZN (n_4532), .A1 (n_4537), .A2 (n_4533));
NAND2_X1 i_4595 (.ZN (n_4531), .A1 (n_4532), .A2 (n_4539));
NAND2_X1 i_4594 (.ZN (n_4530), .A1 (n_4531), .A2 (n_4563));
NAND4_X1 i_4593 (.ZN (n_4529), .A1 (n_4532), .A2 (n_4566), .A3 (n_4564), .A4 (n_4539));
NAND3_X1 i_4592 (.ZN (n_4528), .A1 (n_5829), .A2 (n_5825), .A3 (n_5823));
NAND2_X1 i_4591 (.ZN (n_4527), .A1 (n_5829), .A2 (n_5823));
OAI21_X1 i_4590 (.ZN (n_4526), .A (n_4527), .B1 (n_5828), .B2 (n_5826));
NAND2_X1 i_4589 (.ZN (n_4525), .A1 (n_4526), .A2 (n_4528));
NAND2_X1 i_4588 (.ZN (n_4524), .A1 (n_4529), .A2 (n_4525));
NAND2_X1 i_4587 (.ZN (n_4523), .A1 (n_4524), .A2 (n_4530));
NAND3_X1 i_4586 (.ZN (n_4522), .A1 (n_4523), .A2 (n_4568), .A3 (n_4567));
NAND2_X1 i_4585 (.ZN (n_4521), .A1 (n_4568), .A2 (n_4567));
NAND3_X1 i_4584 (.ZN (n_4520), .A1 (n_4521), .A2 (n_4530), .A3 (n_4524));
INV_X1 i_4583 (.ZN (n_4519), .A (n_5762));
NAND2_X1 i_4582 (.ZN (n_4518), .A1 (n_5791), .A2 (n_5790));
NAND2_X1 i_4581 (.ZN (n_4517), .A1 (n_4518), .A2 (n_4519));
NAND3_X1 i_4580 (.ZN (n_4516), .A1 (n_5762), .A2 (n_5791), .A3 (n_5790));
NAND2_X1 i_4579 (.ZN (n_4515), .A1 (n_4517), .A2 (n_4516));
INV_X1 i_4578 (.ZN (n_4514), .A (n_4515));
AOI21_X1 i_4577 (.ZN (n_4513), .A (n_5764), .B1 (n_5768), .B2 (n_5771));
NAND3_X1 i_4576 (.ZN (n_4512), .A1 (n_5768), .A2 (n_5771), .A3 (n_5764));
INV_X1 i_4575 (.ZN (n_4511), .A (n_4512));
NOR2_X1 i_4574 (.ZN (n_4510), .A1 (n_4513), .A2 (n_4511));
NAND2_X1 i_4573 (.ZN (n_4509), .A1 (n_5807), .A2 (n_5805));
NAND2_X1 i_4572 (.ZN (n_4508), .A1 (n_4509), .A2 (n_5801));
NAND3_X1 i_4571 (.ZN (n_4507), .A1 (n_5807), .A2 (n_5806), .A3 (n_5805));
NAND2_X1 i_4570 (.ZN (n_4506), .A1 (n_4508), .A2 (n_4507));
NAND2_X1 i_4569 (.ZN (n_4505), .A1 (B_imm[13]), .A2 (A_imm[13]));
OAI21_X1 i_4568 (.ZN (n_4504), .A (n_4505), .B1 (n_8860), .B2 (n_7691));
NAND2_X1 i_4567 (.ZN (n_4503), .A1 (B_imm[26]), .A2 (A_imm[0]));
NAND4_X1 i_4566 (.ZN (n_4502), .A1 (B_imm[20]), .A2 (B_imm[13]), .A3 (A_imm[13]), .A4 (A_imm[6]));
NAND2_X1 i_4565 (.ZN (n_4501), .A1 (n_4502), .A2 (n_4503));
NAND4_X1 i_4564 (.ZN (n_4500), .A1 (n_4501), .A2 (B_imm[0]), .A3 (A_imm[27]), .A4 (n_4504));
AOI22_X1 i_4563 (.ZN (n_4499), .A1 (n_4501), .A2 (n_4504), .B1 (A_imm[27]), .B2 (B_imm[0]));
AOI21_X1 i_4562 (.ZN (n_4498), .A (n_5937), .B1 (n_5938), .B2 (n_5936));
NAND3_X1 i_4561 (.ZN (n_4497), .A1 (n_5938), .A2 (n_5937), .A3 (n_5936));
INV_X1 i_4560 (.ZN (n_4496), .A (n_4497));
NOR2_X1 i_4559 (.ZN (n_4495), .A1 (n_4498), .A2 (n_4496));
OAI21_X1 i_4558 (.ZN (n_4494), .A (n_4500), .B1 (n_4499), .B2 (n_4495));
NAND2_X1 i_4557 (.ZN (n_4493), .A1 (n_4506), .A2 (n_4494));
NAND2_X1 i_4556 (.ZN (n_4492), .A1 (B_imm[23]), .A2 (A_imm[3]));
NAND2_X1 i_4555 (.ZN (n_4491), .A1 (A_imm[22]), .A2 (B_imm[3]));
OAI21_X1 i_4554 (.ZN (n_4490), .A (n_4491), .B1 (n_8859), .B2 (n_6577));
NAND2_X1 i_4553 (.ZN (n_4489), .A1 (A_imm[18]), .A2 (B_imm[7]));
INV_X1 i_4552 (.ZN (n_4488), .A (n_4489));
NAND4_X1 i_4551 (.ZN (n_4487), .A1 (A_imm[21]), .A2 (A_imm[22]), .A3 (B_imm[4]), .A4 (B_imm[3]));
INV_X1 i_4550 (.ZN (n_4486), .A (n_4487));
OAI21_X1 i_4549 (.ZN (n_4485), .A (n_4490), .B1 (n_4486), .B2 (n_4488));
NAND2_X1 i_4548 (.ZN (n_4484), .A1 (n_4485), .A2 (n_4492));
NAND2_X1 i_4547 (.ZN (n_4483), .A1 (B_imm[21]), .A2 (A_imm[5]));
OAI21_X1 i_4546 (.ZN (n_4482), .A (n_4483), .B1 (n_4485), .B2 (n_4492));
NAND4_X1 i_4545 (.ZN (n_4481), .A1 (n_4482), .A2 (B_imm[14]), .A3 (A_imm[13]), .A4 (n_4484));
AOI22_X1 i_4544 (.ZN (n_4480), .A1 (n_4484), .A2 (n_4482), .B1 (B_imm[14]), .B2 (A_imm[13]));
NAND2_X1 i_4543 (.ZN (n_4479), .A1 (n_5812), .A2 (n_5810));
XNOR2_X1 i_4542 (.ZN (n_4478), .A (n_4479), .B (n_5811));
OAI21_X1 i_4541 (.ZN (n_4477), .A (n_4481), .B1 (n_4480), .B2 (n_4478));
OAI21_X1 i_4540 (.ZN (n_4476), .A (n_4477), .B1 (n_4506), .B2 (n_4494));
NAND2_X1 i_4539 (.ZN (n_4475), .A1 (n_4476), .A2 (n_4493));
NAND2_X1 i_4538 (.ZN (n_4474), .A1 (n_4510), .A2 (n_4475));
OAI211_X1 i_4537 (.ZN (n_4473), .A (n_4476), .B (n_4493), .C1 (n_4513), .C2 (n_4511));
INV_X1 i_4536 (.ZN (n_4472), .A (n_5778));
NAND2_X1 i_4535 (.ZN (n_4471), .A1 (n_5784), .A2 (n_5777));
NAND2_X1 i_4534 (.ZN (n_4470), .A1 (n_4471), .A2 (n_4472));
NAND3_X1 i_4533 (.ZN (n_4469), .A1 (n_5784), .A2 (n_5777), .A3 (n_5778));
NAND2_X1 i_4532 (.ZN (n_4468), .A1 (n_4470), .A2 (n_4469));
INV_X1 i_4531 (.ZN (n_4467), .A (n_5078));
INV_X1 i_4530 (.ZN (n_4466), .A (n_5077));
OAI21_X1 i_4529 (.ZN (n_4465), .A (n_4467), .B1 (n_4466), .B2 (n_5086));
NAND3_X1 i_4528 (.ZN (n_4464), .A1 (n_5085), .A2 (n_5077), .A3 (n_5078));
NAND2_X1 i_4527 (.ZN (n_4463), .A1 (n_4465), .A2 (n_4464));
NAND2_X1 i_4526 (.ZN (n_4462), .A1 (n_4463), .A2 (n_4468));
NAND4_X1 i_4525 (.ZN (n_4461), .A1 (n_4465), .A2 (n_4470), .A3 (n_4464), .A4 (n_4469));
NAND2_X1 i_4524 (.ZN (n_4460), .A1 (B_imm[6]), .A2 (A_imm[19]));
OAI21_X1 i_4523 (.ZN (n_4459), .A (n_4460), .B1 (n_8893), .B2 (n_8429));
NAND2_X1 i_4522 (.ZN (n_4458), .A1 (B_imm[8]), .A2 (A_imm[17]));
NAND4_X1 i_4521 (.ZN (n_4457), .A1 (A_imm[20]), .A2 (B_imm[6]), .A3 (B_imm[5]), .A4 (A_imm[19]));
NAND2_X1 i_4520 (.ZN (n_4456), .A1 (n_4457), .A2 (n_4458));
AOI22_X1 i_4519 (.ZN (n_4455), .A1 (n_4456), .A2 (n_4459), .B1 (B_imm[19]), .B2 (A_imm[7]));
INV_X1 i_4518 (.ZN (n_4454), .A (n_4455));
NAND4_X1 i_4517 (.ZN (n_4453), .A1 (n_4456), .A2 (B_imm[19]), .A3 (A_imm[7]), .A4 (n_4459));
NAND2_X1 i_4516 (.ZN (n_4452), .A1 (A_imm[24]), .A2 (B_imm[1]));
OAI21_X1 i_4515 (.ZN (n_4451), .A (n_4452), .B1 (n_8907), .B2 (n_6584));
NAND2_X1 i_4514 (.ZN (n_4450), .A1 (B_imm[12]), .A2 (A_imm[13]));
INV_X1 i_4513 (.ZN (n_4449), .A (n_4450));
NAND4_X1 i_4512 (.ZN (n_4448), .A1 (A_imm[23]), .A2 (A_imm[24]), .A3 (B_imm[2]), .A4 (B_imm[1]));
INV_X1 i_4511 (.ZN (n_4447), .A (n_4448));
OAI21_X1 i_4510 (.ZN (n_4446), .A (n_4451), .B1 (n_4447), .B2 (n_4449));
NAND2_X1 i_4509 (.ZN (n_4445), .A1 (n_4453), .A2 (n_4446));
AOI21_X1 i_4508 (.ZN (n_4444), .A (n_5788), .B1 (n_5789), .B2 (n_5787));
NAND3_X1 i_4507 (.ZN (n_4443), .A1 (n_5789), .A2 (n_5788), .A3 (n_5787));
INV_X1 i_4506 (.ZN (n_4442), .A (n_4443));
OAI211_X1 i_4505 (.ZN (n_4441), .A (n_4445), .B (n_4454), .C1 (n_4444), .C2 (n_4442));
NAND2_X1 i_4504 (.ZN (n_4440), .A1 (n_4445), .A2 (n_4454));
NOR2_X1 i_4503 (.ZN (n_4439), .A1 (n_4444), .A2 (n_4442));
NAND2_X1 i_4502 (.ZN (n_4438), .A1 (n_4440), .A2 (n_4439));
INV_X1 i_4501 (.ZN (n_4437), .A (n_4438));
NAND2_X1 i_4500 (.ZN (n_4436), .A1 (n_5783), .A2 (n_5780));
XNOR2_X1 i_4499 (.ZN (n_4435), .A (n_4436), .B (n_5782));
OAI21_X1 i_4498 (.ZN (n_4434), .A (n_4441), .B1 (n_4437), .B2 (n_4435));
NAND2_X1 i_4497 (.ZN (n_4433), .A1 (n_4434), .A2 (n_4461));
NAND2_X1 i_4496 (.ZN (n_4432), .A1 (n_4433), .A2 (n_4462));
NAND2_X1 i_4495 (.ZN (n_4431), .A1 (n_4473), .A2 (n_4432));
NAND2_X1 i_4494 (.ZN (n_4430), .A1 (n_4431), .A2 (n_4474));
NAND2_X1 i_4493 (.ZN (n_4429), .A1 (n_4430), .A2 (n_4514));
NAND3_X1 i_4492 (.ZN (n_4428), .A1 (n_4515), .A2 (n_4431), .A3 (n_4474));
INV_X1 i_4491 (.ZN (n_4427), .A (n_4428));
INV_X1 i_4490 (.ZN (n_4426), .A (n_5052));
NAND2_X1 i_4489 (.ZN (n_4425), .A1 (n_5058), .A2 (n_5056));
NAND2_X1 i_4488 (.ZN (n_4424), .A1 (n_4425), .A2 (n_4426));
NAND3_X1 i_4487 (.ZN (n_4423), .A1 (n_5058), .A2 (n_5056), .A3 (n_5052));
NAND2_X1 i_4486 (.ZN (n_4422), .A1 (n_4424), .A2 (n_4423));
OAI21_X1 i_4485 (.ZN (n_4421), .A (n_4429), .B1 (n_4427), .B2 (n_4422));
NAND2_X1 i_4484 (.ZN (n_4420), .A1 (n_4520), .A2 (n_4421));
NAND2_X1 i_4483 (.ZN (n_4419), .A1 (n_4420), .A2 (n_4522));
NAND2_X1 i_4482 (.ZN (n_4418), .A1 (n_4571), .A2 (n_4419));
NAND3_X1 i_4481 (.ZN (n_4417), .A1 (n_4602), .A2 (n_4574), .A3 (n_4418));
NAND2_X1 i_4480 (.ZN (n_4416), .A1 (n_4418), .A2 (n_4574));
NAND3_X1 i_4479 (.ZN (n_4415), .A1 (n_4416), .A2 (n_4606), .A3 (n_4603));
NAND2_X1 i_4478 (.ZN (n_4414), .A1 (n_4417), .A2 (n_4415));
NAND2_X1 i_4477 (.ZN (n_4413), .A1 (n_4611), .A2 (n_4414));
INV_X1 i_4476 (.ZN (n_4412), .A (n_4414));
NAND3_X1 i_4475 (.ZN (n_4411), .A1 (n_4613), .A2 (n_4412), .A3 (n_4612));
INV_X1 i_4474 (.ZN (n_4410), .A (n_4411));
INV_X1 i_4473 (.ZN (n_4409), .A (n_4577));
NAND3_X1 i_4472 (.ZN (n_4408), .A1 (n_4583), .A2 (n_4409), .A3 (n_4581));
NAND2_X1 i_4471 (.ZN (n_4407), .A1 (n_5958), .A2 (n_5954));
NAND3_X1 i_4470 (.ZN (n_4406), .A1 (n_4407), .A2 (n_5948), .A3 (n_5924));
AOI22_X1 i_4469 (.ZN (n_4405), .A1 (n_4585), .A2 (n_4589), .B1 (n_4598), .B2 (n_4406));
INV_X1 i_4468 (.ZN (n_4404), .A (n_4581));
OAI21_X1 i_4467 (.ZN (n_4403), .A (n_4577), .B1 (n_4404), .B2 (n_4405));
NAND2_X1 i_4466 (.ZN (n_4402), .A1 (n_4403), .A2 (n_4408));
AOI21_X1 i_4465 (.ZN (n_4401), .A (n_4525), .B1 (n_4530), .B2 (n_4529));
INV_X1 i_4464 (.ZN (n_4400), .A (n_4401));
NAND3_X1 i_4463 (.ZN (n_4399), .A1 (n_4530), .A2 (n_4529), .A3 (n_4525));
AOI21_X1 i_4462 (.ZN (n_4398), .A (n_4586), .B1 (n_4589), .B2 (n_4588));
NAND3_X1 i_4461 (.ZN (n_4397), .A1 (n_4589), .A2 (n_4588), .A3 (n_4586));
INV_X1 i_4460 (.ZN (n_4396), .A (n_4397));
NOR2_X1 i_4459 (.ZN (n_4395), .A1 (n_4396), .A2 (n_4398));
NAND3_X1 i_4458 (.ZN (n_4394), .A1 (n_4395), .A2 (n_4400), .A3 (n_4399));
INV_X1 i_4457 (.ZN (n_4393), .A (n_4399));
OAI22_X1 i_4456 (.ZN (n_4392), .A1 (n_4393), .A2 (n_4401), .B1 (n_4396), .B2 (n_4398));
NAND3_X1 i_4455 (.ZN (n_4391), .A1 (n_4539), .A2 (n_4533), .A3 (n_4537));
INV_X1 i_4454 (.ZN (n_4390), .A (n_4533));
NAND2_X1 i_4453 (.ZN (n_4389), .A1 (n_4539), .A2 (n_4537));
NAND2_X1 i_4452 (.ZN (n_4388), .A1 (n_4389), .A2 (n_4390));
NAND2_X1 i_4451 (.ZN (n_4387), .A1 (n_4388), .A2 (n_4391));
INV_X1 i_4450 (.ZN (n_4386), .A (n_4387));
NAND2_X1 i_4449 (.ZN (n_4385), .A1 (n_4805), .A2 (n_4814));
NAND2_X1 i_4448 (.ZN (n_4384), .A1 (n_4385), .A2 (n_4802));
NAND3_X1 i_4447 (.ZN (n_4383), .A1 (n_4384), .A2 (n_4716), .A3 (n_4715));
NAND4_X1 i_4446 (.ZN (n_4382), .A1 (n_4383), .A2 (n_4713), .A3 (n_4692), .A4 (n_4684));
NAND2_X1 i_4445 (.ZN (n_4381), .A1 (n_4684), .A2 (n_4692));
NAND2_X1 i_4444 (.ZN (n_4380), .A1 (n_4713), .A2 (n_4383));
NAND2_X1 i_4443 (.ZN (n_4379), .A1 (n_4380), .A2 (n_4381));
NAND2_X2 i_4442 (.ZN (n_4378), .A1 (n_4379), .A2 (n_4382));
INV_X1 i_4441 (.ZN (n_4377), .A (n_4378));
NAND2_X1 i_4440 (.ZN (n_4376), .A1 (n_4819), .A2 (n_4816));
NAND2_X1 i_4439 (.ZN (n_4375), .A1 (n_4376), .A2 (n_4817));
NAND3_X1 i_4438 (.ZN (n_4374), .A1 (n_4819), .A2 (n_4818), .A3 (n_4816));
NAND2_X1 i_4437 (.ZN (n_4373), .A1 (n_4375), .A2 (n_4374));
INV_X1 i_4436 (.ZN (n_4372), .A (n_4698));
OAI21_X1 i_4435 (.ZN (n_4371), .A (n_4696), .B1 (n_4372), .B2 (n_4694));
NAND3_X1 i_4434 (.ZN (n_4370), .A1 (n_4698), .A2 (n_4695), .A3 (n_4697));
NAND2_X1 i_4433 (.ZN (n_4369), .A1 (n_4371), .A2 (n_4370));
NAND2_X1 i_4432 (.ZN (n_4368), .A1 (n_4369), .A2 (n_4373));
NAND4_X1 i_4431 (.ZN (n_4367), .A1 (n_4371), .A2 (n_4375), .A3 (n_4374), .A4 (n_4370));
INV_X2 i_4430 (.ZN (n_4366), .A (B_imm[1]));
NAND2_X1 i_4429 (.ZN (n_4365), .A1 (B_imm[8]), .A2 (A_imm[16]));
OAI21_X1 i_4428 (.ZN (n_4364), .A (n_4365), .B1 (n_8907), .B2 (n_4366));
NAND2_X1 i_4427 (.ZN (n_4363), .A1 (A_imm[24]), .A2 (B_imm[0]));
NAND4_X1 i_4426 (.ZN (n_4362), .A1 (A_imm[23]), .A2 (B_imm[8]), .A3 (B_imm[1]), .A4 (A_imm[16]));
NAND2_X1 i_4425 (.ZN (n_4361), .A1 (n_4362), .A2 (n_4363));
AOI22_X1 i_4424 (.ZN (n_4360), .A1 (n_4361), .A2 (n_4364), .B1 (B_imm[19]), .B2 (A_imm[6]));
INV_X1 i_4423 (.ZN (n_4359), .A (n_4360));
NAND4_X1 i_4422 (.ZN (n_4358), .A1 (n_4361), .A2 (B_imm[19]), .A3 (A_imm[6]), .A4 (n_4364));
INV_X1 i_4421 (.ZN (n_4357), .A (n_4358));
NAND2_X1 i_4420 (.ZN (n_4356), .A1 (B_imm[12]), .A2 (A_imm[12]));
OAI21_X1 i_4419 (.ZN (n_4355), .A (n_4356), .B1 (n_8849), .B2 (n_8927));
NAND2_X1 i_4418 (.ZN (n_4354), .A1 (B_imm[18]), .A2 (A_imm[6]));
INV_X1 i_4417 (.ZN (n_4353), .A (n_4354));
NAND4_X1 i_4416 (.ZN (n_4352), .A1 (B_imm[11]), .A2 (B_imm[12]), .A3 (A_imm[13]), .A4 (A_imm[12]));
INV_X1 i_4415 (.ZN (n_4351), .A (n_4352));
OAI21_X1 i_4414 (.ZN (n_4350), .A (n_4355), .B1 (n_4351), .B2 (n_4353));
INV_X1 i_4413 (.ZN (n_4349), .A (n_4350));
OAI21_X1 i_4412 (.ZN (n_4348), .A (n_4359), .B1 (n_4349), .B2 (n_4357));
INV_X1 i_4411 (.ZN (n_4347), .A (n_4348));
NAND2_X1 i_4410 (.ZN (n_4346), .A1 (n_4367), .A2 (n_4347));
NAND2_X1 i_4409 (.ZN (n_4345), .A1 (n_4346), .A2 (n_4368));
INV_X1 i_4408 (.ZN (n_4344), .A (n_4685));
NAND2_X1 i_4407 (.ZN (n_4343), .A1 (n_4703), .A2 (n_4705));
NAND2_X1 i_4406 (.ZN (n_4342), .A1 (n_4695), .A2 (n_4697));
NAND4_X1 i_4405 (.ZN (n_4341), .A1 (n_4343), .A2 (n_4342), .A3 (n_4711), .A4 (n_4698));
NAND2_X1 i_4404 (.ZN (n_4340), .A1 (n_4692), .A2 (n_4341));
NAND2_X1 i_4403 (.ZN (n_4339), .A1 (n_4340), .A2 (n_4344));
NAND3_X1 i_4402 (.ZN (n_4338), .A1 (n_4692), .A2 (n_4341), .A3 (n_4685));
NAND2_X1 i_4401 (.ZN (n_4337), .A1 (n_4339), .A2 (n_4338));
NAND2_X1 i_4400 (.ZN (n_4336), .A1 (n_4345), .A2 (n_4337));
NAND4_X1 i_4399 (.ZN (n_4335), .A1 (n_4346), .A2 (n_4339), .A3 (n_4368), .A4 (n_4338));
INV_X1 i_4398 (.ZN (n_4334), .A (n_4499));
INV_X1 i_4397 (.ZN (n_4333), .A (n_4495));
AOI21_X1 i_4396 (.ZN (n_4332), .A (n_4333), .B1 (n_4334), .B2 (n_4500));
NAND3_X1 i_4395 (.ZN (n_4331), .A1 (n_4334), .A2 (n_4500), .A3 (n_4333));
INV_X1 i_4394 (.ZN (n_4330), .A (n_4331));
NOR2_X1 i_4393 (.ZN (n_4329), .A1 (n_4330), .A2 (n_4332));
NAND2_X1 i_4392 (.ZN (n_4328), .A1 (n_4335), .A2 (n_4329));
NAND2_X1 i_4391 (.ZN (n_4327), .A1 (n_4328), .A2 (n_4336));
NAND2_X1 i_4390 (.ZN (n_4326), .A1 (n_4327), .A2 (n_4377));
NAND3_X1 i_4389 (.ZN (n_4325), .A1 (n_4328), .A2 (n_4378), .A3 (n_4336));
NAND2_X1 i_4388 (.ZN (n_4324), .A1 (n_4554), .A2 (n_4553));
XNOR2_X1 i_4387 (.ZN (n_4323), .A (n_4324), .B (n_4547));
NAND2_X2 i_4386 (.ZN (n_4322), .A1 (n_4325), .A2 (n_4323));
NAND2_X1 i_4385 (.ZN (n_4321), .A1 (n_4322), .A2 (n_4326));
NAND2_X1 i_4384 (.ZN (n_4320), .A1 (n_4321), .A2 (n_4386));
NAND3_X1 i_4383 (.ZN (n_4319), .A1 (n_4387), .A2 (n_4326), .A3 (n_4322));
INV_X1 i_4382 (.ZN (n_4318), .A (n_4319));
NAND2_X1 i_4381 (.ZN (n_4317), .A1 (n_4474), .A2 (n_4473));
NAND3_X1 i_4380 (.ZN (n_4316), .A1 (n_4317), .A2 (n_4462), .A3 (n_4433));
NAND3_X1 i_4379 (.ZN (n_4315), .A1 (n_4474), .A2 (n_4473), .A3 (n_4432));
NAND2_X1 i_4378 (.ZN (n_4314), .A1 (n_4316), .A2 (n_4315));
OAI21_X1 i_4377 (.ZN (n_4313), .A (n_4320), .B1 (n_4314), .B2 (n_4318));
NAND2_X2 i_4376 (.ZN (n_4312), .A1 (n_4313), .A2 (n_4392));
NAND2_X1 i_4375 (.ZN (n_4311), .A1 (n_4312), .A2 (n_4394));
NAND2_X1 i_4374 (.ZN (n_4310), .A1 (n_4311), .A2 (n_4402));
NAND4_X2 i_4373 (.ZN (n_4309), .A1 (n_4312), .A2 (n_4408), .A3 (n_4403), .A4 (n_4394));
NAND3_X1 i_4372 (.ZN (n_4308), .A1 (n_4522), .A2 (n_4421), .A3 (n_4520));
INV_X1 i_4371 (.ZN (n_4307), .A (n_4421));
NAND2_X1 i_4370 (.ZN (n_4306), .A1 (n_4520), .A2 (n_4522));
NAND2_X1 i_4369 (.ZN (n_4305), .A1 (n_4306), .A2 (n_4307));
NAND2_X1 i_4368 (.ZN (n_4304), .A1 (n_4305), .A2 (n_4308));
INV_X1 i_4367 (.ZN (n_4303), .A (n_4304));
NAND2_X1 i_4366 (.ZN (n_4302), .A1 (n_4309), .A2 (n_4303));
NAND2_X1 i_4365 (.ZN (n_4301), .A1 (n_4302), .A2 (n_4310));
INV_X1 i_4364 (.ZN (n_4300), .A (n_4419));
NAND2_X1 i_4363 (.ZN (n_4299), .A1 (n_4571), .A2 (n_4574));
NAND2_X1 i_4362 (.ZN (n_4298), .A1 (n_4299), .A2 (n_4300));
NAND3_X1 i_4361 (.ZN (n_4297), .A1 (n_4571), .A2 (n_4419), .A3 (n_4574));
NAND2_X1 i_4360 (.ZN (n_4296), .A1 (n_4298), .A2 (n_4297));
INV_X1 i_4359 (.ZN (n_4295), .A (n_4296));
NAND2_X1 i_4358 (.ZN (n_4294), .A1 (n_4301), .A2 (n_4295));
NAND3_X1 i_4357 (.ZN (n_4293), .A1 (n_4296), .A2 (n_4310), .A3 (n_4302));
NAND3_X1 i_4356 (.ZN (n_4292), .A1 (n_4634), .A2 (n_4633), .A3 (n_4617));
AOI21_X1 i_4355 (.ZN (n_4291), .A (n_4636), .B1 (n_4642), .B2 (n_4664));
INV_X1 i_4354 (.ZN (n_4290), .A (n_4633));
INV_X1 i_4353 (.ZN (n_4289), .A (n_4617));
OAI21_X1 i_4352 (.ZN (n_4288), .A (n_4289), .B1 (n_4290), .B2 (n_4291));
NAND2_X1 i_4351 (.ZN (n_4287), .A1 (n_4288), .A2 (n_4292));
INV_X1 i_4350 (.ZN (n_4286), .A (n_4287));
NAND2_X1 i_4349 (.ZN (n_4285), .A1 (n_4286), .A2 (n_4293));
NAND2_X1 i_4348 (.ZN (n_4284), .A1 (n_4285), .A2 (n_4294));
OAI21_X2 i_4347 (.ZN (n_4283), .A (n_4413), .B1 (n_4410), .B2 (n_4284));
NAND2_X1 i_4346 (.ZN (n_4282), .A1 (n_4416), .A2 (n_4606));
NAND2_X1 i_4345 (.ZN (n_4281), .A1 (n_4282), .A2 (n_4603));
NAND3_X2 i_4344 (.ZN (n_4280), .A1 (n_6124), .A2 (n_6123), .A3 (n_6097));
INV_X1 i_4343 (.ZN (n_4279), .A (n_4280));
AOI21_X1 i_4342 (.ZN (n_4278), .A (n_6097), .B1 (n_6124), .B2 (n_6123));
NAND2_X1 i_4341 (.ZN (n_4277), .A1 (n_5035), .A2 (n_5028));
NAND2_X1 i_4340 (.ZN (n_4276), .A1 (n_4277), .A2 (n_5032));
OAI21_X2 i_4339 (.ZN (n_4275), .A (n_4276), .B1 (n_4278), .B2 (n_4279));
NAND2_X1 i_4338 (.ZN (n_4274), .A1 (n_6124), .A2 (n_6123));
NAND2_X1 i_4337 (.ZN (n_4273), .A1 (n_4274), .A2 (n_6096));
INV_X1 i_4336 (.ZN (n_4272), .A (n_4276));
NAND3_X1 i_4335 (.ZN (n_4271), .A1 (n_4273), .A2 (n_4272), .A3 (n_4280));
NAND3_X1 i_4334 (.ZN (n_4270), .A1 (n_4281), .A2 (n_4275), .A3 (n_4271));
INV_X1 i_4333 (.ZN (n_4269), .A (n_4603));
AOI21_X1 i_4332 (.ZN (n_4268), .A (n_4269), .B1 (n_4606), .B2 (n_4416));
NAND2_X1 i_4331 (.ZN (n_4267), .A1 (n_4271), .A2 (n_4275));
NAND2_X1 i_4330 (.ZN (n_4266), .A1 (n_4267), .A2 (n_4268));
NAND2_X1 i_4329 (.ZN (n_4265), .A1 (n_4266), .A2 (n_4270));
NAND4_X1 i_4328 (.ZN (n_4264), .A1 (n_5748), .A2 (n_5747), .A3 (n_5743), .A4 (n_5742));
INV_X1 i_4327 (.ZN (n_4263), .A (n_5748));
OAI21_X1 i_4326 (.ZN (n_4262), .A (n_5741), .B1 (n_4263), .B2 (n_5746));
NAND2_X1 i_4325 (.ZN (n_4261), .A1 (n_4615), .A2 (n_5019));
NAND2_X1 i_4324 (.ZN (n_4260), .A1 (n_4261), .A2 (n_5015));
NAND3_X1 i_4323 (.ZN (n_4259), .A1 (n_4260), .A2 (n_4264), .A3 (n_4262));
NAND2_X1 i_4322 (.ZN (n_4258), .A1 (n_4262), .A2 (n_4264));
NAND3_X1 i_4321 (.ZN (n_4257), .A1 (n_4261), .A2 (n_5015), .A3 (n_4258));
NAND3_X1 i_4320 (.ZN (n_4256), .A1 (n_4259), .A2 (n_4265), .A3 (n_4257));
INV_X1 i_4319 (.ZN (n_4255), .A (n_4265));
NAND2_X1 i_4318 (.ZN (n_4254), .A1 (n_4259), .A2 (n_4257));
NAND2_X1 i_4317 (.ZN (n_4253), .A1 (n_4254), .A2 (n_4255));
NAND3_X2 i_4316 (.ZN (n_4252), .A1 (n_4283), .A2 (n_4256), .A3 (n_4253));
INV_X1 i_4315 (.ZN (n_4251), .A (n_4271));
NAND3_X1 i_4314 (.ZN (n_4250), .A1 (n_6382), .A2 (n_6094), .A3 (n_6381));
INV_X1 i_4313 (.ZN (n_4249), .A (n_6094));
NAND2_X1 i_4312 (.ZN (n_4248), .A1 (n_6382), .A2 (n_6381));
NAND2_X1 i_4311 (.ZN (n_4247), .A1 (n_4248), .A2 (n_4249));
NAND2_X1 i_4310 (.ZN (n_4246), .A1 (n_4247), .A2 (n_4250));
OAI211_X2 i_4309 (.ZN (n_4245), .A (n_4275), .B (n_4246), .C1 (n_4268), .C2 (n_4251));
INV_X1 i_4308 (.ZN (n_4244), .A (n_4246));
NAND2_X1 i_4307 (.ZN (n_4243), .A1 (n_4281), .A2 (n_4271));
NAND2_X1 i_4306 (.ZN (n_4242), .A1 (n_4243), .A2 (n_4275));
NAND2_X1 i_4305 (.ZN (n_4241), .A1 (n_4242), .A2 (n_4244));
NAND3_X1 i_4304 (.ZN (n_4240), .A1 (n_5733), .A2 (n_5740), .A3 (n_5994));
INV_X1 i_4303 (.ZN (n_4239), .A (n_5994));
INV_X1 i_4302 (.ZN (n_4238), .A (n_5740));
OAI21_X1 i_4301 (.ZN (n_4237), .A (n_4238), .B1 (n_4239), .B2 (n_5995));
NAND2_X2 i_4300 (.ZN (n_4236), .A1 (n_4237), .A2 (n_4240));
NAND3_X1 i_4299 (.ZN (n_4235), .A1 (n_4241), .A2 (n_4245), .A3 (n_4236));
INV_X1 i_4298 (.ZN (n_4234), .A (n_4245));
AOI21_X1 i_4297 (.ZN (n_4233), .A (n_4246), .B1 (n_4243), .B2 (n_4275));
INV_X1 i_4296 (.ZN (n_4232), .A (n_4236));
OAI21_X2 i_4295 (.ZN (n_4231), .A (n_4232), .B1 (n_4234), .B2 (n_4233));
NAND2_X2 i_4294 (.ZN (n_4230), .A1 (n_4255), .A2 (n_4257));
NAND4_X2 i_4293 (.ZN (n_4229), .A1 (n_4231), .A2 (n_4235), .A3 (n_4259), .A4 (n_4230));
NAND3_X1 i_4292 (.ZN (n_4228), .A1 (n_5727), .A2 (n_5737), .A3 (n_5732));
NAND2_X1 i_4291 (.ZN (n_4227), .A1 (n_5737), .A2 (n_5732));
NAND3_X1 i_4290 (.ZN (n_4226), .A1 (n_4227), .A2 (n_5730), .A3 (n_5728));
NAND2_X1 i_4289 (.ZN (n_4225), .A1 (n_4232), .A2 (n_4245));
NAND2_X1 i_4288 (.ZN (n_4224), .A1 (n_4225), .A2 (n_4241));
INV_X1 i_4287 (.ZN (n_4223), .A (n_4224));
NAND3_X2 i_4286 (.ZN (n_4222), .A1 (n_4223), .A2 (n_4226), .A3 (n_4228));
INV_X1 CLOCK_opt_ipo_c559 (.ZN (CLOCK_opt_ipo_n337), .A (n_2773));
INV_X1 i_4283 (.ZN (n_4219), .A (n_4283));
NAND2_X1 i_4282 (.ZN (n_4218), .A1 (n_4253), .A2 (n_4256));
NAND2_X2 i_4281 (.ZN (n_4217), .A1 (n_4218), .A2 (n_4219));
NAND3_X1 i_4280 (.ZN (n_4216), .A1 (n_4287), .A2 (n_4294), .A3 (n_4293));
NAND2_X1 i_4279 (.ZN (n_4215), .A1 (n_4294), .A2 (n_4293));
NAND2_X1 i_4278 (.ZN (n_4214), .A1 (n_4286), .A2 (n_4215));
NAND2_X1 i_4277 (.ZN (n_4213), .A1 (n_4214), .A2 (n_4216));
NAND4_X1 i_4276 (.ZN (n_4212), .A1 (n_4429), .A2 (n_4428), .A3 (n_4424), .A4 (n_4423));
NAND2_X1 i_4275 (.ZN (n_4211), .A1 (n_4429), .A2 (n_4428));
NAND2_X1 i_4274 (.ZN (n_4210), .A1 (n_4211), .A2 (n_4422));
NAND2_X1 i_4273 (.ZN (n_4209), .A1 (n_4210), .A2 (n_4212));
INV_X1 i_4272 (.ZN (n_4208), .A (n_4209));
OAI22_X1 i_4271 (.ZN (n_4207), .A1 (n_4948), .A2 (n_4938), .B1 (n_4936), .B2 (n_4942));
NAND3_X1 i_4270 (.ZN (n_4206), .A1 (n_4207), .A2 (n_4939), .A3 (n_4870));
INV_X2 i_4269 (.ZN (n_4205), .A (n_4206));
AOI21_X1 i_4268 (.ZN (n_4204), .A (n_4870), .B1 (n_4939), .B2 (n_4207));
NOR2_X1 i_4267 (.ZN (n_4203), .A1 (n_4204), .A2 (n_4205));
INV_X1 i_4266 (.ZN (n_4202), .A (n_4494));
NAND3_X1 i_4265 (.ZN (n_4201), .A1 (n_4202), .A2 (n_4508), .A3 (n_4507));
NAND3_X1 i_4264 (.ZN (n_4200), .A1 (n_4201), .A2 (n_4493), .A3 (n_4477));
INV_X1 i_4263 (.ZN (n_4199), .A (n_4477));
NAND2_X1 i_4262 (.ZN (n_4198), .A1 (n_4201), .A2 (n_4493));
NAND2_X1 i_4261 (.ZN (n_4197), .A1 (n_4198), .A2 (n_4199));
NAND2_X1 i_4260 (.ZN (n_4196), .A1 (n_4197), .A2 (n_4200));
INV_X1 i_4259 (.ZN (n_4195), .A (n_4196));
INV_X1 i_4258 (.ZN (n_4194), .A (n_4481));
OAI21_X1 i_4257 (.ZN (n_4193), .A (n_4478), .B1 (n_4194), .B2 (n_4480));
INV_X1 i_4256 (.ZN (n_4192), .A (n_4480));
INV_X1 i_4255 (.ZN (n_4191), .A (n_4478));
NAND3_X1 i_4254 (.ZN (n_4190), .A1 (n_4192), .A2 (n_4481), .A3 (n_4191));
INV_X1 i_4253 (.ZN (n_4189), .A (n_4711));
OAI21_X1 i_4252 (.ZN (n_4188), .A (n_4704), .B1 (n_4189), .B2 (n_4702));
NAND3_X1 i_4251 (.ZN (n_4187), .A1 (n_4711), .A2 (n_4705), .A3 (n_4703));
NAND2_X1 i_4250 (.ZN (n_4186), .A1 (n_4188), .A2 (n_4187));
NAND2_X1 i_4249 (.ZN (n_4185), .A1 (n_4690), .A2 (n_4687));
NAND2_X1 i_4248 (.ZN (n_4184), .A1 (n_4185), .A2 (n_4688));
NAND3_X1 i_4247 (.ZN (n_4183), .A1 (n_4690), .A2 (n_4689), .A3 (n_4687));
NAND2_X1 i_4246 (.ZN (n_4182), .A1 (n_4184), .A2 (n_4183));
NAND2_X1 i_4245 (.ZN (n_4181), .A1 (n_4182), .A2 (n_4186));
NAND4_X1 i_4244 (.ZN (n_4180), .A1 (n_4184), .A2 (n_4188), .A3 (n_4187), .A4 (n_4183));
INV_X1 i_4243 (.ZN (n_4179), .A (n_4504));
INV_X1 i_4242 (.ZN (n_4178), .A (n_4503));
INV_X1 i_4241 (.ZN (n_4177), .A (n_4502));
OAI21_X1 i_4240 (.ZN (n_4176), .A (n_4178), .B1 (n_4179), .B2 (n_4177));
NAND3_X1 i_4239 (.ZN (n_4175), .A1 (n_4504), .A2 (n_4503), .A3 (n_4502));
NAND2_X1 i_4238 (.ZN (n_4174), .A1 (n_4176), .A2 (n_4175));
NAND2_X1 i_4237 (.ZN (n_4173), .A1 (n_4180), .A2 (n_4174));
NAND2_X1 i_4236 (.ZN (n_4172), .A1 (n_4173), .A2 (n_4181));
NAND3_X1 i_4235 (.ZN (n_4171), .A1 (n_4172), .A2 (n_4193), .A3 (n_4190));
NAND2_X1 i_4234 (.ZN (n_4170), .A1 (n_4190), .A2 (n_4193));
NAND3_X1 i_4233 (.ZN (n_4169), .A1 (n_4170), .A2 (n_4181), .A3 (n_4173));
NAND2_X1 i_4232 (.ZN (n_4168), .A1 (n_4487), .A2 (n_4489));
NAND4_X1 i_4231 (.ZN (n_4167), .A1 (n_4168), .A2 (B_imm[23]), .A3 (A_imm[3]), .A4 (n_4490));
AOI21_X1 i_4230 (.ZN (n_4166), .A (n_4483), .B1 (n_4484), .B2 (n_4167));
INV_X1 i_4229 (.ZN (n_4165), .A (n_4166));
NAND3_X1 i_4228 (.ZN (n_4164), .A1 (n_4484), .A2 (n_4167), .A3 (n_4483));
NAND2_X1 i_4227 (.ZN (n_4163), .A1 (n_4165), .A2 (n_4164));
NAND2_X1 i_4226 (.ZN (n_4162), .A1 (B_imm[9]), .A2 (A_imm[15]));
OAI22_X1 i_4225 (.ZN (n_4161), .A1 (n_8927), .A2 (n_8880), .B1 (n_8909), .B2 (n_7691));
NAND2_X1 i_4224 (.ZN (n_4160), .A1 (A_imm[19]), .A2 (B_imm[4]));
NAND4_X1 i_4223 (.ZN (n_4159), .A1 (A_imm[13]), .A2 (B_imm[17]), .A3 (B_imm[10]), .A4 (A_imm[6]));
NAND2_X1 i_4222 (.ZN (n_4158), .A1 (n_4159), .A2 (n_4160));
NAND2_X1 i_4221 (.ZN (n_4157), .A1 (n_4158), .A2 (n_4161));
NAND2_X1 i_4220 (.ZN (n_4156), .A1 (n_4157), .A2 (n_4162));
NAND2_X1 i_4219 (.ZN (n_4155), .A1 (B_imm[24]), .A2 (A_imm[0]));
NAND4_X1 i_4218 (.ZN (n_4154), .A1 (n_4158), .A2 (B_imm[9]), .A3 (A_imm[15]), .A4 (n_4161));
NAND2_X1 i_4217 (.ZN (n_4153), .A1 (n_4154), .A2 (n_4155));
NAND2_X1 i_4216 (.ZN (n_4152), .A1 (B_imm[22]), .A2 (A_imm[2]));
OAI21_X1 i_4215 (.ZN (n_4151), .A (n_4152), .B1 (n_8829), .B2 (n_8645));
NAND2_X1 i_4214 (.ZN (n_4150), .A1 (B_imm[13]), .A2 (A_imm[11]));
NAND4_X1 i_4213 (.ZN (n_4149), .A1 (B_imm[15]), .A2 (B_imm[22]), .A3 (A_imm[9]), .A4 (A_imm[2]));
NAND2_X1 i_4212 (.ZN (n_4148), .A1 (n_4149), .A2 (n_4150));
NAND4_X1 i_4211 (.ZN (n_4147), .A1 (n_4148), .A2 (n_4156), .A3 (n_4153), .A4 (n_4151));
INV_X1 i_4210 (.ZN (n_4146), .A (n_4147));
NAND2_X1 i_4209 (.ZN (n_4145), .A1 (n_4153), .A2 (n_4156));
NAND2_X1 i_4208 (.ZN (n_4144), .A1 (n_4148), .A2 (n_4151));
NAND2_X1 i_4207 (.ZN (n_4143), .A1 (n_4710), .A2 (n_4707));
XNOR2_X1 i_4206 (.ZN (n_4142), .A (n_4143), .B (n_4708));
INV_X1 i_4205 (.ZN (n_4141), .A (n_4142));
AOI21_X1 i_4204 (.ZN (n_4140), .A (n_4141), .B1 (n_4144), .B2 (n_4145));
OAI21_X1 i_4203 (.ZN (n_4139), .A (n_4163), .B1 (n_4140), .B2 (n_4146));
INV_X1 i_4202 (.ZN (n_4138), .A (n_4164));
NOR2_X1 i_4201 (.ZN (n_4137), .A1 (n_4138), .A2 (n_4166));
NAND2_X1 i_4200 (.ZN (n_4136), .A1 (n_4144), .A2 (n_4145));
NAND2_X1 i_4199 (.ZN (n_4135), .A1 (n_4136), .A2 (n_4142));
NAND3_X1 i_4198 (.ZN (n_4134), .A1 (n_4137), .A2 (n_4135), .A3 (n_4147));
INV_X1 i_4197 (.ZN (n_4133), .A (n_4134));
NAND2_X1 i_4196 (.ZN (n_4132), .A1 (B_imm[16]), .A2 (A_imm[7]));
OAI21_X1 i_4195 (.ZN (n_4131), .A (n_4132), .B1 (n_8906), .B2 (n_4366));
NAND2_X1 i_4194 (.ZN (n_4130), .A1 (A_imm[21]), .A2 (B_imm[2]));
NAND4_X1 i_4193 (.ZN (n_4129), .A1 (A_imm[22]), .A2 (B_imm[16]), .A3 (B_imm[1]), .A4 (A_imm[7]));
NAND2_X1 i_4192 (.ZN (n_4128), .A1 (n_4129), .A2 (n_4130));
AOI22_X1 i_4191 (.ZN (n_4127), .A1 (n_4128), .A2 (n_4131), .B1 (B_imm[23]), .B2 (A_imm[1]));
INV_X1 i_4190 (.ZN (n_4126), .A (n_4127));
NAND4_X1 i_4189 (.ZN (n_4125), .A1 (n_4128), .A2 (B_imm[23]), .A3 (A_imm[1]), .A4 (n_4131));
NAND2_X1 i_4188 (.ZN (n_4124), .A1 (B_imm[21]), .A2 (A_imm[3]));
NAND2_X1 i_4187 (.ZN (n_4123), .A1 (n_4125), .A2 (n_4124));
AOI21_X1 i_4186 (.ZN (n_4122), .A (n_4489), .B1 (n_4490), .B2 (n_4487));
INV_X1 i_4185 (.ZN (n_4121), .A (n_4122));
NAND3_X1 i_4184 (.ZN (n_4120), .A1 (n_4490), .A2 (n_4489), .A3 (n_4487));
NAND2_X1 i_4183 (.ZN (n_4119), .A1 (n_4121), .A2 (n_4120));
NAND3_X1 i_4182 (.ZN (n_4118), .A1 (n_4123), .A2 (n_4119), .A3 (n_4126));
INV_X1 i_4181 (.ZN (n_4117), .A (n_4118));
NAND2_X1 i_4180 (.ZN (n_4116), .A1 (n_4123), .A2 (n_4126));
INV_X1 i_4179 (.ZN (n_4115), .A (n_4119));
NAND2_X1 i_4178 (.ZN (n_4114), .A1 (n_4116), .A2 (n_4115));
NAND2_X1 i_4177 (.ZN (n_4113), .A1 (B_imm[14]), .A2 (A_imm[11]));
INV_X1 i_4176 (.ZN (n_4112), .A (n_4113));
AOI21_X1 i_4175 (.ZN (n_4111), .A (n_4117), .B1 (n_4114), .B2 (n_4112));
OAI21_X1 i_4174 (.ZN (n_4110), .A (n_4139), .B1 (n_4133), .B2 (n_4111));
NAND2_X1 i_4173 (.ZN (n_4109), .A1 (n_4169), .A2 (n_4110));
NAND2_X1 i_4172 (.ZN (n_4108), .A1 (n_4109), .A2 (n_4171));
NAND2_X1 i_4171 (.ZN (n_4107), .A1 (n_4108), .A2 (n_4195));
NAND3_X1 i_4170 (.ZN (n_4106), .A1 (n_4196), .A2 (n_4109), .A3 (n_4171));
NAND3_X1 i_4169 (.ZN (n_4105), .A1 (n_4434), .A2 (n_4461), .A3 (n_4462));
INV_X1 i_4168 (.ZN (n_4104), .A (n_4434));
NAND2_X1 i_4167 (.ZN (n_4103), .A1 (n_4461), .A2 (n_4462));
NAND2_X1 i_4166 (.ZN (n_4102), .A1 (n_4103), .A2 (n_4104));
NAND2_X1 i_4165 (.ZN (n_4101), .A1 (n_4102), .A2 (n_4105));
INV_X1 i_4164 (.ZN (n_4100), .A (n_4101));
NAND2_X1 i_4163 (.ZN (n_4099), .A1 (n_4106), .A2 (n_4100));
NAND2_X1 i_4162 (.ZN (n_4098), .A1 (n_4099), .A2 (n_4107));
NAND2_X1 i_4161 (.ZN (n_4097), .A1 (n_4203), .A2 (n_4098));
INV_X1 i_4160 (.ZN (n_4096), .A (n_4441));
OAI21_X1 i_4159 (.ZN (n_4095), .A (n_4435), .B1 (n_4437), .B2 (n_4096));
XNOR2_X1 i_4158 (.ZN (n_4094), .A (n_4436), .B (n_5781));
NAND3_X1 i_4157 (.ZN (n_4093), .A1 (n_4094), .A2 (n_4441), .A3 (n_4438));
NAND2_X1 i_4156 (.ZN (n_4092), .A1 (n_4095), .A2 (n_4093));
INV_X1 i_4155 (.ZN (n_4091), .A (n_4092));
NAND2_X1 i_4154 (.ZN (n_4090), .A1 (B_imm[20]), .A2 (A_imm[4]));
NAND2_X1 i_4153 (.ZN (n_4089), .A1 (B_imm[6]), .A2 (A_imm[17]));
NAND2_X1 i_4152 (.ZN (n_4088), .A1 (A_imm[18]), .A2 (B_imm[5]));
NAND2_X1 i_4151 (.ZN (n_4087), .A1 (n_4089), .A2 (n_4088));
NAND2_X1 i_4150 (.ZN (n_4086), .A1 (A_imm[16]), .A2 (B_imm[7]));
NAND4_X1 i_4149 (.ZN (n_4085), .A1 (B_imm[6]), .A2 (A_imm[18]), .A3 (B_imm[5]), .A4 (A_imm[17]));
NAND2_X1 i_4148 (.ZN (n_4084), .A1 (n_4085), .A2 (n_4086));
NAND2_X1 i_4147 (.ZN (n_4083), .A1 (n_4084), .A2 (n_4087));
NAND2_X1 i_4146 (.ZN (n_4082), .A1 (n_4083), .A2 (n_4090));
NAND4_X1 i_4145 (.ZN (n_4081), .A1 (n_4084), .A2 (B_imm[20]), .A3 (A_imm[4]), .A4 (n_4087));
INV_X1 i_4144 (.ZN (n_4080), .A (n_4081));
NAND2_X1 i_4143 (.ZN (n_4079), .A1 (B_imm[19]), .A2 (A_imm[5]));
INV_X1 i_4142 (.ZN (n_4078), .A (n_4079));
OAI21_X1 i_4141 (.ZN (n_4077), .A (n_4082), .B1 (n_4080), .B2 (n_4078));
INV_X1 i_4140 (.ZN (n_4076), .A (n_4077));
AOI21_X1 i_4139 (.ZN (n_4075), .A (n_4458), .B1 (n_4459), .B2 (n_4457));
NAND3_X1 i_4138 (.ZN (n_4074), .A1 (n_4459), .A2 (n_4458), .A3 (n_4457));
INV_X1 i_4137 (.ZN (n_4073), .A (n_4074));
NOR2_X1 i_4136 (.ZN (n_4072), .A1 (n_4073), .A2 (n_4075));
INV_X1 i_4135 (.ZN (n_4071), .A (n_4072));
NAND2_X1 i_4134 (.ZN (n_4070), .A1 (n_4076), .A2 (n_4071));
INV_X1 i_4133 (.ZN (n_4069), .A (n_4070));
AOI21_X1 i_4132 (.ZN (n_4068), .A (n_4450), .B1 (n_4451), .B2 (n_4448));
NAND3_X1 i_4131 (.ZN (n_4067), .A1 (n_4451), .A2 (n_4450), .A3 (n_4448));
INV_X1 i_4130 (.ZN (n_4066), .A (n_4067));
NOR2_X1 i_4129 (.ZN (n_4065), .A1 (n_4066), .A2 (n_4068));
AOI21_X1 i_4128 (.ZN (n_4064), .A (n_4065), .B1 (n_4077), .B2 (n_4072));
INV_X1 i_4127 (.ZN (n_4063), .A (n_4453));
INV_X1 i_4126 (.ZN (n_4062), .A (n_4446));
OAI21_X1 i_4125 (.ZN (n_4061), .A (n_4062), .B1 (n_4063), .B2 (n_4455));
NAND3_X1 i_4124 (.ZN (n_4060), .A1 (n_4454), .A2 (n_4453), .A3 (n_4446));
NAND2_X1 i_4123 (.ZN (n_4059), .A1 (n_4060), .A2 (n_4061));
OAI21_X1 i_4122 (.ZN (n_4058), .A (n_4059), .B1 (n_4069), .B2 (n_4064));
NAND2_X1 i_4121 (.ZN (n_4057), .A1 (n_4077), .A2 (n_4072));
INV_X1 i_4120 (.ZN (n_4056), .A (n_4065));
NAND2_X1 i_4119 (.ZN (n_4055), .A1 (n_4057), .A2 (n_4056));
INV_X1 i_4118 (.ZN (n_4054), .A (n_4059));
NAND3_X1 i_4117 (.ZN (n_4053), .A1 (n_4055), .A2 (n_4054), .A3 (n_4070));
INV_X1 i_4116 (.ZN (n_4052), .A (n_4896));
NAND2_X1 i_4115 (.ZN (n_4051), .A1 (n_4904), .A2 (n_4895));
NAND2_X1 i_4114 (.ZN (n_4050), .A1 (n_4051), .A2 (n_4052));
NAND3_X1 i_4113 (.ZN (n_4049), .A1 (n_4904), .A2 (n_4896), .A3 (n_4895));
NAND2_X1 i_4112 (.ZN (n_4048), .A1 (n_4050), .A2 (n_4049));
NAND2_X1 i_4111 (.ZN (n_4047), .A1 (n_4053), .A2 (n_4048));
NAND2_X1 i_4110 (.ZN (n_4046), .A1 (n_4047), .A2 (n_4058));
NAND2_X1 i_4109 (.ZN (n_4045), .A1 (n_4046), .A2 (n_4091));
NAND3_X1 i_4108 (.ZN (n_4044), .A1 (n_4092), .A2 (n_4058), .A3 (n_4047));
NAND2_X1 i_4107 (.ZN (n_4043), .A1 (n_4894), .A2 (n_4904));
NAND2_X1 i_4106 (.ZN (n_4042), .A1 (n_4921), .A2 (n_4893));
XNOR2_X1 i_4105 (.ZN (n_4041), .A (n_4042), .B (n_4043));
INV_X1 i_4104 (.ZN (n_4040), .A (n_4041));
NAND2_X1 i_4103 (.ZN (n_4039), .A1 (n_4040), .A2 (n_4044));
INV_X1 i_4102 (.ZN (n_4038), .A (n_4871));
NAND3_X1 i_4101 (.ZN (n_4037), .A1 (n_4890), .A2 (n_4889), .A3 (n_4038));
INV_X1 i_4100 (.ZN (n_4036), .A (n_4037));
AOI21_X1 i_4099 (.ZN (n_4035), .A (n_4038), .B1 (n_4890), .B2 (n_4889));
OAI211_X1 i_4098 (.ZN (n_4034), .A (n_4039), .B (n_4045), .C1 (n_4036), .C2 (n_4035));
NAND2_X1 i_4097 (.ZN (n_4033), .A1 (n_4039), .A2 (n_4045));
NOR2_X1 i_4096 (.ZN (n_4032), .A1 (n_4036), .A2 (n_4035));
NAND2_X1 i_4095 (.ZN (n_4031), .A1 (n_4033), .A2 (n_4032));
NAND3_X1 i_4094 (.ZN (n_4030), .A1 (n_4758), .A2 (n_4756), .A3 (n_4733));
NAND2_X1 i_4093 (.ZN (n_4029), .A1 (n_4758), .A2 (n_4756));
NAND2_X1 i_4092 (.ZN (n_4028), .A1 (n_4029), .A2 (n_4734));
NAND2_X1 i_4091 (.ZN (n_4027), .A1 (n_4028), .A2 (n_4030));
NAND2_X1 i_4090 (.ZN (n_4026), .A1 (n_4031), .A2 (n_4027));
OAI211_X2 i_4089 (.ZN (n_4025), .A (n_4099), .B (n_4107), .C1 (n_4204), .C2 (n_4205));
NAND3_X2 i_4088 (.ZN (n_4024), .A1 (n_4025), .A2 (n_4034), .A3 (n_4026));
NAND2_X1 i_4087 (.ZN (n_4023), .A1 (n_4024), .A2 (n_4097));
NAND2_X1 i_4086 (.ZN (n_4022), .A1 (n_4023), .A2 (n_4208));
NAND3_X2 i_4085 (.ZN (n_4021), .A1 (n_4024), .A2 (n_4209), .A3 (n_4097));
NAND3_X1 i_4084 (.ZN (n_4020), .A1 (n_4667), .A2 (n_4867), .A3 (n_4866));
INV_X1 i_4083 (.ZN (n_4019), .A (n_4667));
NAND2_X1 i_4082 (.ZN (n_4018), .A1 (n_4867), .A2 (n_4866));
NAND2_X1 i_4081 (.ZN (n_4017), .A1 (n_4018), .A2 (n_4019));
NAND2_X2 i_4080 (.ZN (n_4016), .A1 (n_4017), .A2 (n_4020));
INV_X1 i_4079 (.ZN (n_4015), .A (n_4016));
NAND2_X1 i_4078 (.ZN (n_4014), .A1 (n_4021), .A2 (n_4015));
NAND2_X1 i_4077 (.ZN (n_4013), .A1 (n_4014), .A2 (n_4022));
NAND3_X1 i_4076 (.ZN (n_4012), .A1 (n_4664), .A2 (n_4663), .A3 (n_4644));
AOI21_X1 i_4075 (.ZN (n_4011), .A (n_5010), .B1 (n_4666), .B2 (n_4867));
INV_X1 i_4074 (.ZN (n_4010), .A (n_4663));
OAI21_X1 i_4073 (.ZN (n_4009), .A (n_4643), .B1 (n_4010), .B2 (n_4011));
NAND2_X1 i_4072 (.ZN (n_4008), .A1 (n_4009), .A2 (n_4012));
NAND2_X1 i_4071 (.ZN (n_4007), .A1 (n_4008), .A2 (n_4013));
NAND4_X1 i_4070 (.ZN (n_4006), .A1 (n_4009), .A2 (n_4014), .A3 (n_4022), .A4 (n_4012));
NAND3_X1 i_4069 (.ZN (n_4005), .A1 (n_4310), .A2 (n_4309), .A3 (n_4304));
AOI22_X1 i_4068 (.ZN (n_4004), .A1 (n_4312), .A2 (n_4394), .B1 (n_4403), .B2 (n_4408));
INV_X1 i_4067 (.ZN (n_4003), .A (n_4309));
OAI21_X1 i_4066 (.ZN (n_4002), .A (n_4303), .B1 (n_4003), .B2 (n_4004));
NAND2_X2 i_4065 (.ZN (n_4001), .A1 (n_4002), .A2 (n_4005));
NAND2_X1 i_4064 (.ZN (n_4000), .A1 (n_4001), .A2 (n_4006));
NAND2_X1 i_4063 (.ZN (n_3999), .A1 (n_4000), .A2 (n_4007));
NAND2_X2 i_4062 (.ZN (n_3998), .A1 (n_4213), .A2 (n_3999));
INV_X1 i_4061 (.ZN (n_3997), .A (n_3998));
NAND3_X1 i_4060 (.ZN (n_3996), .A1 (n_4413), .A2 (n_4284), .A3 (n_4411));
AOI21_X1 i_4059 (.ZN (n_3995), .A (n_4412), .B1 (n_4612), .B2 (n_4613));
INV_X1 i_4058 (.ZN (n_3994), .A (n_4284));
OAI21_X2 i_4057 (.ZN (n_3993), .A (n_3994), .B1 (n_4410), .B2 (n_3995));
NAND3_X1 i_4056 (.ZN (n_3992), .A1 (n_3993), .A2 (n_3997), .A3 (n_3996));
NAND2_X1 i_4055 (.ZN (n_3991), .A1 (n_4217), .A2 (n_3992));
NAND3_X2 i_4054 (.ZN (n_3990), .A1 (n_3991), .A2 (n_4252), .A3 (n_4221));
INV_X1 i_4053 (.ZN (n_3989), .A (n_4222));
NAND2_X1 i_4052 (.ZN (n_3988), .A1 (n_4231), .A2 (n_4235));
NAND2_X1 i_4051 (.ZN (n_3987), .A1 (n_4230), .A2 (n_4259));
NAND2_X1 i_4050 (.ZN (n_3986), .A1 (n_3988), .A2 (n_3987));
NAND2_X1 i_4049 (.ZN (n_3985), .A1 (n_4226), .A2 (n_4228));
NAND2_X1 i_4048 (.ZN (n_3984), .A1 (n_3985), .A2 (n_4224));
OAI21_X1 i_4047 (.ZN (n_3983), .A (n_3984), .B1 (n_3986), .B2 (n_3989));
INV_X1 i_4046 (.ZN (n_3982), .A (n_3983));
NAND2_X2 i_4045 (.ZN (n_3981), .A1 (n_3990), .A2 (n_3982));
NAND2_X1 i_4044 (.ZN (n_3980), .A1 (n_3981), .A2 (n_5109));
NAND3_X1 i_4043 (.ZN (n_3979), .A1 (n_4110), .A2 (n_4171), .A3 (n_4169));
INV_X1 i_4042 (.ZN (n_3978), .A (n_4110));
NAND2_X1 i_4041 (.ZN (n_3977), .A1 (n_4169), .A2 (n_4171));
NAND2_X1 i_4040 (.ZN (n_3976), .A1 (n_3977), .A2 (n_3978));
NAND2_X1 i_4039 (.ZN (n_3975), .A1 (n_3976), .A2 (n_3979));
AOI21_X1 i_4038 (.ZN (n_3974), .A (n_4763), .B1 (n_4770), .B2 (n_4767));
NAND3_X1 i_4037 (.ZN (n_3973), .A1 (n_4767), .A2 (n_4770), .A3 (n_4763));
INV_X1 i_4036 (.ZN (n_3972), .A (n_3973));
NOR2_X1 i_4035 (.ZN (n_3971), .A1 (n_3972), .A2 (n_3974));
INV_X1 i_4034 (.ZN (n_3970), .A (n_3971));
NAND2_X1 i_4033 (.ZN (n_3969), .A1 (B_imm[14]), .A2 (A_imm[10]));
NAND2_X1 i_4032 (.ZN (n_3968), .A1 (B_imm[15]), .A2 (A_imm[8]));
NAND2_X1 i_4031 (.ZN (n_3967), .A1 (A_imm[21]), .A2 (B_imm[1]));
OAI21_X2 i_4030 (.ZN (n_3966), .A (n_3967), .B1 (n_8956), .B2 (n_6577));
NAND2_X1 i_4029 (.ZN (n_3965), .A1 (A_imm[12]), .A2 (B_imm[10]));
INV_X1 i_4028 (.ZN (n_3964), .A (n_3965));
NAND4_X1 i_4027 (.ZN (n_3963), .A1 (A_imm[18]), .A2 (A_imm[21]), .A3 (B_imm[4]), .A4 (B_imm[1]));
INV_X1 i_4026 (.ZN (n_3962), .A (n_3963));
OAI21_X1 i_4025 (.ZN (n_3961), .A (n_3966), .B1 (n_3962), .B2 (n_3964));
NAND2_X1 i_4024 (.ZN (n_3960), .A1 (n_3961), .A2 (n_3968));
NAND2_X1 i_4023 (.ZN (n_3959), .A1 (B_imm[13]), .A2 (A_imm[10]));
OAI21_X1 i_4022 (.ZN (n_3958), .A (n_3959), .B1 (n_3961), .B2 (n_3968));
NAND2_X1 i_4021 (.ZN (n_3957), .A1 (n_3958), .A2 (n_3960));
NAND2_X1 i_4020 (.ZN (n_3956), .A1 (n_3957), .A2 (n_3969));
NAND4_X1 i_4019 (.ZN (n_3955), .A1 (n_3958), .A2 (B_imm[14]), .A3 (A_imm[10]), .A4 (n_3960));
INV_X1 i_4018 (.ZN (n_3954), .A (n_3955));
INV_X1 i_4017 (.ZN (n_3953), .A (n_4778));
OAI21_X1 i_4016 (.ZN (n_3952), .A (n_4776), .B1 (n_3953), .B2 (n_4774));
NAND3_X1 i_4015 (.ZN (n_3951), .A1 (n_4778), .A2 (n_4777), .A3 (n_4775));
NAND2_X1 i_4014 (.ZN (n_3950), .A1 (n_3952), .A2 (n_3951));
OAI21_X1 i_4013 (.ZN (n_3949), .A (n_3956), .B1 (n_3954), .B2 (n_3950));
NAND2_X1 i_4012 (.ZN (n_3948), .A1 (B_imm[21]), .A2 (A_imm[2]));
NAND2_X1 i_4011 (.ZN (n_3947), .A1 (A_imm[17]), .A2 (B_imm[5]));
NAND2_X1 i_4010 (.ZN (n_3946), .A1 (B_imm[16]), .A2 (A_imm[6]));
NAND2_X1 i_4009 (.ZN (n_3945), .A1 (n_3946), .A2 (n_3947));
NAND2_X1 i_4008 (.ZN (n_3944), .A1 (A_imm[22]), .A2 (B_imm[0]));
INV_X1 i_4007 (.ZN (n_3943), .A (n_3944));
NAND4_X1 i_4006 (.ZN (n_3942), .A1 (B_imm[16]), .A2 (A_imm[17]), .A3 (B_imm[5]), .A4 (A_imm[6]));
INV_X1 i_4005 (.ZN (n_3941), .A (n_3942));
OAI21_X1 i_4004 (.ZN (n_3940), .A (n_3945), .B1 (n_3941), .B2 (n_3943));
NAND2_X1 i_4003 (.ZN (n_3939), .A1 (n_3940), .A2 (n_3948));
NAND2_X1 i_4002 (.ZN (n_3938), .A1 (B_imm[22]), .A2 (A_imm[1]));
OAI21_X1 i_4001 (.ZN (n_3937), .A (n_3938), .B1 (n_3940), .B2 (n_3948));
NAND2_X1 i_4000 (.ZN (n_3936), .A1 (n_3937), .A2 (n_3939));
NAND2_X1 i_3999 (.ZN (n_3935), .A1 (B_imm[12]), .A2 (A_imm[11]));
OAI21_X1 i_3998 (.ZN (n_3934), .A (n_3935), .B1 (n_8849), .B2 (n_8752));
AOI22_X1 i_3997 (.ZN (n_3933), .A1 (A_imm[15]), .A2 (B_imm[7]), .B1 (B_imm[17]), .B2 (A_imm[5]));
NAND2_X1 i_3996 (.ZN (n_3932), .A1 (A_imm[19]), .A2 (B_imm[3]));
NAND4_X1 i_3995 (.ZN (n_3931), .A1 (A_imm[15]), .A2 (B_imm[17]), .A3 (B_imm[7]), .A4 (A_imm[5]));
AOI21_X1 i_3994 (.ZN (n_3930), .A (n_3933), .B1 (n_3932), .B2 (n_3931));
NAND4_X1 i_3993 (.ZN (n_3929), .A1 (B_imm[11]), .A2 (B_imm[12]), .A3 (A_imm[12]), .A4 (A_imm[11]));
INV_X1 i_3992 (.ZN (n_3928), .A (n_3929));
OAI21_X1 i_3991 (.ZN (n_3927), .A (n_3934), .B1 (n_3928), .B2 (n_3930));
NAND2_X1 i_3990 (.ZN (n_3926), .A1 (n_3936), .A2 (n_3927));
INV_X1 i_3989 (.ZN (n_3925), .A (n_3927));
NAND3_X1 i_3988 (.ZN (n_3924), .A1 (n_3925), .A2 (n_3937), .A3 (n_3939));
NAND2_X1 i_3987 (.ZN (n_3923), .A1 (n_4797), .A2 (n_4795));
XNOR2_X1 i_3986 (.ZN (n_3922), .A (n_3923), .B (n_4796));
NAND2_X1 i_3985 (.ZN (n_3921), .A1 (n_3924), .A2 (n_3922));
NAND2_X1 i_3984 (.ZN (n_3920), .A1 (n_3921), .A2 (n_3926));
NAND2_X2 i_3983 (.ZN (n_3919), .A1 (n_3949), .A2 (n_3920));
INV_X1 i_3982 (.ZN (n_3918), .A (n_3919));
INV_X1 i_3981 (.ZN (n_3917), .A (n_3949));
INV_X1 i_3980 (.ZN (n_3916), .A (n_3920));
OAI21_X1 i_3979 (.ZN (n_3915), .A (n_4349), .B1 (n_4357), .B2 (n_4360));
NAND3_X1 i_3978 (.ZN (n_3914), .A1 (n_4359), .A2 (n_4358), .A3 (n_4350));
NAND2_X1 i_3977 (.ZN (n_3913), .A1 (n_3915), .A2 (n_3914));
AOI21_X1 i_3976 (.ZN (n_3912), .A (n_3913), .B1 (n_3917), .B2 (n_3916));
OAI21_X1 i_3975 (.ZN (n_3911), .A (n_3970), .B1 (n_3912), .B2 (n_3918));
INV_X1 i_3974 (.ZN (n_3910), .A (n_3913));
OAI21_X1 i_3973 (.ZN (n_3909), .A (n_3910), .B1 (n_3949), .B2 (n_3920));
NAND3_X1 i_3972 (.ZN (n_3908), .A1 (n_3909), .A2 (n_3971), .A3 (n_3919));
NAND2_X1 i_3971 (.ZN (n_3907), .A1 (n_4367), .A2 (n_4368));
XNOR2_X1 i_3970 (.ZN (n_3906), .A (n_3907), .B (n_4347));
INV_X1 i_3969 (.ZN (n_3905), .A (n_3906));
NAND2_X1 i_3968 (.ZN (n_3904), .A1 (n_3905), .A2 (n_3908));
NAND3_X1 i_3967 (.ZN (n_3903), .A1 (n_4336), .A2 (n_4335), .A3 (n_4329));
INV_X1 i_3966 (.ZN (n_3902), .A (n_4329));
NAND2_X1 i_3965 (.ZN (n_3901), .A1 (n_4336), .A2 (n_4335));
NAND2_X1 i_3964 (.ZN (n_3900), .A1 (n_3901), .A2 (n_3902));
NAND4_X1 i_3963 (.ZN (n_3899), .A1 (n_3904), .A2 (n_3911), .A3 (n_3903), .A4 (n_3900));
INV_X1 i_3962 (.ZN (n_3898), .A (n_3908));
OAI21_X1 i_3961 (.ZN (n_3897), .A (n_3911), .B1 (n_3898), .B2 (n_3906));
NAND2_X1 i_3960 (.ZN (n_3896), .A1 (n_3900), .A2 (n_3903));
NAND2_X1 i_3959 (.ZN (n_3895), .A1 (n_3897), .A2 (n_3896));
NAND3_X1 i_3958 (.ZN (n_3894), .A1 (n_3899), .A2 (n_3895), .A3 (n_3975));
INV_X1 i_3957 (.ZN (n_3893), .A (n_3975));
NAND2_X1 i_3956 (.ZN (n_3892), .A1 (n_3899), .A2 (n_3895));
NAND2_X1 i_3955 (.ZN (n_3891), .A1 (n_3892), .A2 (n_3893));
NAND2_X1 i_3954 (.ZN (n_3890), .A1 (n_3891), .A2 (n_3894));
INV_X1 i_3953 (.ZN (n_3889), .A (n_4781));
NAND3_X1 i_3952 (.ZN (n_3888), .A1 (n_3889), .A2 (n_4803), .A3 (n_4801));
NAND3_X1 i_3951 (.ZN (n_3887), .A1 (n_3888), .A2 (n_4780), .A3 (n_4761));
INV_X1 i_3950 (.ZN (n_3886), .A (n_3887));
AOI21_X1 i_3949 (.ZN (n_3885), .A (n_4761), .B1 (n_3888), .B2 (n_4780));
NOR2_X1 i_3948 (.ZN (n_3884), .A1 (n_3886), .A2 (n_3885));
INV_X1 i_3947 (.ZN (n_3883), .A (n_3884));
INV_X1 i_3946 (.ZN (n_3882), .A (n_4822));
NAND2_X1 i_3945 (.ZN (n_3881), .A1 (n_4838), .A2 (n_4837));
NAND2_X1 i_3944 (.ZN (n_3880), .A1 (n_3881), .A2 (n_3882));
NAND3_X1 i_3943 (.ZN (n_3879), .A1 (n_4838), .A2 (n_4837), .A3 (n_4822));
NAND2_X1 i_3942 (.ZN (n_3878), .A1 (n_3880), .A2 (n_3879));
INV_X1 i_3941 (.ZN (n_3877), .A (n_4791));
NAND4_X1 i_3940 (.ZN (n_3876), .A1 (n_4794), .A2 (B_imm[23]), .A3 (A_imm[2]), .A4 (n_4797));
NAND2_X1 i_3939 (.ZN (n_3875), .A1 (n_4792), .A2 (n_3876));
NAND2_X1 i_3938 (.ZN (n_3874), .A1 (n_3875), .A2 (n_3877));
NAND3_X1 i_3937 (.ZN (n_3873), .A1 (n_4792), .A2 (n_4791), .A3 (n_3876));
NAND2_X1 i_3936 (.ZN (n_3872), .A1 (n_3874), .A2 (n_3873));
NAND2_X1 i_3935 (.ZN (n_3871), .A1 (n_4901), .A2 (n_4898));
NAND2_X1 i_3934 (.ZN (n_3870), .A1 (n_3871), .A2 (n_4899));
NAND3_X1 i_3933 (.ZN (n_3869), .A1 (n_4901), .A2 (n_4898), .A3 (n_4900));
NAND2_X1 i_3932 (.ZN (n_3868), .A1 (n_3870), .A2 (n_3869));
NAND2_X1 i_3931 (.ZN (n_3867), .A1 (n_3872), .A2 (n_3868));
INV_X1 i_3930 (.ZN (n_3866), .A (n_4773));
NAND2_X1 i_3929 (.ZN (n_3865), .A1 (n_4779), .A2 (n_4772));
NAND2_X1 i_3928 (.ZN (n_3864), .A1 (n_3865), .A2 (n_3866));
NAND3_X1 i_3927 (.ZN (n_3863), .A1 (n_4779), .A2 (n_4773), .A3 (n_4772));
NAND2_X1 i_3926 (.ZN (n_3862), .A1 (n_3864), .A2 (n_3863));
NAND4_X1 i_3925 (.ZN (n_3861), .A1 (n_3874), .A2 (n_3870), .A3 (n_3873), .A4 (n_3869));
NAND2_X1 i_3924 (.ZN (n_3860), .A1 (n_3861), .A2 (n_3862));
NAND2_X1 i_3923 (.ZN (n_3859), .A1 (n_3860), .A2 (n_3867));
AOI21_X1 i_3922 (.ZN (n_3858), .A (n_4908), .B1 (n_4909), .B2 (n_4907));
NAND3_X1 i_3921 (.ZN (n_3857), .A1 (n_4909), .A2 (n_4908), .A3 (n_4907));
INV_X1 i_3920 (.ZN (n_3856), .A (n_3857));
NAND2_X1 i_3919 (.ZN (n_3855), .A1 (A_imm[20]), .A2 (B_imm[3]));
OAI21_X1 i_3918 (.ZN (n_3854), .A (n_3855), .B1 (n_8947), .B2 (n_8946));
NAND2_X1 i_3917 (.ZN (n_3853), .A1 (A_imm[23]), .A2 (B_imm[0]));
NAND4_X1 i_3916 (.ZN (n_3852), .A1 (B_imm[8]), .A2 (A_imm[20]), .A3 (B_imm[3]), .A4 (A_imm[15]));
NAND2_X1 i_3915 (.ZN (n_3851), .A1 (n_3852), .A2 (n_3853));
INV_X1 i_3914 (.ZN (n_3850), .A (n_4919));
NAND2_X1 i_3913 (.ZN (n_3849), .A1 (n_4920), .A2 (n_4918));
NAND2_X1 i_3912 (.ZN (n_3848), .A1 (n_3849), .A2 (n_3850));
NAND3_X1 i_3911 (.ZN (n_3847), .A1 (n_4920), .A2 (n_4919), .A3 (n_4918));
NAND2_X1 i_3910 (.ZN (n_3846), .A1 (n_3848), .A2 (n_3847));
NAND3_X1 i_3909 (.ZN (n_3845), .A1 (n_3846), .A2 (n_3851), .A3 (n_3854));
INV_X1 i_3908 (.ZN (n_3844), .A (n_3845));
OAI22_X1 i_3907 (.ZN (n_3843), .A1 (n_8347), .A2 (n_8971), .B1 (n_8423), .B2 (n_8293));
NAND2_X1 i_3906 (.ZN (n_3842), .A1 (B_imm[23]), .A2 (A_imm[0]));
NAND4_X1 i_3905 (.ZN (n_3841), .A1 (B_imm[9]), .A2 (B_imm[18]), .A3 (A_imm[14]), .A4 (A_imm[5]));
NAND2_X1 i_3904 (.ZN (n_3840), .A1 (n_3841), .A2 (n_3842));
NAND2_X1 i_3903 (.ZN (n_3839), .A1 (n_3840), .A2 (n_3843));
INV_X1 i_3902 (.ZN (n_3838), .A (n_3839));
NAND2_X1 i_3901 (.ZN (n_3837), .A1 (n_3851), .A2 (n_3854));
INV_X1 i_3900 (.ZN (n_3836), .A (n_3846));
NAND2_X1 i_3899 (.ZN (n_3835), .A1 (n_3837), .A2 (n_3836));
NAND2_X1 i_3898 (.ZN (n_3834), .A1 (n_3838), .A2 (n_3835));
INV_X1 i_3897 (.ZN (n_3833), .A (n_3834));
OAI22_X1 i_3896 (.ZN (n_3832), .A1 (n_3833), .A2 (n_3844), .B1 (n_3858), .B2 (n_3856));
NOR2_X1 i_3895 (.ZN (n_3831), .A1 (n_3856), .A2 (n_3858));
NAND3_X1 i_3894 (.ZN (n_3830), .A1 (n_3831), .A2 (n_3834), .A3 (n_3845));
INV_X1 i_3893 (.ZN (n_3829), .A (n_4914));
NAND2_X1 i_3892 (.ZN (n_3828), .A1 (n_4915), .A2 (n_4913));
XNOR2_X1 i_3891 (.ZN (n_3827), .A (n_3828), .B (n_3829));
NAND2_X1 i_3890 (.ZN (n_3826), .A1 (n_3830), .A2 (n_3827));
NAND2_X1 i_3889 (.ZN (n_3825), .A1 (n_3826), .A2 (n_3832));
NAND2_X1 i_3888 (.ZN (n_3824), .A1 (n_3825), .A2 (n_3859));
NAND4_X1 i_3887 (.ZN (n_3823), .A1 (n_3826), .A2 (n_3860), .A3 (n_3867), .A4 (n_3832));
INV_X1 i_3886 (.ZN (n_3822), .A (n_4785));
OAI21_X1 i_3885 (.ZN (n_3821), .A (n_4782), .B1 (n_4784), .B2 (n_3822));
INV_X1 i_3884 (.ZN (n_3820), .A (n_4784));
INV_X1 i_3883 (.ZN (n_3819), .A (n_4782));
NAND3_X1 i_3882 (.ZN (n_3818), .A1 (n_3820), .A2 (n_4785), .A3 (n_3819));
NAND2_X1 i_3881 (.ZN (n_3817), .A1 (n_3821), .A2 (n_3818));
INV_X1 i_3880 (.ZN (n_3816), .A (n_3817));
NAND2_X1 i_3879 (.ZN (n_3815), .A1 (n_3823), .A2 (n_3816));
AOI21_X1 i_3878 (.ZN (n_3814), .A (n_3878), .B1 (n_3815), .B2 (n_3824));
INV_X1 i_3877 (.ZN (n_3813), .A (n_3814));
INV_X1 i_3876 (.ZN (n_3812), .A (n_3823));
OAI211_X1 i_3875 (.ZN (n_3811), .A (n_3878), .B (n_3824), .C1 (n_3812), .C2 (n_3817));
NAND3_X1 i_3874 (.ZN (n_3810), .A1 (n_3813), .A2 (n_3883), .A3 (n_3811));
INV_X1 i_3873 (.ZN (n_3809), .A (n_3811));
OAI21_X1 i_3872 (.ZN (n_3808), .A (n_3884), .B1 (n_3814), .B2 (n_3809));
NAND2_X1 i_3871 (.ZN (n_3807), .A1 (n_3808), .A2 (n_3810));
NAND3_X1 i_3870 (.ZN (n_3806), .A1 (n_3911), .A2 (n_3908), .A3 (n_3906));
INV_X1 i_3869 (.ZN (n_3805), .A (n_3974));
AOI22_X1 i_3868 (.ZN (n_3804), .A1 (n_3909), .A2 (n_3919), .B1 (n_3805), .B2 (n_3973));
OAI21_X1 i_3867 (.ZN (n_3803), .A (n_3905), .B1 (n_3804), .B2 (n_3898));
INV_X1 i_3866 (.ZN (n_3802), .A (n_3827));
NAND3_X1 i_3865 (.ZN (n_3801), .A1 (n_3832), .A2 (n_3830), .A3 (n_3802));
AOI21_X1 i_3864 (.ZN (n_3800), .A (n_3844), .B1 (n_3838), .B2 (n_3835));
NOR2_X1 i_3863 (.ZN (n_3799), .A1 (n_3800), .A2 (n_3831));
INV_X1 i_3862 (.ZN (n_3798), .A (n_3830));
OAI21_X1 i_3861 (.ZN (n_3797), .A (n_3827), .B1 (n_3799), .B2 (n_3798));
NAND2_X1 i_3860 (.ZN (n_3796), .A1 (n_3797), .A2 (n_3801));
INV_X1 i_3859 (.ZN (n_3795), .A (n_3835));
OAI21_X1 i_3858 (.ZN (n_3794), .A (n_3838), .B1 (n_3795), .B2 (n_3844));
NAND3_X1 i_3857 (.ZN (n_3793), .A1 (n_3835), .A2 (n_3839), .A3 (n_3845));
NAND2_X1 i_3856 (.ZN (n_3792), .A1 (n_3794), .A2 (n_3793));
OAI22_X1 i_3855 (.ZN (n_3791), .A1 (n_8860), .A2 (n_6677), .B1 (n_8973), .B2 (n_8645));
OAI22_X1 i_3854 (.ZN (n_3790), .A1 (n_6817), .A2 (n_8956), .B1 (n_8859), .B2 (n_6740));
NAND2_X1 i_3853 (.ZN (n_3789), .A1 (B_imm[6]), .A2 (A_imm[15]));
NAND4_X1 i_3852 (.ZN (n_3788), .A1 (A_imm[18]), .A2 (A_imm[21]), .A3 (B_imm[3]), .A4 (B_imm[0]));
NAND2_X1 i_3851 (.ZN (n_3787), .A1 (n_3788), .A2 (n_3789));
NAND2_X1 i_3850 (.ZN (n_3786), .A1 (n_3787), .A2 (n_3790));
NAND4_X1 i_3849 (.ZN (n_3785), .A1 (B_imm[20]), .A2 (B_imm[13]), .A3 (A_imm[9]), .A4 (A_imm[2]));
NAND2_X1 i_3848 (.ZN (n_3784), .A1 (n_3785), .A2 (n_3786));
AOI21_X1 i_3847 (.ZN (n_3783), .A (n_3853), .B1 (n_3854), .B2 (n_3852));
NAND3_X1 i_3846 (.ZN (n_3782), .A1 (n_3854), .A2 (n_3853), .A3 (n_3852));
INV_X1 i_3845 (.ZN (n_3781), .A (n_3782));
OAI211_X1 i_3844 (.ZN (n_3780), .A (n_3784), .B (n_3791), .C1 (n_3781), .C2 (n_3783));
NAND2_X1 i_3843 (.ZN (n_3779), .A1 (n_3784), .A2 (n_3791));
NOR2_X1 i_3842 (.ZN (n_3778), .A1 (n_3781), .A2 (n_3783));
NAND2_X1 i_3841 (.ZN (n_3777), .A1 (n_3779), .A2 (n_3778));
NAND2_X1 i_3840 (.ZN (n_3776), .A1 (n_4087), .A2 (n_4085));
XNOR2_X1 i_3839 (.ZN (n_3775), .A (n_3776), .B (n_4086));
INV_X1 i_3838 (.ZN (n_3774), .A (n_3775));
NAND2_X1 i_3837 (.ZN (n_3773), .A1 (n_3777), .A2 (n_3774));
NAND2_X1 i_3836 (.ZN (n_3772), .A1 (n_3773), .A2 (n_3780));
NAND2_X1 i_3835 (.ZN (n_3771), .A1 (n_3772), .A2 (n_3792));
NAND4_X1 i_3834 (.ZN (n_3770), .A1 (n_3773), .A2 (n_3794), .A3 (n_3793), .A4 (n_3780));
NAND3_X1 i_3833 (.ZN (n_3769), .A1 (n_3926), .A2 (n_3924), .A3 (n_3922));
INV_X1 i_3832 (.ZN (n_3768), .A (n_3922));
NAND2_X1 i_3831 (.ZN (n_3767), .A1 (n_3926), .A2 (n_3924));
NAND2_X1 i_3830 (.ZN (n_3766), .A1 (n_3767), .A2 (n_3768));
NAND2_X1 i_3829 (.ZN (n_3765), .A1 (n_3766), .A2 (n_3769));
NAND2_X1 i_3828 (.ZN (n_3764), .A1 (n_3765), .A2 (n_3770));
NAND2_X1 i_3827 (.ZN (n_3763), .A1 (n_3764), .A2 (n_3771));
NAND2_X1 i_3826 (.ZN (n_3762), .A1 (n_3763), .A2 (n_3796));
NAND4_X2 i_3825 (.ZN (n_3761), .A1 (n_3764), .A2 (n_3797), .A3 (n_3801), .A4 (n_3771));
INV_X1 i_3824 (.ZN (n_3760), .A (n_3761));
INV_X1 i_3823 (.ZN (n_3759), .A (n_3862));
NAND3_X1 i_3822 (.ZN (n_3758), .A1 (n_3867), .A2 (n_3861), .A3 (n_3759));
INV_X1 i_3821 (.ZN (n_3757), .A (n_3758));
AOI21_X1 i_3820 (.ZN (n_3756), .A (n_3759), .B1 (n_3867), .B2 (n_3861));
NOR2_X1 i_3819 (.ZN (n_3755), .A1 (n_3757), .A2 (n_3756));
OAI21_X1 i_3818 (.ZN (n_3754), .A (n_3762), .B1 (n_3760), .B2 (n_3755));
NAND3_X2 i_3817 (.ZN (n_3753), .A1 (n_3754), .A2 (n_3806), .A3 (n_3803));
NAND2_X1 i_3816 (.ZN (n_3752), .A1 (n_3803), .A2 (n_3806));
INV_X1 i_3815 (.ZN (n_3751), .A (n_3754));
NAND2_X2 i_3814 (.ZN (n_3750), .A1 (n_3752), .A2 (n_3751));
NAND2_X1 i_3813 (.ZN (n_3749), .A1 (n_3917), .A2 (n_3916));
NAND3_X1 i_3812 (.ZN (n_3748), .A1 (n_3749), .A2 (n_3919), .A3 (n_3910));
NAND2_X1 i_3811 (.ZN (n_3747), .A1 (n_3749), .A2 (n_3919));
NAND2_X1 i_3810 (.ZN (n_3746), .A1 (n_3747), .A2 (n_3913));
NAND2_X1 i_3809 (.ZN (n_3745), .A1 (n_3746), .A2 (n_3748));
INV_X1 i_3808 (.ZN (n_3744), .A (n_3950));
NAND3_X1 i_3807 (.ZN (n_3743), .A1 (n_3956), .A2 (n_3955), .A3 (n_3744));
NAND2_X1 i_3806 (.ZN (n_3742), .A1 (n_3956), .A2 (n_3955));
NAND2_X1 i_3805 (.ZN (n_3741), .A1 (n_3742), .A2 (n_3950));
NAND2_X1 i_3804 (.ZN (n_3740), .A1 (n_3741), .A2 (n_3743));
INV_X1 i_3803 (.ZN (n_3739), .A (n_3934));
OAI21_X1 i_3802 (.ZN (n_3738), .A (n_3930), .B1 (n_3739), .B2 (n_3928));
INV_X1 i_3801 (.ZN (n_3737), .A (n_3930));
NAND3_X1 i_3800 (.ZN (n_3736), .A1 (n_3934), .A2 (n_3737), .A3 (n_3929));
NAND2_X1 i_3799 (.ZN (n_3735), .A1 (n_3738), .A2 (n_3736));
INV_X1 i_3798 (.ZN (n_3734), .A (n_3842));
NAND2_X1 i_3797 (.ZN (n_3733), .A1 (n_3843), .A2 (n_3841));
NAND2_X1 i_3796 (.ZN (n_3732), .A1 (n_3733), .A2 (n_3734));
NAND3_X1 i_3795 (.ZN (n_3731), .A1 (n_3843), .A2 (n_3842), .A3 (n_3841));
NAND2_X1 i_3794 (.ZN (n_3730), .A1 (n_3732), .A2 (n_3731));
NAND2_X1 i_3793 (.ZN (n_3729), .A1 (n_3730), .A2 (n_3735));
NAND2_X1 i_3792 (.ZN (n_3728), .A1 (B_imm[19]), .A2 (A_imm[3]));
OAI22_X1 i_3791 (.ZN (n_3727), .A1 (n_4366), .A2 (n_8893), .B1 (n_8858), .B2 (n_8429));
NAND2_X1 i_3790 (.ZN (n_3726), .A1 (B_imm[8]), .A2 (A_imm[13]));
NAND4_X1 i_3789 (.ZN (n_3725), .A1 (A_imm[20]), .A2 (A_imm[16]), .A3 (B_imm[5]), .A4 (B_imm[1]));
NAND2_X1 i_3788 (.ZN (n_3724), .A1 (n_3725), .A2 (n_3726));
NAND2_X1 i_3787 (.ZN (n_3723), .A1 (n_3724), .A2 (n_3727));
NAND2_X1 i_3786 (.ZN (n_3722), .A1 (n_3723), .A2 (n_3728));
INV_X1 i_3785 (.ZN (n_3721), .A (n_3722));
NAND2_X1 i_3784 (.ZN (n_3720), .A1 (B_imm[12]), .A2 (A_imm[9]));
OAI21_X1 i_3783 (.ZN (n_3719), .A (n_3720), .B1 (n_8849), .B2 (n_8751));
INV_X2 i_3782 (.ZN (n_3718), .A (A_imm[3]));
OAI22_X1 i_3781 (.ZN (n_3717), .A1 (n_8927), .A2 (n_8573), .B1 (n_8909), .B2 (n_3718));
NAND2_X1 i_3780 (.ZN (n_3716), .A1 (A_imm[15]), .A2 (B_imm[5]));
INV_X1 i_3779 (.ZN (n_3715), .A (n_3716));
NAND4_X1 i_3778 (.ZN (n_3714), .A1 (A_imm[13]), .A2 (B_imm[17]), .A3 (B_imm[7]), .A4 (A_imm[3]));
INV_X1 i_3777 (.ZN (n_3713), .A (n_3714));
OAI21_X1 i_3776 (.ZN (n_3712), .A (n_3717), .B1 (n_3713), .B2 (n_3715));
INV_X1 i_3775 (.ZN (n_3711), .A (n_3712));
NAND4_X1 i_3774 (.ZN (n_3710), .A1 (B_imm[11]), .A2 (B_imm[12]), .A3 (A_imm[10]), .A4 (A_imm[9]));
INV_X1 i_3773 (.ZN (n_3709), .A (n_3710));
OAI21_X1 i_3772 (.ZN (n_3708), .A (n_3719), .B1 (n_3711), .B2 (n_3709));
INV_X1 i_3771 (.ZN (n_3707), .A (n_3728));
INV_X1 i_3770 (.ZN (n_3706), .A (n_3723));
NAND2_X1 i_3769 (.ZN (n_3705), .A1 (n_3706), .A2 (n_3707));
AOI21_X1 i_3768 (.ZN (n_3704), .A (n_3721), .B1 (n_3705), .B2 (n_3708));
NAND4_X1 i_3767 (.ZN (n_3703), .A1 (n_3732), .A2 (n_3738), .A3 (n_3736), .A4 (n_3731));
NAND2_X1 i_3766 (.ZN (n_3702), .A1 (n_3703), .A2 (n_3704));
NAND2_X1 i_3765 (.ZN (n_3701), .A1 (n_3702), .A2 (n_3729));
NAND2_X1 i_3764 (.ZN (n_3700), .A1 (n_3740), .A2 (n_3701));
NAND4_X1 i_3763 (.ZN (n_3699), .A1 (n_3741), .A2 (n_3702), .A3 (n_3743), .A4 (n_3729));
NAND2_X1 i_3762 (.ZN (n_3698), .A1 (A_imm[16]), .A2 (B_imm[6]));
OAI21_X1 i_3761 (.ZN (n_3697), .A (n_3698), .B1 (n_8893), .B2 (n_6584));
NAND2_X1 i_3760 (.ZN (n_3696), .A1 (B_imm[8]), .A2 (A_imm[14]));
INV_X1 i_3759 (.ZN (n_3695), .A (n_3696));
NAND4_X1 i_3758 (.ZN (n_3694), .A1 (A_imm[20]), .A2 (A_imm[16]), .A3 (B_imm[6]), .A4 (B_imm[2]));
INV_X1 i_3757 (.ZN (n_3693), .A (n_3694));
OAI21_X1 i_3756 (.ZN (n_3692), .A (n_3697), .B1 (n_3693), .B2 (n_3695));
INV_X1 i_3755 (.ZN (n_3691), .A (n_3692));
OAI22_X1 i_3754 (.ZN (n_3690), .A1 (n_8525), .A2 (n_6678), .B1 (n_8860), .B2 (n_3718));
NAND4_X1 i_3753 (.ZN (n_3689), .A1 (B_imm[19]), .A2 (B_imm[20]), .A3 (A_imm[4]), .A4 (A_imm[3]));
NAND2_X1 i_3752 (.ZN (n_3688), .A1 (n_3690), .A2 (n_3689));
NAND2_X1 i_3751 (.ZN (n_3687), .A1 (n_3688), .A2 (n_3691));
NAND3_X1 i_3750 (.ZN (n_3686), .A1 (n_3690), .A2 (n_3692), .A3 (n_3689));
NAND2_X1 i_3749 (.ZN (n_3685), .A1 (n_3687), .A2 (n_3686));
NAND2_X1 i_3748 (.ZN (n_3684), .A1 (n_3942), .A2 (n_3944));
NAND4_X1 i_3747 (.ZN (n_3683), .A1 (n_3684), .A2 (B_imm[21]), .A3 (A_imm[2]), .A4 (n_3945));
NAND2_X1 i_3746 (.ZN (n_3682), .A1 (n_3939), .A2 (n_3683));
NAND3_X1 i_3745 (.ZN (n_3681), .A1 (n_3682), .A2 (B_imm[22]), .A3 (A_imm[1]));
NAND3_X1 i_3744 (.ZN (n_3680), .A1 (n_3939), .A2 (n_3683), .A3 (n_3938));
NAND2_X1 i_3743 (.ZN (n_3679), .A1 (n_3681), .A2 (n_3680));
NAND2_X1 i_3742 (.ZN (n_3678), .A1 (n_3685), .A2 (n_3679));
NAND4_X1 i_3741 (.ZN (n_3677), .A1 (n_3687), .A2 (n_3680), .A3 (n_3686), .A4 (n_3681));
NAND2_X1 i_3740 (.ZN (n_3676), .A1 (n_3963), .A2 (n_3965));
NAND4_X1 i_3739 (.ZN (n_3675), .A1 (n_3676), .A2 (B_imm[15]), .A3 (A_imm[8]), .A4 (n_3966));
NAND2_X1 i_3738 (.ZN (n_3674), .A1 (n_3960), .A2 (n_3675));
NAND3_X1 i_3737 (.ZN (n_3673), .A1 (n_3674), .A2 (B_imm[13]), .A3 (A_imm[10]));
NAND3_X1 i_3736 (.ZN (n_3672), .A1 (n_3960), .A2 (n_3675), .A3 (n_3959));
NAND2_X1 i_3735 (.ZN (n_3671), .A1 (n_3673), .A2 (n_3672));
NAND2_X1 i_3734 (.ZN (n_3670), .A1 (n_3677), .A2 (n_3671));
NAND2_X1 i_3733 (.ZN (n_3669), .A1 (n_3670), .A2 (n_3678));
NAND2_X1 i_3732 (.ZN (n_3668), .A1 (n_3699), .A2 (n_3669));
NAND2_X1 i_3731 (.ZN (n_3667), .A1 (n_3668), .A2 (n_3700));
NAND2_X1 i_3730 (.ZN (n_3666), .A1 (n_3667), .A2 (n_3745));
NAND4_X1 i_3729 (.ZN (n_3665), .A1 (n_3746), .A2 (n_3668), .A3 (n_3748), .A4 (n_3700));
INV_X1 i_3728 (.ZN (n_3664), .A (n_3665));
AOI22_X1 i_3727 (.ZN (n_3663), .A1 (n_4148), .A2 (n_4151), .B1 (n_4153), .B2 (n_4156));
OAI21_X1 i_3726 (.ZN (n_3662), .A (n_4141), .B1 (n_4146), .B2 (n_3663));
NAND3_X1 i_3725 (.ZN (n_3661), .A1 (n_4136), .A2 (n_4147), .A3 (n_4142));
NAND2_X1 i_3724 (.ZN (n_3660), .A1 (n_3662), .A2 (n_3661));
NAND2_X1 i_3723 (.ZN (n_3659), .A1 (n_3689), .A2 (n_3692));
INV_X1 i_3722 (.ZN (n_3658), .A (n_4363));
NAND2_X1 i_3721 (.ZN (n_3657), .A1 (n_4364), .A2 (n_4362));
NAND2_X1 i_3720 (.ZN (n_3656), .A1 (n_3657), .A2 (n_3658));
NAND3_X1 i_3719 (.ZN (n_3655), .A1 (n_4364), .A2 (n_4363), .A3 (n_4362));
NAND2_X1 i_3718 (.ZN (n_3654), .A1 (n_3656), .A2 (n_3655));
NAND3_X1 i_3717 (.ZN (n_3653), .A1 (n_3654), .A2 (n_3690), .A3 (n_3659));
INV_X1 i_3716 (.ZN (n_3652), .A (n_3653));
NAND2_X1 i_3715 (.ZN (n_3651), .A1 (n_3659), .A2 (n_3690));
AOI21_X1 i_3714 (.ZN (n_3650), .A (n_4363), .B1 (n_4364), .B2 (n_4362));
INV_X1 i_3713 (.ZN (n_3649), .A (n_3655));
NOR2_X1 i_3712 (.ZN (n_3648), .A1 (n_3649), .A2 (n_3650));
INV_X1 i_3711 (.ZN (n_3647), .A (n_4355));
OAI21_X1 i_3710 (.ZN (n_3646), .A (n_4353), .B1 (n_3647), .B2 (n_4351));
NAND3_X1 i_3709 (.ZN (n_3645), .A1 (n_4355), .A2 (n_4354), .A3 (n_4352));
AOI22_X1 i_3708 (.ZN (n_3644), .A1 (n_3651), .A2 (n_3648), .B1 (n_3646), .B2 (n_3645));
NOR2_X1 i_3707 (.ZN (n_3643), .A1 (n_3644), .A2 (n_3652));
NAND2_X1 i_3706 (.ZN (n_3642), .A1 (n_3660), .A2 (n_3643));
NAND2_X1 i_3705 (.ZN (n_3641), .A1 (n_3651), .A2 (n_3648));
INV_X1 i_3704 (.ZN (n_3640), .A (n_3641));
NAND2_X1 i_3703 (.ZN (n_3639), .A1 (n_3646), .A2 (n_3645));
INV_X1 i_3702 (.ZN (n_3638), .A (n_3639));
OAI21_X1 i_3701 (.ZN (n_3637), .A (n_3653), .B1 (n_3640), .B2 (n_3638));
NAND3_X1 i_3700 (.ZN (n_3636), .A1 (n_3637), .A2 (n_3662), .A3 (n_3661));
AOI21_X1 i_3699 (.ZN (n_3635), .A (n_4150), .B1 (n_4151), .B2 (n_4149));
NAND3_X1 i_3698 (.ZN (n_3634), .A1 (n_4151), .A2 (n_4150), .A3 (n_4149));
INV_X1 i_3697 (.ZN (n_3633), .A (n_3634));
NAND2_X1 i_3696 (.ZN (n_3632), .A1 (n_4154), .A2 (n_4156));
NAND3_X1 i_3695 (.ZN (n_3631), .A1 (n_3632), .A2 (B_imm[24]), .A3 (A_imm[0]));
NAND3_X1 i_3694 (.ZN (n_3630), .A1 (n_4156), .A2 (n_4154), .A3 (n_4155));
NAND2_X1 i_3693 (.ZN (n_3629), .A1 (n_3631), .A2 (n_3630));
OAI21_X1 i_3692 (.ZN (n_3628), .A (n_3629), .B1 (n_3635), .B2 (n_3633));
INV_X1 i_3691 (.ZN (n_3627), .A (n_3635));
NAND4_X1 i_3690 (.ZN (n_3626), .A1 (n_3627), .A2 (n_3631), .A3 (n_3634), .A4 (n_3630));
OAI22_X1 i_3689 (.ZN (n_3625), .A1 (n_8880), .A2 (n_8926), .B1 (n_8909), .B2 (n_6678));
NAND2_X1 i_3688 (.ZN (n_3624), .A1 (A_imm[14]), .A2 (B_imm[7]));
NAND4_X1 i_3687 (.ZN (n_3623), .A1 (B_imm[10]), .A2 (A_imm[11]), .A3 (B_imm[17]), .A4 (A_imm[4]));
NAND2_X1 i_3686 (.ZN (n_3622), .A1 (n_3623), .A2 (n_3624));
NAND2_X1 i_3685 (.ZN (n_3621), .A1 (n_3622), .A2 (n_3625));
OAI21_X1 i_3684 (.ZN (n_3620), .A (n_3621), .B1 (n_8795), .B2 (n_8751));
NAND2_X1 i_3683 (.ZN (n_3619), .A1 (B_imm[11]), .A2 (A_imm[11]));
INV_X1 i_3682 (.ZN (n_3618), .A (n_3619));
NAND4_X1 i_3681 (.ZN (n_3617), .A1 (B_imm[12]), .A2 (n_3622), .A3 (A_imm[10]), .A4 (n_3625));
INV_X1 i_3680 (.ZN (n_3616), .A (n_3617));
OAI21_X1 i_3679 (.ZN (n_3615), .A (n_3620), .B1 (n_3616), .B2 (n_3618));
INV_X1 i_3678 (.ZN (n_3614), .A (n_3615));
NAND2_X1 i_3677 (.ZN (n_3613), .A1 (n_4161), .A2 (n_4159));
NAND3_X1 i_3676 (.ZN (n_3612), .A1 (n_3613), .A2 (B_imm[4]), .A3 (A_imm[19]));
NAND3_X1 i_3675 (.ZN (n_3611), .A1 (n_4161), .A2 (n_4160), .A3 (n_4159));
NAND2_X1 i_3674 (.ZN (n_3610), .A1 (n_3612), .A2 (n_3611));
NAND2_X1 i_3673 (.ZN (n_3609), .A1 (n_3614), .A2 (n_3610));
NAND2_X1 i_3672 (.ZN (n_3608), .A1 (B_imm[18]), .A2 (A_imm[4]));
OAI21_X1 i_3671 (.ZN (n_3607), .A (n_3608), .B1 (n_8347), .B2 (n_8927));
NAND2_X1 i_3670 (.ZN (n_3606), .A1 (A_imm[19]), .A2 (B_imm[2]));
OAI21_X1 i_3669 (.ZN (n_3605), .A (n_3606), .B1 (n_8955), .B2 (n_6577));
NAND2_X1 i_3668 (.ZN (n_3604), .A1 (B_imm[16]), .A2 (A_imm[5]));
INV_X1 i_3667 (.ZN (n_3603), .A (n_3604));
NAND4_X1 i_3666 (.ZN (n_3602), .A1 (A_imm[17]), .A2 (A_imm[19]), .A3 (B_imm[4]), .A4 (B_imm[2]));
INV_X1 i_3665 (.ZN (n_3601), .A (n_3602));
OAI21_X1 i_3664 (.ZN (n_3600), .A (n_3605), .B1 (n_3601), .B2 (n_3603));
INV_X1 i_3663 (.ZN (n_3599), .A (n_3600));
NAND4_X1 i_3662 (.ZN (n_3598), .A1 (B_imm[9]), .A2 (B_imm[18]), .A3 (A_imm[13]), .A4 (A_imm[4]));
INV_X1 i_3661 (.ZN (n_3597), .A (n_3598));
OAI21_X1 i_3660 (.ZN (n_3596), .A (n_3607), .B1 (n_3599), .B2 (n_3597));
INV_X1 i_3659 (.ZN (n_3595), .A (n_3596));
NAND3_X1 i_3658 (.ZN (n_3594), .A1 (n_3615), .A2 (n_3612), .A3 (n_3611));
NAND2_X1 i_3657 (.ZN (n_3593), .A1 (n_3594), .A2 (n_3595));
NAND2_X1 i_3656 (.ZN (n_3592), .A1 (n_3593), .A2 (n_3609));
NAND2_X1 i_3655 (.ZN (n_3591), .A1 (n_3592), .A2 (n_3626));
NAND2_X1 i_3654 (.ZN (n_3590), .A1 (n_3591), .A2 (n_3628));
NAND3_X1 i_3653 (.ZN (n_3589), .A1 (n_3642), .A2 (n_3636), .A3 (n_3590));
NAND2_X1 i_3652 (.ZN (n_3588), .A1 (n_3636), .A2 (n_3642));
INV_X1 i_3651 (.ZN (n_3587), .A (n_3590));
NAND2_X1 i_3650 (.ZN (n_3586), .A1 (n_3588), .A2 (n_3587));
NAND2_X1 i_3649 (.ZN (n_3585), .A1 (n_3586), .A2 (n_3589));
OAI21_X2 i_3648 (.ZN (n_3584), .A (n_3666), .B1 (n_3664), .B2 (n_3585));
NAND2_X2 i_3647 (.ZN (n_3583), .A1 (n_3750), .A2 (n_3584));
NAND2_X1 i_3646 (.ZN (n_3582), .A1 (n_3583), .A2 (n_3753));
NAND2_X2 i_3645 (.ZN (n_3581), .A1 (n_3582), .A2 (n_3807));
INV_X1 i_3644 (.ZN (n_3580), .A (n_3807));
NAND3_X2 i_3643 (.ZN (n_3579), .A1 (n_3580), .A2 (n_3583), .A3 (n_3753));
NAND3_X1 i_3642 (.ZN (n_3578), .A1 (n_3581), .A2 (n_3890), .A3 (n_3579));
INV_X1 i_3641 (.ZN (n_3577), .A (n_3578));
AOI21_X1 i_3640 (.ZN (n_3576), .A (n_3890), .B1 (n_3581), .B2 (n_3579));
INV_X1 i_3639 (.ZN (n_3575), .A (n_4048));
NAND2_X1 i_3638 (.ZN (n_3574), .A1 (n_4058), .A2 (n_4053));
NAND2_X1 i_3637 (.ZN (n_3573), .A1 (n_3574), .A2 (n_3575));
NAND3_X1 i_3636 (.ZN (n_3572), .A1 (n_4058), .A2 (n_4053), .A3 (n_4048));
NAND2_X1 i_3635 (.ZN (n_3571), .A1 (n_3573), .A2 (n_3572));
INV_X1 i_3634 (.ZN (n_3570), .A (n_3571));
AOI21_X1 i_3633 (.ZN (n_3569), .A (n_4112), .B1 (n_4114), .B2 (n_4118));
NAND3_X1 i_3632 (.ZN (n_3568), .A1 (n_4114), .A2 (n_4118), .A3 (n_4112));
INV_X1 i_3631 (.ZN (n_3567), .A (n_3568));
NOR2_X1 i_3630 (.ZN (n_3566), .A1 (n_3567), .A2 (n_3569));
AOI22_X1 i_3629 (.ZN (n_3565), .A1 (n_4084), .A2 (n_4087), .B1 (B_imm[20]), .B2 (A_imm[4]));
OAI21_X1 i_3628 (.ZN (n_3564), .A (n_4078), .B1 (n_4080), .B2 (n_3565));
NAND3_X1 i_3627 (.ZN (n_3563), .A1 (n_4082), .A2 (n_4081), .A3 (n_4079));
NAND2_X1 i_3626 (.ZN (n_3562), .A1 (n_3564), .A2 (n_3563));
INV_X1 i_3625 (.ZN (n_3561), .A (n_4125));
INV_X1 i_3624 (.ZN (n_3560), .A (n_4124));
OAI21_X1 i_3623 (.ZN (n_3559), .A (n_3560), .B1 (n_3561), .B2 (n_4127));
NAND3_X1 i_3622 (.ZN (n_3558), .A1 (n_4126), .A2 (n_4125), .A3 (n_4124));
NAND2_X1 i_3621 (.ZN (n_3557), .A1 (n_3559), .A2 (n_3558));
NAND2_X1 i_3620 (.ZN (n_3556), .A1 (n_3562), .A2 (n_3557));
NAND4_X1 i_3619 (.ZN (n_3555), .A1 (n_3564), .A2 (n_3559), .A3 (n_3558), .A4 (n_3563));
INV_X1 i_3618 (.ZN (n_3554), .A (A_imm[0]));
NAND2_X1 i_3617 (.ZN (n_3553), .A1 (B_imm[21]), .A2 (A_imm[1]));
OAI21_X1 i_3616 (.ZN (n_3552), .A (n_3553), .B1 (n_8958), .B2 (n_3554));
NAND2_X1 i_3615 (.ZN (n_3551), .A1 (B_imm[15]), .A2 (A_imm[7]));
NAND4_X1 i_3614 (.ZN (n_3550), .A1 (B_imm[22]), .A2 (B_imm[21]), .A3 (A_imm[1]), .A4 (A_imm[0]));
NAND2_X1 i_3613 (.ZN (n_3549), .A1 (n_3550), .A2 (n_3551));
AOI21_X1 i_3612 (.ZN (n_3548), .A (n_4130), .B1 (n_4131), .B2 (n_4129));
NAND3_X1 i_3611 (.ZN (n_3547), .A1 (n_4131), .A2 (n_4130), .A3 (n_4129));
INV_X1 i_3610 (.ZN (n_3546), .A (n_3547));
OAI211_X1 i_3609 (.ZN (n_3545), .A (n_3549), .B (n_3552), .C1 (n_3548), .C2 (n_3546));
NAND2_X1 i_3608 (.ZN (n_3544), .A1 (B_imm[14]), .A2 (A_imm[9]));
INV_X1 i_3607 (.ZN (n_3543), .A (n_3551));
INV_X1 i_3606 (.ZN (n_3542), .A (n_3550));
OAI21_X1 i_3605 (.ZN (n_3541), .A (n_3552), .B1 (n_3542), .B2 (n_3543));
NOR2_X1 i_3604 (.ZN (n_3540), .A1 (n_3546), .A2 (n_3548));
NAND2_X1 i_3603 (.ZN (n_3539), .A1 (n_3541), .A2 (n_3540));
INV_X1 i_3602 (.ZN (n_3538), .A (n_3539));
OAI21_X1 i_3601 (.ZN (n_3537), .A (n_3545), .B1 (n_3538), .B2 (n_3544));
NAND2_X1 i_3600 (.ZN (n_3536), .A1 (n_3537), .A2 (n_3555));
NAND2_X1 i_3599 (.ZN (n_3535), .A1 (n_3536), .A2 (n_3556));
NAND2_X1 i_3598 (.ZN (n_3534), .A1 (n_3535), .A2 (n_3566));
OAI211_X1 i_3597 (.ZN (n_3533), .A (n_3536), .B (n_3556), .C1 (n_3569), .C2 (n_3567));
AOI21_X1 i_3596 (.ZN (n_3532), .A (n_4056), .B1 (n_4070), .B2 (n_4057));
NAND3_X1 i_3595 (.ZN (n_3531), .A1 (n_4070), .A2 (n_4057), .A3 (n_4056));
INV_X1 i_3594 (.ZN (n_3530), .A (n_3531));
NOR2_X1 i_3593 (.ZN (n_3529), .A1 (n_3530), .A2 (n_3532));
NAND2_X1 i_3592 (.ZN (n_3528), .A1 (n_3533), .A2 (n_3529));
NAND2_X1 i_3591 (.ZN (n_3527), .A1 (n_3528), .A2 (n_3534));
NAND2_X1 i_3590 (.ZN (n_3526), .A1 (n_3527), .A2 (n_3570));
NAND3_X1 i_3589 (.ZN (n_3525), .A1 (n_3571), .A2 (n_3534), .A3 (n_3528));
INV_X1 i_3588 (.ZN (n_3524), .A (n_3525));
NAND3_X1 i_3587 (.ZN (n_3523), .A1 (n_3824), .A2 (n_3823), .A3 (n_3816));
NAND2_X1 i_3586 (.ZN (n_3522), .A1 (n_3823), .A2 (n_3824));
NAND2_X1 i_3585 (.ZN (n_3521), .A1 (n_3522), .A2 (n_3817));
NAND2_X1 i_3584 (.ZN (n_3520), .A1 (n_3521), .A2 (n_3523));
OAI21_X1 i_3583 (.ZN (n_3519), .A (n_3526), .B1 (n_3524), .B2 (n_3520));
NAND3_X1 i_3582 (.ZN (n_3518), .A1 (n_4045), .A2 (n_4044), .A3 (n_4041));
INV_X1 i_3581 (.ZN (n_3517), .A (n_3518));
AOI21_X1 i_3580 (.ZN (n_3516), .A (n_4041), .B1 (n_4045), .B2 (n_4044));
INV_X1 i_3579 (.ZN (n_3515), .A (n_3636));
NAND2_X1 i_3578 (.ZN (n_3514), .A1 (n_4181), .A2 (n_4180));
NAND3_X1 i_3577 (.ZN (n_3513), .A1 (n_3514), .A2 (n_4176), .A3 (n_4175));
NAND3_X1 i_3576 (.ZN (n_3512), .A1 (n_4181), .A2 (n_4180), .A3 (n_4174));
NAND2_X1 i_3575 (.ZN (n_3511), .A1 (n_3513), .A2 (n_3512));
INV_X1 i_3574 (.ZN (n_3510), .A (n_3511));
AOI22_X1 i_3573 (.ZN (n_3509), .A1 (n_3660), .A2 (n_3643), .B1 (n_3591), .B2 (n_3628));
OAI21_X1 i_3572 (.ZN (n_3508), .A (n_3510), .B1 (n_3509), .B2 (n_3515));
NAND2_X1 i_3571 (.ZN (n_3507), .A1 (n_3642), .A2 (n_3590));
NAND3_X1 i_3570 (.ZN (n_3506), .A1 (n_3507), .A2 (n_3636), .A3 (n_3511));
INV_X1 i_3569 (.ZN (n_3505), .A (n_4114));
OAI21_X1 i_3568 (.ZN (n_3504), .A (n_4118), .B1 (n_3505), .B2 (n_4113));
NAND3_X1 i_3567 (.ZN (n_3503), .A1 (n_3504), .A2 (n_4139), .A3 (n_4134));
INV_X1 i_3566 (.ZN (n_3502), .A (n_3503));
AOI21_X1 i_3565 (.ZN (n_3501), .A (n_3504), .B1 (n_4139), .B2 (n_4134));
NOR2_X1 i_3564 (.ZN (n_3500), .A1 (n_3502), .A2 (n_3501));
NAND2_X1 i_3563 (.ZN (n_3499), .A1 (n_3506), .A2 (n_3500));
NAND2_X1 i_3562 (.ZN (n_3498), .A1 (n_3499), .A2 (n_3508));
OAI21_X2 i_3561 (.ZN (n_3497), .A (n_3498), .B1 (n_3517), .B2 (n_3516));
NAND2_X1 i_3560 (.ZN (n_3496), .A1 (n_4045), .A2 (n_4044));
NAND2_X1 i_3559 (.ZN (n_3495), .A1 (n_3496), .A2 (n_4040));
NAND4_X1 i_3558 (.ZN (n_3494), .A1 (n_3495), .A2 (n_3518), .A3 (n_3508), .A4 (n_3499));
NAND3_X1 i_3557 (.ZN (n_3493), .A1 (n_3497), .A2 (n_3519), .A3 (n_3494));
INV_X1 i_3556 (.ZN (n_3492), .A (n_3519));
NAND2_X1 i_3555 (.ZN (n_3491), .A1 (n_3494), .A2 (n_3497));
NAND2_X1 i_3554 (.ZN (n_3490), .A1 (n_3491), .A2 (n_3492));
NAND2_X1 i_3553 (.ZN (n_3489), .A1 (n_3490), .A2 (n_3493));
INV_X1 i_3552 (.ZN (n_3488), .A (n_3489));
NAND3_X1 i_3551 (.ZN (n_3487), .A1 (n_3526), .A2 (n_3525), .A3 (n_3520));
INV_X1 i_3550 (.ZN (n_3486), .A (n_3520));
NAND2_X1 i_3549 (.ZN (n_3485), .A1 (n_3526), .A2 (n_3525));
NAND2_X1 i_3548 (.ZN (n_3484), .A1 (n_3485), .A2 (n_3486));
NAND2_X1 i_3547 (.ZN (n_3483), .A1 (n_3484), .A2 (n_3487));
INV_X1 i_3546 (.ZN (n_3482), .A (n_3501));
NAND2_X1 i_3545 (.ZN (n_3481), .A1 (n_3482), .A2 (n_3503));
NAND3_X1 i_3544 (.ZN (n_3480), .A1 (n_3508), .A2 (n_3506), .A3 (n_3481));
INV_X1 i_3543 (.ZN (n_3479), .A (n_3480));
AOI21_X1 i_3542 (.ZN (n_3478), .A (n_3481), .B1 (n_3508), .B2 (n_3506));
NOR2_X1 i_3541 (.ZN (n_3477), .A1 (n_3479), .A2 (n_3478));
INV_X1 i_3540 (.ZN (n_3476), .A (n_3477));
NAND2_X1 i_3539 (.ZN (n_3475), .A1 (n_3483), .A2 (n_3476));
NAND3_X1 i_3538 (.ZN (n_3474), .A1 (n_3484), .A2 (n_3477), .A3 (n_3487));
INV_X1 i_3537 (.ZN (n_3473), .A (n_3474));
NAND3_X1 i_3536 (.ZN (n_3472), .A1 (n_3534), .A2 (n_3533), .A3 (n_3529));
INV_X1 i_3535 (.ZN (n_3471), .A (n_3529));
NAND2_X1 i_3534 (.ZN (n_3470), .A1 (n_3534), .A2 (n_3533));
NAND2_X1 i_3533 (.ZN (n_3469), .A1 (n_3470), .A2 (n_3471));
NAND3_X1 i_3532 (.ZN (n_3468), .A1 (n_3653), .A2 (n_3641), .A3 (n_3638));
INV_X1 i_3531 (.ZN (n_3467), .A (n_3468));
AOI21_X1 i_3530 (.ZN (n_3466), .A (n_3638), .B1 (n_3641), .B2 (n_3653));
AOI21_X1 i_3529 (.ZN (n_3465), .A (n_3944), .B1 (n_3945), .B2 (n_3942));
NAND3_X1 i_3528 (.ZN (n_3464), .A1 (n_3945), .A2 (n_3942), .A3 (n_3944));
INV_X1 i_3527 (.ZN (n_3463), .A (n_3464));
AOI21_X1 i_3526 (.ZN (n_3462), .A (n_3965), .B1 (n_3966), .B2 (n_3963));
NAND3_X1 i_3525 (.ZN (n_3461), .A1 (n_3966), .A2 (n_3965), .A3 (n_3963));
INV_X1 i_3524 (.ZN (n_3460), .A (n_3461));
OAI22_X1 i_3523 (.ZN (n_3459), .A1 (n_3460), .A2 (n_3462), .B1 (n_3463), .B2 (n_3465));
NAND2_X1 i_3522 (.ZN (n_3458), .A1 (B_imm[14]), .A2 (A_imm[8]));
INV_X1 i_3521 (.ZN (n_3457), .A (n_3465));
INV_X1 i_3520 (.ZN (n_3456), .A (n_3462));
NAND4_X1 i_3519 (.ZN (n_3455), .A1 (n_3456), .A2 (n_3457), .A3 (n_3464), .A4 (n_3461));
INV_X1 i_3518 (.ZN (n_3454), .A (n_3455));
OAI21_X1 i_3517 (.ZN (n_3453), .A (n_3459), .B1 (n_3454), .B2 (n_3458));
NAND2_X1 i_3516 (.ZN (n_3452), .A1 (B_imm[21]), .A2 (A_imm[0]));
OAI21_X1 i_3515 (.ZN (n_3451), .A (n_3452), .B1 (n_8829), .B2 (n_7691));
NAND2_X1 i_3514 (.ZN (n_3450), .A1 (B_imm[13]), .A2 (A_imm[8]));
NAND4_X1 i_3513 (.ZN (n_3449), .A1 (B_imm[15]), .A2 (B_imm[21]), .A3 (A_imm[6]), .A4 (A_imm[0]));
NAND2_X1 i_3512 (.ZN (n_3448), .A1 (n_3449), .A2 (n_3450));
INV_X1 i_3511 (.ZN (n_3447), .A (n_3931));
OAI211_X1 i_3510 (.ZN (n_3446), .A (B_imm[3]), .B (A_imm[19]), .C1 (n_3447), .C2 (n_3933));
INV_X1 i_3509 (.ZN (n_3445), .A (n_3933));
NAND3_X1 i_3508 (.ZN (n_3444), .A1 (n_3445), .A2 (n_3932), .A3 (n_3931));
NAND2_X1 i_3507 (.ZN (n_3443), .A1 (n_3446), .A2 (n_3444));
NAND3_X1 i_3506 (.ZN (n_3442), .A1 (n_3448), .A2 (n_3451), .A3 (n_3443));
NAND2_X1 i_3505 (.ZN (n_3441), .A1 (B_imm[18]), .A2 (A_imm[3]));
NAND2_X1 i_3504 (.ZN (n_3440), .A1 (A_imm[19]), .A2 (B_imm[1]));
OAI21_X1 i_3503 (.ZN (n_3439), .A (n_3440), .B1 (n_8751), .B2 (n_8880));
NAND2_X1 i_3502 (.ZN (n_3438), .A1 (A_imm[17]), .A2 (B_imm[3]));
INV_X1 i_3501 (.ZN (n_3437), .A (n_3438));
NAND4_X1 i_3500 (.ZN (n_3436), .A1 (A_imm[10]), .A2 (A_imm[19]), .A3 (B_imm[10]), .A4 (B_imm[1]));
INV_X1 i_3499 (.ZN (n_3435), .A (n_3436));
OAI21_X1 i_3498 (.ZN (n_3434), .A (n_3439), .B1 (n_3435), .B2 (n_3437));
NAND2_X1 i_3497 (.ZN (n_3433), .A1 (n_3434), .A2 (n_3441));
NAND2_X1 i_3496 (.ZN (n_3432), .A1 (B_imm[9]), .A2 (A_imm[12]));
OAI21_X1 i_3495 (.ZN (n_3431), .A (n_3432), .B1 (n_3434), .B2 (n_3441));
NAND2_X1 i_3494 (.ZN (n_3430), .A1 (n_3431), .A2 (n_3433));
AOI21_X1 i_3493 (.ZN (n_3429), .A (n_3443), .B1 (n_3448), .B2 (n_3451));
OAI21_X1 i_3492 (.ZN (n_3428), .A (n_3442), .B1 (n_3429), .B2 (n_3430));
NAND2_X2 i_3491 (.ZN (n_3427), .A1 (n_3428), .A2 (n_3453));
INV_X1 i_3490 (.ZN (n_3426), .A (n_3427));
INV_X1 i_3489 (.ZN (n_3425), .A (n_3453));
INV_X1 i_3488 (.ZN (n_3424), .A (n_3428));
NAND2_X1 i_3487 (.ZN (n_3423), .A1 (n_3424), .A2 (n_3425));
OAI22_X1 i_3486 (.ZN (n_3422), .A1 (n_6584), .A2 (n_8956), .B1 (n_8908), .B2 (n_6678));
NAND2_X1 i_3485 (.ZN (n_3421), .A1 (B_imm[6]), .A2 (A_imm[14]));
NAND4_X1 i_3484 (.ZN (n_3420), .A1 (A_imm[18]), .A2 (B_imm[16]), .A3 (B_imm[2]), .A4 (A_imm[4]));
NAND2_X1 i_3483 (.ZN (n_3419), .A1 (n_3420), .A2 (n_3421));
NAND2_X1 i_3482 (.ZN (n_3418), .A1 (n_3419), .A2 (n_3422));
OAI21_X1 i_3481 (.ZN (n_3417), .A (n_3418), .B1 (n_8860), .B2 (n_6836));
NAND2_X1 i_3480 (.ZN (n_3416), .A1 (B_imm[19]), .A2 (A_imm[2]));
NAND4_X2 i_3479 (.ZN (n_3415), .A1 (n_3419), .A2 (n_3422), .A3 (B_imm[20]), .A4 (A_imm[1]));
NAND2_X1 i_3478 (.ZN (n_3414), .A1 (n_3415), .A2 (n_3416));
AOI21_X1 i_3477 (.ZN (n_3413), .A (n_3696), .B1 (n_3697), .B2 (n_3694));
NAND3_X1 i_3476 (.ZN (n_3412), .A1 (n_3697), .A2 (n_3696), .A3 (n_3694));
INV_X1 i_3475 (.ZN (n_3411), .A (n_3412));
OAI211_X2 i_3474 (.ZN (n_3410), .A (n_3414), .B (n_3417), .C1 (n_3413), .C2 (n_3411));
NAND2_X1 i_3473 (.ZN (n_3409), .A1 (n_3414), .A2 (n_3417));
NOR2_X1 i_3472 (.ZN (n_3408), .A1 (n_3411), .A2 (n_3413));
NAND2_X2 i_3471 (.ZN (n_3407), .A1 (n_3409), .A2 (n_3408));
INV_X1 i_3470 (.ZN (n_3406), .A (n_3620));
OAI21_X1 i_3469 (.ZN (n_3405), .A (n_3618), .B1 (n_3406), .B2 (n_3616));
NAND3_X1 i_3468 (.ZN (n_3404), .A1 (n_3620), .A2 (n_3619), .A3 (n_3617));
NAND2_X1 i_3467 (.ZN (n_3403), .A1 (n_3405), .A2 (n_3404));
NAND2_X2 i_3466 (.ZN (n_3402), .A1 (n_3407), .A2 (n_3403));
NAND2_X1 i_3465 (.ZN (n_3401), .A1 (n_3402), .A2 (n_3410));
NAND2_X1 i_3464 (.ZN (n_3400), .A1 (n_3423), .A2 (n_3401));
INV_X1 i_3463 (.ZN (n_3399), .A (n_3400));
OAI22_X1 i_3462 (.ZN (n_3398), .A1 (n_3399), .A2 (n_3426), .B1 (n_3467), .B2 (n_3466));
NOR2_X1 i_3461 (.ZN (n_3397), .A1 (n_3467), .A2 (n_3466));
NAND3_X1 i_3460 (.ZN (n_3396), .A1 (n_3397), .A2 (n_3400), .A3 (n_3427));
INV_X1 i_3459 (.ZN (n_3395), .A (n_3396));
NAND3_X1 i_3458 (.ZN (n_3394), .A1 (n_3628), .A2 (n_3626), .A3 (n_3592));
INV_X1 i_3457 (.ZN (n_3393), .A (n_3592));
NAND2_X1 i_3456 (.ZN (n_3392), .A1 (n_3628), .A2 (n_3626));
NAND2_X1 i_3455 (.ZN (n_3391), .A1 (n_3392), .A2 (n_3393));
NAND2_X1 i_3454 (.ZN (n_3390), .A1 (n_3391), .A2 (n_3394));
OAI21_X1 i_3453 (.ZN (n_3389), .A (n_3398), .B1 (n_3395), .B2 (n_3390));
NAND3_X1 i_3452 (.ZN (n_3388), .A1 (n_3389), .A2 (n_3472), .A3 (n_3469));
INV_X1 i_3451 (.ZN (n_3387), .A (n_3388));
NAND2_X1 i_3450 (.ZN (n_3386), .A1 (n_3469), .A2 (n_3472));
INV_X1 i_3449 (.ZN (n_3385), .A (n_3466));
AOI22_X1 i_3448 (.ZN (n_3384), .A1 (n_3400), .A2 (n_3427), .B1 (n_3385), .B2 (n_3468));
INV_X1 i_3447 (.ZN (n_3383), .A (n_3390));
AOI21_X1 i_3446 (.ZN (n_3382), .A (n_3384), .B1 (n_3396), .B2 (n_3383));
NAND2_X1 i_3445 (.ZN (n_3381), .A1 (n_3386), .A2 (n_3382));
INV_X1 i_3444 (.ZN (n_3380), .A (n_3755));
NAND3_X1 i_3443 (.ZN (n_3379), .A1 (n_3762), .A2 (n_3761), .A3 (n_3380));
INV_X1 i_3442 (.ZN (n_3378), .A (n_3379));
AOI21_X1 i_3441 (.ZN (n_3377), .A (n_3380), .B1 (n_3761), .B2 (n_3762));
NOR2_X1 i_3440 (.ZN (n_3376), .A1 (n_3378), .A2 (n_3377));
AOI21_X1 i_3439 (.ZN (n_3375), .A (n_3387), .B1 (n_3381), .B2 (n_3376));
OAI21_X1 i_3438 (.ZN (n_3374), .A (n_3475), .B1 (n_3473), .B2 (n_3375));
NAND2_X1 i_3437 (.ZN (n_3373), .A1 (n_3374), .A2 (n_3488));
INV_X1 i_3436 (.ZN (n_3372), .A (n_3381));
INV_X1 i_3435 (.ZN (n_3371), .A (n_3377));
NAND2_X1 i_3434 (.ZN (n_3370), .A1 (n_3371), .A2 (n_3379));
OAI21_X1 i_3433 (.ZN (n_3369), .A (n_3388), .B1 (n_3372), .B2 (n_3370));
NAND2_X1 i_3432 (.ZN (n_3368), .A1 (n_3474), .A2 (n_3369));
NAND3_X1 i_3431 (.ZN (n_3367), .A1 (n_3489), .A2 (n_3475), .A3 (n_3368));
OAI211_X1 i_3430 (.ZN (n_3366), .A (n_3373), .B (n_3367), .C1 (n_3577), .C2 (n_3576));
INV_X1 i_3429 (.ZN (n_3365), .A (n_3890));
AOI21_X1 i_3428 (.ZN (n_3364), .A (n_3580), .B1 (n_3583), .B2 (n_3753));
INV_X1 i_3427 (.ZN (n_3363), .A (n_3579));
OAI21_X1 i_3426 (.ZN (n_3362), .A (n_3365), .B1 (n_3363), .B2 (n_3364));
NAND2_X1 i_3425 (.ZN (n_3361), .A1 (n_3362), .A2 (n_3578));
INV_X1 i_3424 (.ZN (n_3360), .A (n_3361));
NAND2_X1 i_3423 (.ZN (n_3359), .A1 (n_3373), .A2 (n_3367));
NAND2_X2 i_3422 (.ZN (n_3358), .A1 (n_3360), .A2 (n_3359));
NAND2_X1 i_3421 (.ZN (n_3357), .A1 (n_3358), .A2 (n_3366));
NAND3_X1 i_3420 (.ZN (n_3356), .A1 (n_3750), .A2 (n_3584), .A3 (n_3753));
INV_X1 i_3419 (.ZN (n_3355), .A (n_3584));
NAND2_X1 i_3418 (.ZN (n_3354), .A1 (n_3750), .A2 (n_3753));
NAND2_X1 i_3417 (.ZN (n_3353), .A1 (n_3354), .A2 (n_3355));
NAND2_X1 i_3416 (.ZN (n_3352), .A1 (n_3353), .A2 (n_3356));
INV_X1 i_3415 (.ZN (n_3351), .A (n_3352));
NAND3_X1 i_3414 (.ZN (n_3350), .A1 (n_3423), .A2 (n_3401), .A3 (n_3427));
NOR2_X1 i_3413 (.ZN (n_3349), .A1 (n_3428), .A2 (n_3453));
OAI211_X1 i_3412 (.ZN (n_3348), .A (n_3410), .B (n_3402), .C1 (n_3426), .C2 (n_3349));
AOI21_X1 i_3411 (.ZN (n_3347), .A (n_3712), .B1 (n_3719), .B2 (n_3710));
NAND3_X1 i_3410 (.ZN (n_3346), .A1 (n_3719), .A2 (n_3712), .A3 (n_3710));
INV_X1 i_3409 (.ZN (n_3345), .A (n_3346));
OAI22_X1 i_3408 (.ZN (n_3344), .A1 (n_8525), .A2 (n_6836), .B1 (n_8860), .B2 (n_3554));
NAND2_X1 i_3407 (.ZN (n_3343), .A1 (B_imm[6]), .A2 (A_imm[13]));
OAI21_X1 i_3406 (.ZN (n_3342), .A (n_3343), .B1 (n_8858), .B2 (n_6817));
OAI22_X1 i_3405 (.ZN (n_3341), .A1 (n_8880), .A2 (n_8511), .B1 (n_8909), .B2 (n_6836));
NAND2_X1 i_3404 (.ZN (n_3340), .A1 (B_imm[7]), .A2 (A_imm[11]));
INV_X1 i_3403 (.ZN (n_3339), .A (n_3340));
NAND4_X1 i_3402 (.ZN (n_3338), .A1 (B_imm[10]), .A2 (B_imm[17]), .A3 (A_imm[8]), .A4 (A_imm[1]));
INV_X1 i_3401 (.ZN (n_3337), .A (n_3338));
OAI21_X1 i_3400 (.ZN (n_3336), .A (n_3341), .B1 (n_3337), .B2 (n_3339));
INV_X1 i_3399 (.ZN (n_3335), .A (n_3336));
NAND4_X1 i_3398 (.ZN (n_3334), .A1 (A_imm[16]), .A2 (B_imm[6]), .A3 (B_imm[3]), .A4 (A_imm[13]));
INV_X1 i_3397 (.ZN (n_3333), .A (n_3334));
OAI21_X1 i_3396 (.ZN (n_3332), .A (n_3342), .B1 (n_3335), .B2 (n_3333));
NAND4_X1 i_3395 (.ZN (n_3331), .A1 (B_imm[19]), .A2 (B_imm[20]), .A3 (A_imm[1]), .A4 (A_imm[0]));
NAND2_X1 i_3394 (.ZN (n_3330), .A1 (n_3332), .A2 (n_3331));
OAI211_X2 i_3393 (.ZN (n_3329), .A (n_3344), .B (n_3330), .C1 (n_3345), .C2 (n_3347));
NOR2_X1 i_3392 (.ZN (n_3328), .A1 (n_3345), .A2 (n_3347));
NAND2_X1 i_3391 (.ZN (n_3327), .A1 (n_3330), .A2 (n_3344));
NAND2_X1 i_3390 (.ZN (n_3326), .A1 (n_3328), .A2 (n_3327));
INV_X1 i_3389 (.ZN (n_3325), .A (n_3432));
INV_X1 i_3388 (.ZN (n_3324), .A (n_3441));
INV_X1 i_3387 (.ZN (n_3323), .A (n_3434));
NAND2_X1 i_3386 (.ZN (n_3322), .A1 (n_3323), .A2 (n_3324));
NAND2_X1 i_3385 (.ZN (n_3321), .A1 (n_3322), .A2 (n_3433));
NAND2_X1 i_3384 (.ZN (n_3320), .A1 (n_3321), .A2 (n_3325));
NAND3_X1 i_3383 (.ZN (n_3319), .A1 (n_3322), .A2 (n_3433), .A3 (n_3432));
NAND2_X1 i_3382 (.ZN (n_3318), .A1 (n_3320), .A2 (n_3319));
NAND2_X1 i_3381 (.ZN (n_3317), .A1 (n_3326), .A2 (n_3318));
NAND2_X1 i_3380 (.ZN (n_3316), .A1 (B_imm[14]), .A2 (A_imm[7]));
OAI22_X2 i_3379 (.ZN (n_3315), .A1 (n_4366), .A2 (n_8956), .B1 (n_8908), .B2 (n_3718));
NAND2_X1 i_3378 (.ZN (n_3314), .A1 (A_imm[12]), .A2 (B_imm[7]));
NAND4_X1 i_3377 (.ZN (n_3313), .A1 (A_imm[18]), .A2 (B_imm[16]), .A3 (B_imm[1]), .A4 (A_imm[3]));
NAND2_X1 i_3376 (.ZN (n_3312), .A1 (n_3313), .A2 (n_3314));
NAND2_X1 i_3375 (.ZN (n_3311), .A1 (n_3312), .A2 (n_3315));
OAI21_X1 i_3374 (.ZN (n_3310), .A (n_3311), .B1 (n_8829), .B2 (n_8293));
NAND2_X1 i_3373 (.ZN (n_3309), .A1 (B_imm[13]), .A2 (A_imm[7]));
NAND4_X1 i_3372 (.ZN (n_3308), .A1 (n_3312), .A2 (B_imm[15]), .A3 (A_imm[5]), .A4 (n_3315));
NAND2_X1 i_3371 (.ZN (n_3307), .A1 (n_3308), .A2 (n_3309));
NAND2_X1 i_3370 (.ZN (n_3306), .A1 (n_3307), .A2 (n_3310));
NAND2_X1 i_3369 (.ZN (n_3305), .A1 (n_3306), .A2 (n_3316));
NAND4_X1 i_3368 (.ZN (n_3304), .A1 (n_3307), .A2 (B_imm[14]), .A3 (A_imm[7]), .A4 (n_3310));
INV_X1 i_3367 (.ZN (n_3303), .A (n_3304));
NAND2_X1 i_3366 (.ZN (n_3302), .A1 (n_3727), .A2 (n_3725));
NAND3_X1 i_3365 (.ZN (n_3301), .A1 (n_3302), .A2 (B_imm[8]), .A3 (A_imm[13]));
NAND3_X1 i_3364 (.ZN (n_3300), .A1 (n_3727), .A2 (n_3726), .A3 (n_3725));
NAND2_X1 i_3363 (.ZN (n_3299), .A1 (n_3301), .A2 (n_3300));
OAI21_X1 i_3362 (.ZN (n_3298), .A (n_3305), .B1 (n_3303), .B2 (n_3299));
NAND3_X2 i_3361 (.ZN (n_3297), .A1 (n_3298), .A2 (n_3329), .A3 (n_3317));
NAND2_X1 i_3360 (.ZN (n_3296), .A1 (n_3317), .A2 (n_3329));
INV_X1 i_3359 (.ZN (n_3295), .A (n_3298));
NAND2_X1 i_3358 (.ZN (n_3294), .A1 (n_3296), .A2 (n_3295));
INV_X1 i_3357 (.ZN (n_3293), .A (n_3442));
OAI211_X1 i_3356 (.ZN (n_3292), .A (n_3433), .B (n_3431), .C1 (n_3429), .C2 (n_3293));
INV_X1 i_3355 (.ZN (n_3291), .A (n_3429));
NAND3_X1 i_3354 (.ZN (n_3290), .A1 (n_3291), .A2 (n_3442), .A3 (n_3430));
NAND2_X1 i_3353 (.ZN (n_3289), .A1 (n_3292), .A2 (n_3290));
INV_X1 i_3352 (.ZN (n_3288), .A (n_3289));
NAND2_X1 i_3351 (.ZN (n_3287), .A1 (n_3294), .A2 (n_3288));
NAND4_X2 i_3350 (.ZN (n_3286), .A1 (n_3348), .A2 (n_3287), .A3 (n_3350), .A4 (n_3297));
INV_X1 i_3349 (.ZN (n_3285), .A (n_3286));
NAND2_X1 i_3348 (.ZN (n_3284), .A1 (n_3348), .A2 (n_3350));
NAND2_X1 i_3347 (.ZN (n_3283), .A1 (n_3287), .A2 (n_3297));
INV_X1 i_3346 (.ZN (n_3282), .A (n_3671));
NAND3_X1 i_3345 (.ZN (n_3281), .A1 (n_3678), .A2 (n_3677), .A3 (n_3282));
INV_X1 i_3344 (.ZN (n_3280), .A (n_3281));
AOI21_X1 i_3343 (.ZN (n_3279), .A (n_3282), .B1 (n_3677), .B2 (n_3678));
NOR2_X1 i_3342 (.ZN (n_3278), .A1 (n_3280), .A2 (n_3279));
AOI21_X1 i_3341 (.ZN (n_3277), .A (n_3278), .B1 (n_3283), .B2 (n_3284));
NAND3_X1 i_3340 (.ZN (n_3276), .A1 (n_3777), .A2 (n_3780), .A3 (n_3775));
INV_X1 i_3339 (.ZN (n_3275), .A (n_3276));
AOI21_X1 i_3338 (.ZN (n_3274), .A (n_3775), .B1 (n_3777), .B2 (n_3780));
NAND2_X1 i_3337 (.ZN (n_3273), .A1 (n_3791), .A2 (n_3785));
NAND3_X1 i_3336 (.ZN (n_3272), .A1 (n_3273), .A2 (n_3790), .A3 (n_3787));
NAND3_X1 i_3335 (.ZN (n_3271), .A1 (n_3791), .A2 (n_3786), .A3 (n_3785));
NAND2_X1 i_3334 (.ZN (n_3270), .A1 (n_3272), .A2 (n_3271));
OAI22_X2 i_3333 (.ZN (n_3269), .A1 (n_8892), .A2 (n_6740), .B1 (n_8946), .B2 (n_6577));
NAND2_X1 i_3332 (.ZN (n_3268), .A1 (A_imm[17]), .A2 (B_imm[2]));
NAND4_X1 i_3331 (.ZN (n_3267), .A1 (A_imm[19]), .A2 (B_imm[4]), .A3 (B_imm[0]), .A4 (A_imm[15]));
NAND2_X1 i_3330 (.ZN (n_3266), .A1 (n_3267), .A2 (n_3268));
NAND2_X1 i_3329 (.ZN (n_3265), .A1 (n_3266), .A2 (n_3269));
OAI21_X1 i_3328 (.ZN (n_3264), .A (n_3265), .B1 (n_8423), .B2 (n_6677));
NAND2_X1 i_3327 (.ZN (n_3263), .A1 (B_imm[9]), .A2 (A_imm[11]));
NAND4_X1 i_3326 (.ZN (n_3262), .A1 (n_3266), .A2 (n_3269), .A3 (B_imm[18]), .A4 (A_imm[2]));
NAND2_X1 i_3325 (.ZN (n_3261), .A1 (n_3262), .A2 (n_3263));
INV_X1 i_3324 (.ZN (n_3260), .A (n_3605));
OAI21_X1 i_3323 (.ZN (n_3259), .A (n_3603), .B1 (n_3260), .B2 (n_3601));
NAND3_X1 i_3322 (.ZN (n_3258), .A1 (n_3605), .A2 (n_3604), .A3 (n_3602));
NAND2_X1 i_3321 (.ZN (n_3257), .A1 (n_3259), .A2 (n_3258));
NAND3_X1 i_3320 (.ZN (n_3256), .A1 (n_3261), .A2 (n_3257), .A3 (n_3264));
INV_X1 i_3319 (.ZN (n_3255), .A (n_3256));
NAND2_X1 i_3318 (.ZN (n_3254), .A1 (n_3261), .A2 (n_3264));
INV_X1 i_3317 (.ZN (n_3253), .A (n_3257));
AOI21_X1 i_3316 (.ZN (n_3252), .A (n_3789), .B1 (n_3790), .B2 (n_3788));
NAND3_X1 i_3315 (.ZN (n_3251), .A1 (n_3790), .A2 (n_3789), .A3 (n_3788));
INV_X1 i_3314 (.ZN (n_3250), .A (n_3251));
NOR2_X2 i_3313 (.ZN (n_3249), .A1 (n_3252), .A2 (n_3250));
AOI21_X1 i_3312 (.ZN (n_3248), .A (n_3249), .B1 (n_3254), .B2 (n_3253));
OAI21_X1 i_3311 (.ZN (n_3247), .A (n_3270), .B1 (n_3248), .B2 (n_3255));
NAND2_X1 i_3310 (.ZN (n_3246), .A1 (n_3254), .A2 (n_3253));
INV_X1 i_3309 (.ZN (n_3245), .A (n_3249));
NAND2_X1 i_3308 (.ZN (n_3244), .A1 (n_3246), .A2 (n_3245));
NAND4_X1 i_3307 (.ZN (n_3243), .A1 (n_3244), .A2 (n_3272), .A3 (n_3271), .A4 (n_3256));
INV_X1 i_3306 (.ZN (n_3242), .A (n_3708));
INV_X1 i_3305 (.ZN (n_3241), .A (n_3705));
OAI21_X1 i_3304 (.ZN (n_3240), .A (n_3242), .B1 (n_3721), .B2 (n_3241));
NAND3_X1 i_3303 (.ZN (n_3239), .A1 (n_3705), .A2 (n_3722), .A3 (n_3708));
NAND2_X1 i_3302 (.ZN (n_3238), .A1 (n_3240), .A2 (n_3239));
NAND2_X1 i_3301 (.ZN (n_3237), .A1 (n_3243), .A2 (n_3238));
NAND2_X1 i_3300 (.ZN (n_3236), .A1 (n_3237), .A2 (n_3247));
OAI21_X1 i_3299 (.ZN (n_3235), .A (n_3236), .B1 (n_3275), .B2 (n_3274));
NOR2_X1 i_3298 (.ZN (n_3234), .A1 (n_3275), .A2 (n_3274));
NAND3_X1 i_3297 (.ZN (n_3233), .A1 (n_3237), .A2 (n_3234), .A3 (n_3247));
INV_X1 i_3296 (.ZN (n_3232), .A (n_3233));
OAI21_X1 i_3295 (.ZN (n_3231), .A (n_3722), .B1 (n_3242), .B2 (n_3241));
AOI21_X1 i_3294 (.ZN (n_3230), .A (n_3231), .B1 (n_3703), .B2 (n_3729));
NAND3_X1 i_3293 (.ZN (n_3229), .A1 (n_3729), .A2 (n_3231), .A3 (n_3703));
INV_X1 i_3292 (.ZN (n_3228), .A (n_3229));
NOR2_X1 i_3291 (.ZN (n_3227), .A1 (n_3228), .A2 (n_3230));
OAI21_X2 i_3290 (.ZN (n_3226), .A (n_3235), .B1 (n_3232), .B2 (n_3227));
OAI21_X2 i_3289 (.ZN (n_3225), .A (n_3226), .B1 (n_3277), .B2 (n_3285));
NAND2_X1 i_3288 (.ZN (n_3224), .A1 (n_3284), .A2 (n_3283));
INV_X1 i_3287 (.ZN (n_3223), .A (n_3278));
NAND2_X1 i_3286 (.ZN (n_3222), .A1 (n_3224), .A2 (n_3223));
INV_X1 i_3285 (.ZN (n_3221), .A (n_3226));
NAND3_X2 i_3284 (.ZN (n_3220), .A1 (n_3222), .A2 (n_3286), .A3 (n_3221));
NAND2_X1 i_3283 (.ZN (n_3219), .A1 (n_3700), .A2 (n_3699));
XNOR2_X1 i_3282 (.ZN (n_3218), .A (n_3219), .B (n_3669));
NAND2_X2 i_3281 (.ZN (n_3217), .A1 (n_3220), .A2 (n_3218));
NAND2_X1 i_3280 (.ZN (n_3216), .A1 (n_3217), .A2 (n_3225));
NAND3_X1 i_3279 (.ZN (n_3215), .A1 (n_3537), .A2 (n_3556), .A3 (n_3555));
NAND2_X1 i_3278 (.ZN (n_3214), .A1 (n_3556), .A2 (n_3555));
OAI211_X1 i_3277 (.ZN (n_3213), .A (n_3214), .B (n_3545), .C1 (n_3544), .C2 (n_3538));
NAND2_X1 i_3276 (.ZN (n_3212), .A1 (n_3213), .A2 (n_3215));
INV_X1 i_3275 (.ZN (n_3211), .A (n_3212));
NAND2_X1 i_3274 (.ZN (n_3210), .A1 (n_3594), .A2 (n_3609));
NAND2_X1 i_3273 (.ZN (n_3209), .A1 (n_3210), .A2 (n_3595));
NAND3_X1 i_3272 (.ZN (n_3208), .A1 (n_3609), .A2 (n_3594), .A3 (n_3596));
INV_X1 i_3271 (.ZN (n_3207), .A (n_3607));
OAI21_X1 i_3270 (.ZN (n_3206), .A (n_3599), .B1 (n_3207), .B2 (n_3597));
NAND3_X1 i_3269 (.ZN (n_3205), .A1 (n_3607), .A2 (n_3600), .A3 (n_3598));
NAND2_X1 i_3268 (.ZN (n_3204), .A1 (n_3206), .A2 (n_3205));
OAI22_X1 i_3267 (.ZN (n_3203), .A1 (n_6740), .A2 (n_8893), .B1 (n_8858), .B2 (n_6577));
NAND2_X1 i_3266 (.ZN (n_3202), .A1 (B_imm[8]), .A2 (A_imm[12]));
NAND4_X1 i_3265 (.ZN (n_3201), .A1 (A_imm[20]), .A2 (A_imm[16]), .A3 (B_imm[4]), .A4 (B_imm[0]));
NAND2_X1 i_3264 (.ZN (n_3200), .A1 (n_3201), .A2 (n_3202));
AOI21_X1 i_3263 (.ZN (n_3199), .A (n_3624), .B1 (n_3625), .B2 (n_3623));
NAND3_X1 i_3262 (.ZN (n_3198), .A1 (n_3625), .A2 (n_3624), .A3 (n_3623));
INV_X1 i_3261 (.ZN (n_3197), .A (n_3198));
OAI211_X1 i_3260 (.ZN (n_3196), .A (n_3200), .B (n_3203), .C1 (n_3199), .C2 (n_3197));
OAI22_X2 i_3259 (.ZN (n_3195), .A1 (n_8971), .A2 (n_8429), .B1 (n_8909), .B2 (n_6677));
NAND2_X1 i_3258 (.ZN (n_3194), .A1 (A_imm[9]), .A2 (B_imm[10]));
NAND4_X1 i_3257 (.ZN (n_3193), .A1 (A_imm[14]), .A2 (B_imm[17]), .A3 (B_imm[5]), .A4 (A_imm[2]));
NAND2_X1 i_3256 (.ZN (n_3192), .A1 (n_3193), .A2 (n_3194));
NAND2_X1 i_3255 (.ZN (n_3191), .A1 (n_3192), .A2 (n_3195));
OAI21_X1 i_3254 (.ZN (n_3190), .A (n_3191), .B1 (n_8795), .B2 (n_8511));
NAND2_X1 i_3253 (.ZN (n_3189), .A1 (B_imm[11]), .A2 (A_imm[9]));
INV_X1 i_3252 (.ZN (n_3188), .A (n_3189));
NAND4_X1 i_3251 (.ZN (n_3187), .A1 (n_3192), .A2 (B_imm[12]), .A3 (n_3195), .A4 (A_imm[8]));
INV_X1 i_3250 (.ZN (n_3186), .A (n_3187));
OAI21_X1 i_3249 (.ZN (n_3185), .A (n_3190), .B1 (n_3186), .B2 (n_3188));
NAND2_X1 i_3248 (.ZN (n_3184), .A1 (n_3200), .A2 (n_3203));
NOR2_X1 i_3247 (.ZN (n_3183), .A1 (n_3199), .A2 (n_3197));
NAND2_X1 i_3246 (.ZN (n_3182), .A1 (n_3184), .A2 (n_3183));
INV_X1 i_3245 (.ZN (n_3181), .A (n_3182));
OAI21_X1 i_3244 (.ZN (n_3180), .A (n_3196), .B1 (n_3181), .B2 (n_3185));
NAND2_X1 i_3243 (.ZN (n_3179), .A1 (n_3180), .A2 (n_3204));
INV_X1 i_3242 (.ZN (n_3178), .A (n_3185));
NAND2_X1 i_3241 (.ZN (n_3177), .A1 (n_3178), .A2 (n_3182));
NAND4_X1 i_3240 (.ZN (n_3176), .A1 (n_3177), .A2 (n_3206), .A3 (n_3205), .A4 (n_3196));
INV_X1 i_3239 (.ZN (n_3175), .A (n_3552));
OAI21_X1 i_3238 (.ZN (n_3174), .A (n_3543), .B1 (n_3175), .B2 (n_3542));
NAND3_X1 i_3237 (.ZN (n_3173), .A1 (n_3552), .A2 (n_3551), .A3 (n_3550));
NAND2_X1 i_3236 (.ZN (n_3172), .A1 (n_3174), .A2 (n_3173));
NAND2_X1 i_3235 (.ZN (n_3171), .A1 (n_3176), .A2 (n_3172));
AOI22_X1 i_3234 (.ZN (n_3170), .A1 (n_3171), .A2 (n_3179), .B1 (n_3209), .B2 (n_3208));
INV_X1 i_3233 (.ZN (n_3169), .A (n_3170));
AOI21_X1 i_3232 (.ZN (n_3168), .A (n_3596), .B1 (n_3594), .B2 (n_3609));
INV_X1 i_3231 (.ZN (n_3167), .A (n_3208));
NOR2_X1 i_3230 (.ZN (n_3166), .A1 (n_3167), .A2 (n_3168));
NAND3_X1 i_3229 (.ZN (n_3165), .A1 (n_3166), .A2 (n_3179), .A3 (n_3171));
INV_X1 i_3228 (.ZN (n_3164), .A (n_3544));
NAND2_X1 i_3227 (.ZN (n_3163), .A1 (n_3545), .A2 (n_3539));
XNOR2_X1 i_3226 (.ZN (n_3162), .A (n_3163), .B (n_3164));
NAND2_X1 i_3225 (.ZN (n_3161), .A1 (n_3162), .A2 (n_3165));
NAND2_X1 i_3224 (.ZN (n_3160), .A1 (n_3161), .A2 (n_3169));
NAND2_X1 i_3223 (.ZN (n_3159), .A1 (n_3160), .A2 (n_3211));
NAND3_X1 i_3222 (.ZN (n_3158), .A1 (n_3212), .A2 (n_3169), .A3 (n_3161));
INV_X1 i_3221 (.ZN (n_3157), .A (n_3158));
NAND3_X1 i_3220 (.ZN (n_3156), .A1 (n_3771), .A2 (n_3765), .A3 (n_3770));
NAND2_X1 i_3219 (.ZN (n_3155), .A1 (n_3771), .A2 (n_3770));
NAND3_X1 i_3218 (.ZN (n_3154), .A1 (n_3155), .A2 (n_3769), .A3 (n_3766));
NAND2_X1 i_3217 (.ZN (n_3153), .A1 (n_3154), .A2 (n_3156));
OAI21_X1 i_3216 (.ZN (n_3152), .A (n_3159), .B1 (n_3157), .B2 (n_3153));
NAND2_X1 i_3215 (.ZN (n_3151), .A1 (n_3216), .A2 (n_3152));
INV_X1 i_3214 (.ZN (n_3150), .A (n_3152));
NAND3_X2 i_3213 (.ZN (n_3149), .A1 (n_3217), .A2 (n_3225), .A3 (n_3150));
NAND3_X1 i_3212 (.ZN (n_3148), .A1 (n_3666), .A2 (n_3665), .A3 (n_3585));
NAND2_X1 i_3211 (.ZN (n_3147), .A1 (n_3666), .A2 (n_3665));
NAND3_X1 i_3210 (.ZN (n_3146), .A1 (n_3147), .A2 (n_3589), .A3 (n_3586));
NAND2_X1 i_3209 (.ZN (n_3145), .A1 (n_3146), .A2 (n_3148));
NAND2_X1 i_3208 (.ZN (n_3144), .A1 (n_3149), .A2 (n_3145));
NAND2_X1 i_3207 (.ZN (n_3143), .A1 (n_3144), .A2 (n_3151));
NAND2_X1 i_3206 (.ZN (n_3142), .A1 (n_3143), .A2 (n_3351));
NAND3_X1 i_3205 (.ZN (n_3141), .A1 (n_3144), .A2 (n_3352), .A3 (n_3151));
NAND3_X1 i_3204 (.ZN (n_3140), .A1 (n_3475), .A2 (n_3369), .A3 (n_3474));
NAND2_X1 i_3203 (.ZN (n_3139), .A1 (n_3475), .A2 (n_3474));
NAND2_X1 i_3202 (.ZN (n_3138), .A1 (n_3139), .A2 (n_3375));
NAND3_X1 i_3201 (.ZN (n_3137), .A1 (n_3141), .A2 (n_3140), .A3 (n_3138));
NAND2_X1 i_3200 (.ZN (n_3136), .A1 (n_3137), .A2 (n_3142));
NAND2_X2 i_3199 (.ZN (n_3135), .A1 (n_3357), .A2 (n_3136));
NAND3_X1 i_3198 (.ZN (n_3134), .A1 (n_4326), .A2 (n_4325), .A3 (n_4323));
INV_X1 i_3197 (.ZN (n_3133), .A (n_3134));
AOI21_X1 i_3196 (.ZN (n_3132), .A (n_4323), .B1 (n_4326), .B2 (n_4325));
NAND2_X1 i_3195 (.ZN (n_3131), .A1 (n_3811), .A2 (n_3884));
NAND2_X1 i_3194 (.ZN (n_3130), .A1 (n_3131), .A2 (n_3813));
INV_X1 i_3193 (.ZN (n_3129), .A (n_3130));
OAI21_X2 i_3192 (.ZN (n_3128), .A (n_3129), .B1 (n_3133), .B2 (n_3132));
INV_X1 i_3191 (.ZN (n_3127), .A (n_4323));
NAND2_X1 i_3190 (.ZN (n_3126), .A1 (n_4326), .A2 (n_4325));
NAND2_X1 i_3189 (.ZN (n_3125), .A1 (n_3126), .A2 (n_3127));
NAND3_X1 i_3188 (.ZN (n_3124), .A1 (n_3125), .A2 (n_3130), .A3 (n_3134));
NAND2_X1 i_3187 (.ZN (n_3123), .A1 (n_3895), .A2 (n_3893));
NAND2_X1 i_3186 (.ZN (n_3122), .A1 (n_3123), .A2 (n_3899));
NAND3_X1 i_3185 (.ZN (n_3121), .A1 (n_3128), .A2 (n_3124), .A3 (n_3122));
NAND2_X1 i_3184 (.ZN (n_3120), .A1 (n_3128), .A2 (n_3124));
INV_X1 i_3183 (.ZN (n_3119), .A (n_3122));
NAND2_X1 i_3182 (.ZN (n_3118), .A1 (n_3120), .A2 (n_3119));
NAND2_X1 i_3181 (.ZN (n_3117), .A1 (n_3118), .A2 (n_3121));
NAND2_X1 i_3180 (.ZN (n_3116), .A1 (n_3579), .A2 (n_3890));
NAND3_X1 i_3179 (.ZN (n_3115), .A1 (n_3117), .A2 (n_3581), .A3 (n_3116));
INV_X1 i_3178 (.ZN (n_3114), .A (n_3117));
NAND2_X1 i_3177 (.ZN (n_3113), .A1 (n_3116), .A2 (n_3581));
NAND2_X1 i_3176 (.ZN (n_3112), .A1 (n_3113), .A2 (n_3114));
NAND3_X1 i_3175 (.ZN (n_3111), .A1 (n_4107), .A2 (n_4106), .A3 (n_4101));
INV_X1 i_3174 (.ZN (n_3110), .A (n_3111));
AOI21_X1 i_3173 (.ZN (n_3109), .A (n_4101), .B1 (n_4107), .B2 (n_4106));
NOR2_X1 i_3172 (.ZN (n_3108), .A1 (n_3110), .A2 (n_3109));
NAND2_X1 i_3171 (.ZN (n_3107), .A1 (n_3494), .A2 (n_3519));
NAND3_X2 i_3170 (.ZN (n_3106), .A1 (n_3108), .A2 (n_3107), .A3 (n_3497));
INV_X1 i_3169 (.ZN (n_3105), .A (n_3108));
NAND2_X1 i_3168 (.ZN (n_3104), .A1 (n_3107), .A2 (n_3497));
NAND2_X1 i_3167 (.ZN (n_3103), .A1 (n_3104), .A2 (n_3105));
NAND3_X1 i_3166 (.ZN (n_3102), .A1 (n_4031), .A2 (n_4034), .A3 (n_4027));
INV_X1 i_3165 (.ZN (n_3101), .A (n_4027));
NAND2_X1 i_3164 (.ZN (n_3100), .A1 (n_4034), .A2 (n_4031));
NAND2_X1 i_3163 (.ZN (n_3099), .A1 (n_3100), .A2 (n_3101));
NAND2_X1 i_3162 (.ZN (n_3098), .A1 (n_3099), .A2 (n_3102));
NAND3_X1 i_3161 (.ZN (n_3097), .A1 (n_3103), .A2 (n_3106), .A3 (n_3098));
INV_X1 i_3160 (.ZN (n_3096), .A (n_3097));
AOI21_X1 i_3159 (.ZN (n_3095), .A (n_3098), .B1 (n_3103), .B2 (n_3106));
OAI211_X1 i_3158 (.ZN (n_3094), .A (n_3112), .B (n_3115), .C1 (n_3096), .C2 (n_3095));
NAND2_X1 i_3157 (.ZN (n_3093), .A1 (n_3112), .A2 (n_3115));
INV_X1 i_3156 (.ZN (n_3092), .A (n_3106));
AOI21_X1 i_3155 (.ZN (n_3091), .A (n_3108), .B1 (n_3497), .B2 (n_3107));
INV_X1 i_3154 (.ZN (n_3090), .A (n_3098));
OAI21_X1 i_3153 (.ZN (n_3089), .A (n_3090), .B1 (n_3092), .B2 (n_3091));
NAND2_X1 i_3152 (.ZN (n_3088), .A1 (n_3089), .A2 (n_3097));
INV_X1 i_3151 (.ZN (n_3087), .A (n_3088));
NAND2_X1 i_3150 (.ZN (n_3086), .A1 (n_3087), .A2 (n_3093));
NAND2_X1 i_3149 (.ZN (n_3085), .A1 (n_3086), .A2 (n_3094));
NAND3_X1 i_3148 (.ZN (n_3084), .A1 (n_3367), .A2 (n_3362), .A3 (n_3578));
NAND2_X1 i_3147 (.ZN (n_3083), .A1 (n_3084), .A2 (n_3373));
NAND2_X2 i_3146 (.ZN (n_3082), .A1 (n_3085), .A2 (n_3083));
INV_X2 i_3145 (.ZN (n_3081), .A (n_3082));
INV_X1 i_3144 (.ZN (n_3080), .A (n_3083));
NAND3_X1 i_3143 (.ZN (n_3079), .A1 (n_3086), .A2 (n_3094), .A3 (n_3080));
INV_X1 i_3142 (.ZN (n_3078), .A (n_3079));
OAI21_X4 i_3141 (.ZN (n_3077), .A (n_3135), .B1 (n_3081), .B2 (n_3078));
NAND2_X1 i_3140 (.ZN (n_3076), .A1 (n_3138), .A2 (n_3140));
NAND3_X1 i_3139 (.ZN (n_3075), .A1 (n_3076), .A2 (n_3142), .A3 (n_3141));
INV_X1 i_3138 (.ZN (n_3074), .A (n_3076));
NAND2_X1 i_3137 (.ZN (n_3073), .A1 (n_3142), .A2 (n_3141));
NAND2_X1 i_3136 (.ZN (n_3072), .A1 (n_3073), .A2 (n_3074));
NAND3_X1 i_3135 (.ZN (n_3071), .A1 (n_3370), .A2 (n_3388), .A3 (n_3381));
OAI21_X1 i_3134 (.ZN (n_3070), .A (n_3376), .B1 (n_3372), .B2 (n_3387));
NAND2_X1 i_3133 (.ZN (n_3069), .A1 (n_3070), .A2 (n_3071));
NAND3_X1 i_3132 (.ZN (n_3068), .A1 (n_3398), .A2 (n_3396), .A3 (n_3390));
OAI21_X2 i_3131 (.ZN (n_3067), .A (n_3383), .B1 (n_3395), .B2 (n_3384));
NAND2_X2 i_3130 (.ZN (n_3066), .A1 (n_3067), .A2 (n_3068));
NAND3_X1 i_3129 (.ZN (n_3065), .A1 (n_3169), .A2 (n_3162), .A3 (n_3165));
INV_X1 i_3128 (.ZN (n_3064), .A (n_3165));
INV_X1 i_3127 (.ZN (n_3063), .A (n_3162));
OAI21_X1 i_3126 (.ZN (n_3062), .A (n_3063), .B1 (n_3064), .B2 (n_3170));
NAND2_X1 i_3125 (.ZN (n_3061), .A1 (n_3459), .A2 (n_3455));
NAND3_X1 i_3124 (.ZN (n_3060), .A1 (n_3061), .A2 (B_imm[14]), .A3 (A_imm[8]));
NAND3_X1 i_3123 (.ZN (n_3059), .A1 (n_3455), .A2 (n_3459), .A3 (n_3458));
NAND2_X1 i_3122 (.ZN (n_3058), .A1 (n_3060), .A2 (n_3059));
NAND2_X1 i_3121 (.ZN (n_3057), .A1 (n_3451), .A2 (n_3449));
NAND3_X1 i_3120 (.ZN (n_3056), .A1 (n_3057), .A2 (B_imm[13]), .A3 (A_imm[8]));
NAND3_X1 i_3119 (.ZN (n_3055), .A1 (n_3451), .A2 (n_3450), .A3 (n_3449));
NAND2_X1 i_3118 (.ZN (n_3054), .A1 (n_3056), .A2 (n_3055));
OAI22_X1 i_3117 (.ZN (n_3053), .A1 (n_8795), .A2 (n_8644), .B1 (n_8947), .B2 (n_8926));
NAND2_X1 i_3116 (.ZN (n_3052), .A1 (B_imm[11]), .A2 (A_imm[8]));
NAND4_X1 i_3115 (.ZN (n_3051), .A1 (B_imm[12]), .A2 (B_imm[8]), .A3 (A_imm[11]), .A4 (A_imm[7]));
NAND2_X1 i_3114 (.ZN (n_3050), .A1 (n_3051), .A2 (n_3052));
NAND2_X1 i_3113 (.ZN (n_3049), .A1 (n_3717), .A2 (n_3714));
NAND2_X1 i_3112 (.ZN (n_3048), .A1 (n_3049), .A2 (n_3715));
NAND3_X1 i_3111 (.ZN (n_3047), .A1 (n_3717), .A2 (n_3716), .A3 (n_3714));
NAND2_X1 i_3110 (.ZN (n_3046), .A1 (n_3048), .A2 (n_3047));
NAND3_X1 i_3109 (.ZN (n_3045), .A1 (n_3046), .A2 (n_3053), .A3 (n_3050));
OAI22_X1 i_3108 (.ZN (n_3044), .A1 (n_8927), .A2 (n_8429), .B1 (n_8971), .B2 (n_6577));
NAND2_X1 i_3107 (.ZN (n_3043), .A1 (A_imm[15]), .A2 (B_imm[3]));
NAND4_X1 i_3106 (.ZN (n_3042), .A1 (A_imm[13]), .A2 (B_imm[5]), .A3 (B_imm[4]), .A4 (A_imm[14]));
NAND2_X1 i_3105 (.ZN (n_3041), .A1 (n_3042), .A2 (n_3043));
NAND2_X1 i_3104 (.ZN (n_3040), .A1 (n_3041), .A2 (n_3044));
OAI21_X1 i_3103 (.ZN (n_3039), .A (n_3040), .B1 (n_8423), .B2 (n_6836));
NAND2_X1 i_3102 (.ZN (n_3038), .A1 (B_imm[9]), .A2 (A_imm[10]));
INV_X1 i_3101 (.ZN (n_3037), .A (n_3038));
NAND4_X1 i_3100 (.ZN (n_3036), .A1 (n_3041), .A2 (n_3044), .A3 (B_imm[18]), .A4 (A_imm[1]));
INV_X1 i_3099 (.ZN (n_3035), .A (n_3036));
OAI21_X2 i_3098 (.ZN (n_3034), .A (n_3039), .B1 (n_3035), .B2 (n_3037));
INV_X1 i_3097 (.ZN (n_3033), .A (n_3034));
NAND2_X1 i_3096 (.ZN (n_3032), .A1 (n_3050), .A2 (n_3053));
NAND3_X1 i_3095 (.ZN (n_3031), .A1 (n_3032), .A2 (n_3048), .A3 (n_3047));
NAND2_X2 i_3094 (.ZN (n_3030), .A1 (n_3031), .A2 (n_3033));
NAND2_X2 i_3093 (.ZN (n_3029), .A1 (n_3030), .A2 (n_3045));
NAND2_X1 i_3092 (.ZN (n_3028), .A1 (n_3029), .A2 (n_3054));
AOI21_X1 i_3091 (.ZN (n_3027), .A (n_3416), .B1 (n_3417), .B2 (n_3415));
NAND3_X1 i_3090 (.ZN (n_3026), .A1 (n_3417), .A2 (n_3416), .A3 (n_3415));
INV_X1 i_3089 (.ZN (n_3025), .A (n_3026));
OAI22_X1 i_3088 (.ZN (n_3024), .A1 (n_3029), .A2 (n_3054), .B1 (n_3027), .B2 (n_3025));
NAND2_X1 i_3087 (.ZN (n_3023), .A1 (n_3024), .A2 (n_3028));
NAND2_X1 i_3086 (.ZN (n_3022), .A1 (n_3023), .A2 (n_3058));
INV_X1 i_3085 (.ZN (n_3021), .A (n_3058));
NAND3_X2 i_3084 (.ZN (n_3020), .A1 (n_3024), .A2 (n_3021), .A3 (n_3028));
INV_X1 i_3083 (.ZN (n_3019), .A (n_3020));
INV_X1 i_3082 (.ZN (n_3018), .A (n_3403));
NAND3_X1 i_3081 (.ZN (n_3017), .A1 (n_3407), .A2 (n_3410), .A3 (n_3018));
INV_X1 i_3080 (.ZN (n_3016), .A (n_3017));
AOI21_X1 i_3079 (.ZN (n_3015), .A (n_3018), .B1 (n_3410), .B2 (n_3407));
NOR2_X1 i_3078 (.ZN (n_3014), .A1 (n_3016), .A2 (n_3015));
OAI21_X2 i_3077 (.ZN (n_3013), .A (n_3022), .B1 (n_3019), .B2 (n_3014));
NAND3_X1 i_3076 (.ZN (n_3012), .A1 (n_3013), .A2 (n_3065), .A3 (n_3062));
NAND2_X1 i_3075 (.ZN (n_3011), .A1 (n_3062), .A2 (n_3065));
INV_X1 i_3074 (.ZN (n_3010), .A (n_3013));
NAND2_X2 i_3073 (.ZN (n_3009), .A1 (n_3011), .A2 (n_3010));
NAND4_X1 i_3072 (.ZN (n_3008), .A1 (n_3179), .A2 (n_3176), .A3 (n_3174), .A4 (n_3173));
NAND2_X1 i_3071 (.ZN (n_3007), .A1 (n_3179), .A2 (n_3176));
NAND2_X1 i_3070 (.ZN (n_3006), .A1 (n_3007), .A2 (n_3172));
NAND2_X1 i_3069 (.ZN (n_3005), .A1 (n_3006), .A2 (n_3008));
AOI21_X1 i_3068 (.ZN (n_3004), .A (n_3421), .B1 (n_3422), .B2 (n_3420));
NAND3_X1 i_3067 (.ZN (n_3003), .A1 (n_3422), .A2 (n_3421), .A3 (n_3420));
INV_X1 i_3066 (.ZN (n_3002), .A (n_3003));
AOI21_X1 i_3065 (.ZN (n_3001), .A (n_3438), .B1 (n_3439), .B2 (n_3436));
NAND3_X1 i_3064 (.ZN (n_3000), .A1 (n_3439), .A2 (n_3438), .A3 (n_3436));
INV_X1 i_3063 (.ZN (n_2999), .A (n_3000));
OAI22_X1 i_3062 (.ZN (n_2998), .A1 (n_3004), .A2 (n_3002), .B1 (n_2999), .B2 (n_3001));
INV_X1 i_3061 (.ZN (n_2997), .A (n_3004));
INV_X1 i_3060 (.ZN (n_2996), .A (n_3001));
NAND4_X1 i_3059 (.ZN (n_2995), .A1 (n_2997), .A2 (n_3003), .A3 (n_2996), .A4 (n_3000));
INV_X1 i_3058 (.ZN (n_2994), .A (n_2995));
OAI22_X1 i_3057 (.ZN (n_2993), .A1 (n_8908), .A2 (n_6677), .B1 (n_8955), .B2 (n_4366));
NAND2_X1 i_3056 (.ZN (n_2992), .A1 (A_imm[18]), .A2 (B_imm[0]));
NAND4_X1 i_3055 (.ZN (n_2991), .A1 (B_imm[16]), .A2 (A_imm[17]), .A3 (B_imm[1]), .A4 (A_imm[2]));
NAND2_X1 i_3054 (.ZN (n_2990), .A1 (n_2991), .A2 (n_2992));
NAND2_X1 i_3053 (.ZN (n_2989), .A1 (n_2990), .A2 (n_2993));
OAI21_X1 i_3052 (.ZN (n_2988), .A (n_2989), .B1 (n_8829), .B2 (n_6678));
NAND2_X1 i_3051 (.ZN (n_2987), .A1 (B_imm[13]), .A2 (A_imm[6]));
NAND4_X1 i_3050 (.ZN (n_2986), .A1 (n_2990), .A2 (n_2993), .A3 (B_imm[15]), .A4 (A_imm[4]));
NAND2_X1 i_3049 (.ZN (n_2985), .A1 (n_2986), .A2 (n_2987));
NAND2_X1 i_3048 (.ZN (n_2984), .A1 (n_2985), .A2 (n_2988));
OAI21_X1 i_3047 (.ZN (n_2983), .A (n_2998), .B1 (n_2984), .B2 (n_2994));
INV_X1 i_3046 (.ZN (n_2982), .A (n_3196));
OAI21_X1 i_3045 (.ZN (n_2981), .A (n_3178), .B1 (n_3181), .B2 (n_2982));
NAND3_X1 i_3044 (.ZN (n_2980), .A1 (n_3182), .A2 (n_3196), .A3 (n_3185));
NAND2_X1 i_3043 (.ZN (n_2979), .A1 (n_2981), .A2 (n_2980));
NAND2_X1 i_3042 (.ZN (n_2978), .A1 (n_2979), .A2 (n_2983));
INV_X1 i_3041 (.ZN (n_2977), .A (n_2984));
NAND2_X1 i_3040 (.ZN (n_2976), .A1 (n_2977), .A2 (n_2995));
NAND4_X1 i_3039 (.ZN (n_2975), .A1 (n_2981), .A2 (n_2976), .A3 (n_2998), .A4 (n_2980));
AOI21_X1 i_3038 (.ZN (n_2974), .A (n_3202), .B1 (n_3203), .B2 (n_3201));
NAND3_X1 i_3037 (.ZN (n_2973), .A1 (n_3203), .A2 (n_3202), .A3 (n_3201));
INV_X1 i_3036 (.ZN (n_2972), .A (n_2973));
OAI211_X1 i_3035 (.ZN (n_2971), .A (B_imm[14]), .B (A_imm[6]), .C1 (n_2974), .C2 (n_2972));
NOR2_X1 i_3034 (.ZN (n_2970), .A1 (n_2974), .A2 (n_2972));
OAI21_X1 i_3033 (.ZN (n_2969), .A (n_2970), .B1 (n_7913), .B2 (n_7691));
NAND2_X1 i_3032 (.ZN (n_2968), .A1 (n_3190), .A2 (n_3187));
NAND2_X1 i_3031 (.ZN (n_2967), .A1 (n_2968), .A2 (n_3188));
NAND3_X1 i_3030 (.ZN (n_2966), .A1 (n_3190), .A2 (n_3189), .A3 (n_3187));
NAND2_X1 i_3029 (.ZN (n_2965), .A1 (n_2967), .A2 (n_2966));
NAND2_X1 i_3028 (.ZN (n_2964), .A1 (n_2969), .A2 (n_2965));
NAND2_X1 i_3027 (.ZN (n_2963), .A1 (n_2964), .A2 (n_2971));
NAND2_X1 i_3026 (.ZN (n_2962), .A1 (n_2963), .A2 (n_2975));
NAND2_X1 i_3025 (.ZN (n_2961), .A1 (n_2962), .A2 (n_2978));
NAND2_X1 i_3024 (.ZN (n_2960), .A1 (n_2961), .A2 (n_3005));
NAND4_X1 i_3023 (.ZN (n_2959), .A1 (n_2962), .A2 (n_3006), .A3 (n_3008), .A4 (n_2978));
NAND4_X1 i_3022 (.ZN (n_2958), .A1 (n_3247), .A2 (n_3243), .A3 (n_3240), .A4 (n_3239));
NAND2_X1 i_3021 (.ZN (n_2957), .A1 (n_3247), .A2 (n_3243));
NAND2_X1 i_3020 (.ZN (n_2956), .A1 (n_2957), .A2 (n_3238));
NAND2_X1 i_3019 (.ZN (n_2955), .A1 (n_2958), .A2 (n_2956));
NAND2_X1 i_3018 (.ZN (n_2954), .A1 (n_2955), .A2 (n_2959));
NAND2_X2 i_3017 (.ZN (n_2953), .A1 (n_2954), .A2 (n_2960));
NAND2_X2 i_3016 (.ZN (n_2952), .A1 (n_3009), .A2 (n_2953));
NAND2_X1 i_3015 (.ZN (n_2951), .A1 (n_2952), .A2 (n_3012));
NAND2_X2 i_3014 (.ZN (n_2950), .A1 (n_2951), .A2 (n_3066));
INV_X1 i_3013 (.ZN (n_2949), .A (n_3066));
NAND3_X1 i_3012 (.ZN (n_2948), .A1 (n_2952), .A2 (n_2949), .A3 (n_3012));
NAND3_X1 i_3011 (.ZN (n_2947), .A1 (n_3159), .A2 (n_3158), .A3 (n_3153));
INV_X1 i_3010 (.ZN (n_2946), .A (n_3153));
NAND2_X1 i_3009 (.ZN (n_2945), .A1 (n_3159), .A2 (n_3158));
NAND2_X1 i_3008 (.ZN (n_2944), .A1 (n_2945), .A2 (n_2946));
NAND2_X1 i_3007 (.ZN (n_2943), .A1 (n_2944), .A2 (n_2947));
NAND2_X1 i_3006 (.ZN (n_2942), .A1 (n_2948), .A2 (n_2943));
NAND2_X1 i_3005 (.ZN (n_2941), .A1 (n_2942), .A2 (n_2950));
NAND2_X2 i_3004 (.ZN (n_2940), .A1 (n_2941), .A2 (n_3069));
NAND4_X2 i_3003 (.ZN (n_2939), .A1 (n_2942), .A2 (n_3070), .A3 (n_2950), .A4 (n_3071));
NAND3_X1 i_3002 (.ZN (n_2938), .A1 (n_3151), .A2 (n_3149), .A3 (n_3145));
AOI21_X1 i_3001 (.ZN (n_2937), .A (n_3150), .B1 (n_3217), .B2 (n_3225));
INV_X1 i_3000 (.ZN (n_2936), .A (n_3149));
INV_X1 i_2999 (.ZN (n_2935), .A (n_3145));
OAI21_X2 i_2998 (.ZN (n_2934), .A (n_2935), .B1 (n_2936), .B2 (n_2937));
NAND3_X2 i_2997 (.ZN (n_2933), .A1 (n_2934), .A2 (n_2939), .A3 (n_2938));
AOI22_X2 i_2996 (.ZN (n_2932), .A1 (n_3072), .A2 (n_3075), .B1 (n_2940), .B2 (n_2933));
INV_X2 i_2995 (.ZN (n_2931), .A (n_2932));
NAND4_X1 i_2994 (.ZN (n_2930), .A1 (n_3358), .A2 (n_3366), .A3 (n_3142), .A4 (n_3137));
NAND2_X2 i_2993 (.ZN (n_2929), .A1 (n_3135), .A2 (n_2930));
NAND2_X4 i_2992 (.ZN (n_2928), .A1 (n_2929), .A2 (n_2931));
NAND2_X1 i_2991 (.ZN (n_2927), .A1 (n_2934), .A2 (n_2938));
NAND3_X1 i_2990 (.ZN (n_2926), .A1 (n_2927), .A2 (n_2940), .A3 (n_2939));
NAND2_X1 i_2989 (.ZN (n_2925), .A1 (n_2940), .A2 (n_2939));
NAND3_X1 i_2988 (.ZN (n_2924), .A1 (n_2925), .A2 (n_2938), .A3 (n_2934));
NAND2_X1 i_2987 (.ZN (n_2923), .A1 (n_2926), .A2 (n_2924));
INV_X1 i_2986 (.ZN (n_2922), .A (n_3218));
NAND3_X1 i_2985 (.ZN (n_2921), .A1 (n_3225), .A2 (n_3220), .A3 (n_2922));
NAND2_X1 i_2984 (.ZN (n_2920), .A1 (n_3225), .A2 (n_3220));
NAND2_X2 i_2983 (.ZN (n_2919), .A1 (n_2920), .A2 (n_3218));
NAND2_X1 i_2982 (.ZN (n_2918), .A1 (n_2919), .A2 (n_2921));
INV_X1 i_2981 (.ZN (n_2917), .A (n_3227));
NAND3_X1 i_2980 (.ZN (n_2916), .A1 (n_3235), .A2 (n_2917), .A3 (n_3233));
INV_X1 i_2979 (.ZN (n_2915), .A (n_3274));
AOI22_X1 i_2978 (.ZN (n_2914), .A1 (n_3237), .A2 (n_3247), .B1 (n_2915), .B2 (n_3276));
OAI21_X1 i_2977 (.ZN (n_2913), .A (n_3227), .B1 (n_3232), .B2 (n_2914));
NAND2_X1 i_2976 (.ZN (n_2912), .A1 (n_2913), .A2 (n_2916));
INV_X1 i_2975 (.ZN (n_2911), .A (n_2912));
AOI21_X1 i_2974 (.ZN (n_2910), .A (n_3289), .B1 (n_3294), .B2 (n_3297));
NAND3_X1 i_2973 (.ZN (n_2909), .A1 (n_3294), .A2 (n_3297), .A3 (n_3289));
INV_X1 i_2972 (.ZN (n_2908), .A (n_2909));
NOR2_X1 i_2971 (.ZN (n_2907), .A1 (n_2908), .A2 (n_2910));
INV_X1 i_2970 (.ZN (n_2906), .A (n_3299));
NAND3_X1 i_2969 (.ZN (n_2905), .A1 (n_3305), .A2 (n_3304), .A3 (n_2906));
NAND2_X1 i_2968 (.ZN (n_2904), .A1 (n_3305), .A2 (n_3304));
NAND2_X1 i_2967 (.ZN (n_2903), .A1 (n_2904), .A2 (n_3299));
NAND2_X1 i_2966 (.ZN (n_2902), .A1 (n_2903), .A2 (n_2905));
NAND2_X1 i_2965 (.ZN (n_2901), .A1 (n_3264), .A2 (n_3262));
NAND3_X1 i_2964 (.ZN (n_2900), .A1 (n_2901), .A2 (B_imm[9]), .A3 (A_imm[11]));
NAND3_X1 i_2963 (.ZN (n_2899), .A1 (n_3264), .A2 (n_3263), .A3 (n_3262));
NAND2_X1 i_2962 (.ZN (n_2898), .A1 (n_2900), .A2 (n_2899));
INV_X1 i_2961 (.ZN (n_2897), .A (n_3194));
NAND2_X1 i_2960 (.ZN (n_2896), .A1 (n_3195), .A2 (n_3193));
NAND2_X1 i_2959 (.ZN (n_2895), .A1 (n_2896), .A2 (n_2897));
NAND3_X1 i_2958 (.ZN (n_2894), .A1 (n_3195), .A2 (n_3194), .A3 (n_3193));
NAND2_X1 i_2957 (.ZN (n_2893), .A1 (n_2895), .A2 (n_2894));
NAND3_X1 i_2956 (.ZN (n_2892), .A1 (n_2893), .A2 (B_imm[19]), .A3 (A_imm[0]));
OAI211_X1 i_2955 (.ZN (n_2891), .A (n_2895), .B (n_2894), .C1 (n_8525), .C2 (n_3554));
AOI22_X1 i_2954 (.ZN (n_2890), .A1 (B_imm[12]), .A2 (A_imm[6]), .B1 (B_imm[8]), .B2 (A_imm[10]));
NAND2_X1 i_2953 (.ZN (n_2889), .A1 (B_imm[11]), .A2 (A_imm[7]));
NAND4_X1 i_2952 (.ZN (n_2888), .A1 (B_imm[12]), .A2 (B_imm[8]), .A3 (A_imm[10]), .A4 (A_imm[6]));
AOI21_X1 i_2951 (.ZN (n_2887), .A (n_2890), .B1 (n_2889), .B2 (n_2888));
NAND2_X1 i_2950 (.ZN (n_2886), .A1 (n_2887), .A2 (n_2891));
NAND2_X1 i_2949 (.ZN (n_2885), .A1 (n_2886), .A2 (n_2892));
NAND2_X1 i_2948 (.ZN (n_2884), .A1 (n_2898), .A2 (n_2885));
INV_X1 i_2947 (.ZN (n_2883), .A (n_3332));
NAND2_X1 i_2946 (.ZN (n_2882), .A1 (n_3344), .A2 (n_3331));
NAND2_X1 i_2945 (.ZN (n_2881), .A1 (n_2882), .A2 (n_2883));
NAND3_X1 i_2944 (.ZN (n_2880), .A1 (n_3344), .A2 (n_3332), .A3 (n_3331));
NAND2_X1 i_2943 (.ZN (n_2879), .A1 (n_2881), .A2 (n_2880));
NAND4_X1 i_2942 (.ZN (n_2878), .A1 (n_2900), .A2 (n_2886), .A3 (n_2899), .A4 (n_2892));
NAND2_X1 i_2941 (.ZN (n_2877), .A1 (n_2878), .A2 (n_2879));
NAND2_X1 i_2940 (.ZN (n_2876), .A1 (n_2877), .A2 (n_2884));
NAND2_X1 i_2939 (.ZN (n_2875), .A1 (n_2902), .A2 (n_2876));
NAND4_X1 i_2938 (.ZN (n_2874), .A1 (n_2903), .A2 (n_2877), .A3 (n_2905), .A4 (n_2884));
OAI22_X2 i_2937 (.ZN (n_2873), .A1 (n_6577), .A2 (n_8927), .B1 (n_8946), .B2 (n_6584));
NAND2_X1 i_2936 (.ZN (n_2872), .A1 (A_imm[10]), .A2 (B_imm[7]));
NAND4_X1 i_2935 (.ZN (n_2871), .A1 (A_imm[13]), .A2 (A_imm[15]), .A3 (B_imm[4]), .A4 (B_imm[2]));
NAND2_X1 i_2934 (.ZN (n_2870), .A1 (n_2871), .A2 (n_2872));
NAND2_X1 i_2933 (.ZN (n_2869), .A1 (n_2870), .A2 (n_2873));
OAI21_X1 i_2932 (.ZN (n_2868), .A (n_2869), .B1 (n_8423), .B2 (n_3554));
NAND2_X1 i_2931 (.ZN (n_2867), .A1 (B_imm[9]), .A2 (A_imm[9]));
NAND4_X1 i_2930 (.ZN (n_2866), .A1 (n_2870), .A2 (n_2873), .A3 (B_imm[18]), .A4 (A_imm[0]));
NAND2_X1 i_2929 (.ZN (n_2865), .A1 (n_2866), .A2 (n_2867));
NAND2_X1 i_2928 (.ZN (n_2864), .A1 (B_imm[6]), .A2 (A_imm[12]));
OAI21_X1 i_2927 (.ZN (n_2863), .A (n_2864), .B1 (n_8858), .B2 (n_6584));
OAI22_X1 i_2926 (.ZN (n_2862), .A1 (n_8880), .A2 (n_8644), .B1 (n_8909), .B2 (n_3554));
NAND2_X1 i_2925 (.ZN (n_2861), .A1 (A_imm[14]), .A2 (B_imm[3]));
INV_X1 i_2924 (.ZN (n_2860), .A (n_2861));
NAND4_X1 i_2923 (.ZN (n_2859), .A1 (B_imm[10]), .A2 (B_imm[17]), .A3 (A_imm[7]), .A4 (A_imm[0]));
INV_X1 i_2922 (.ZN (n_2858), .A (n_2859));
OAI21_X1 i_2921 (.ZN (n_2857), .A (n_2862), .B1 (n_2858), .B2 (n_2860));
NAND4_X1 i_2920 (.ZN (n_2856), .A1 (A_imm[16]), .A2 (B_imm[6]), .A3 (A_imm[12]), .A4 (B_imm[2]));
NAND2_X1 i_2919 (.ZN (n_2855), .A1 (n_2856), .A2 (n_2857));
NAND2_X1 i_2918 (.ZN (n_2854), .A1 (n_2855), .A2 (n_2863));
INV_X1 i_2917 (.ZN (n_2853), .A (n_2854));
NAND3_X1 i_2916 (.ZN (n_2852), .A1 (n_2865), .A2 (n_2868), .A3 (n_2853));
AOI22_X1 i_2915 (.ZN (n_2851), .A1 (n_2865), .A2 (n_2868), .B1 (n_2863), .B2 (n_2855));
NAND2_X1 i_2914 (.ZN (n_2850), .A1 (n_3269), .A2 (n_3267));
INV_X1 i_2913 (.ZN (n_2849), .A (n_2850));
NOR2_X1 i_2912 (.ZN (n_2848), .A1 (n_2849), .A2 (n_3268));
NAND2_X1 i_2911 (.ZN (n_2847), .A1 (n_2849), .A2 (n_3268));
INV_X1 i_2910 (.ZN (n_2846), .A (n_2847));
NOR2_X1 i_2909 (.ZN (n_2845), .A1 (n_2846), .A2 (n_2848));
OAI21_X2 i_2908 (.ZN (n_2844), .A (n_2852), .B1 (n_2851), .B2 (n_2845));
INV_X1 i_2907 (.ZN (n_2843), .A (n_3309));
NAND2_X1 i_2906 (.ZN (n_2842), .A1 (n_3310), .A2 (n_3308));
NAND2_X1 i_2905 (.ZN (n_2841), .A1 (n_2842), .A2 (n_2843));
NAND3_X1 i_2904 (.ZN (n_2840), .A1 (n_3310), .A2 (n_3309), .A3 (n_3308));
NAND2_X1 i_2903 (.ZN (n_2839), .A1 (n_2841), .A2 (n_2840));
NOR2_X1 i_2902 (.ZN (n_2838), .A1 (n_2844), .A2 (n_2839));
NAND2_X1 i_2901 (.ZN (n_2837), .A1 (n_2844), .A2 (n_2839));
NAND2_X1 i_2900 (.ZN (n_2836), .A1 (n_3315), .A2 (n_3313));
NAND3_X1 i_2899 (.ZN (n_2835), .A1 (n_2836), .A2 (B_imm[7]), .A3 (A_imm[12]));
NAND3_X1 i_2898 (.ZN (n_2834), .A1 (n_3315), .A2 (n_3314), .A3 (n_3313));
OAI211_X1 i_2897 (.ZN (n_2833), .A (n_2835), .B (n_2834), .C1 (n_7913), .C2 (n_8293));
NAND2_X1 i_2896 (.ZN (n_2832), .A1 (n_2835), .A2 (n_2834));
NAND3_X1 i_2895 (.ZN (n_2831), .A1 (n_2832), .A2 (B_imm[14]), .A3 (A_imm[5]));
OAI22_X1 i_2894 (.ZN (n_2830), .A1 (n_8908), .A2 (n_6836), .B1 (n_8955), .B2 (n_6740));
NAND2_X1 i_2893 (.ZN (n_2829), .A1 (A_imm[12]), .A2 (B_imm[5]));
NAND4_X1 i_2892 (.ZN (n_2828), .A1 (B_imm[16]), .A2 (A_imm[17]), .A3 (B_imm[0]), .A4 (A_imm[1]));
NAND2_X1 i_2891 (.ZN (n_2827), .A1 (n_2828), .A2 (n_2829));
NAND2_X1 i_2890 (.ZN (n_2826), .A1 (n_2827), .A2 (n_2830));
OAI21_X1 i_2889 (.ZN (n_2825), .A (n_2826), .B1 (n_8829), .B2 (n_3718));
NAND2_X1 i_2888 (.ZN (n_2824), .A1 (B_imm[13]), .A2 (A_imm[5]));
INV_X1 i_2887 (.ZN (n_2823), .A (n_2824));
NAND4_X1 i_2886 (.ZN (n_2822), .A1 (n_2827), .A2 (n_2830), .A3 (B_imm[15]), .A4 (A_imm[3]));
INV_X1 i_2885 (.ZN (n_2821), .A (n_2822));
OAI21_X1 i_2884 (.ZN (n_2820), .A (n_2825), .B1 (n_2821), .B2 (n_2823));
NAND2_X1 i_2883 (.ZN (n_2819), .A1 (n_2831), .A2 (n_2820));
NAND2_X1 i_2882 (.ZN (n_2818), .A1 (n_2819), .A2 (n_2833));
AOI21_X1 i_2881 (.ZN (n_2817), .A (n_2838), .B1 (n_2837), .B2 (n_2818));
NAND2_X1 i_2880 (.ZN (n_2816), .A1 (n_2874), .A2 (n_2817));
NAND2_X1 i_2879 (.ZN (n_2815), .A1 (n_2816), .A2 (n_2875));
NAND2_X1 i_2878 (.ZN (n_2814), .A1 (n_2907), .A2 (n_2815));
OAI211_X1 i_2877 (.ZN (n_2813), .A (n_2816), .B (n_2875), .C1 (n_2908), .C2 (n_2910));
AOI21_X1 i_2876 (.ZN (n_2812), .A (n_3318), .B1 (n_3329), .B2 (n_3326));
NAND3_X1 i_2875 (.ZN (n_2811), .A1 (n_3326), .A2 (n_3318), .A3 (n_3329));
INV_X1 i_2874 (.ZN (n_2810), .A (n_2811));
NOR2_X1 i_2873 (.ZN (n_2809), .A1 (n_2810), .A2 (n_2812));
NAND3_X1 i_2872 (.ZN (n_2808), .A1 (n_3246), .A2 (n_3256), .A3 (n_3249));
INV_X1 i_2871 (.ZN (n_2807), .A (n_2808));
AOI21_X1 i_2870 (.ZN (n_2806), .A (n_3249), .B1 (n_3246), .B2 (n_3256));
OAI21_X1 i_2869 (.ZN (n_2805), .A (n_2809), .B1 (n_2807), .B2 (n_2806));
NOR2_X1 i_2868 (.ZN (n_2804), .A1 (n_2806), .A2 (n_2807));
OAI21_X1 i_2867 (.ZN (n_2803), .A (n_2804), .B1 (n_2812), .B2 (n_2810));
INV_X1 i_2866 (.ZN (n_2802), .A (n_2803));
NAND4_X1 i_2865 (.ZN (n_2801), .A1 (n_3030), .A2 (n_3056), .A3 (n_3055), .A4 (n_3045));
NOR2_X1 i_2864 (.ZN (n_2800), .A1 (n_3025), .A2 (n_3027));
NAND3_X1 i_2863 (.ZN (n_2799), .A1 (n_3028), .A2 (n_2801), .A3 (n_2800));
INV_X1 i_2862 (.ZN (n_2798), .A (n_2799));
AOI21_X1 i_2861 (.ZN (n_2797), .A (n_2800), .B1 (n_3028), .B2 (n_2801));
NOR2_X1 i_2860 (.ZN (n_2796), .A1 (n_2798), .A2 (n_2797));
OAI21_X1 i_2859 (.ZN (n_2795), .A (n_2805), .B1 (n_2796), .B2 (n_2802));
NAND2_X2 i_2858 (.ZN (n_2794), .A1 (n_2813), .A2 (n_2795));
NAND2_X1 i_2857 (.ZN (n_2793), .A1 (n_2794), .A2 (n_2814));
NAND2_X1 i_2856 (.ZN (n_2792), .A1 (n_2793), .A2 (n_2911));
NAND3_X2 i_2855 (.ZN (n_2791), .A1 (n_2794), .A2 (n_2912), .A3 (n_2814));
NAND3_X1 i_2854 (.ZN (n_2790), .A1 (n_3224), .A2 (n_3286), .A3 (n_3223));
INV_X1 i_2853 (.ZN (n_2789), .A (n_2790));
AOI21_X1 i_2852 (.ZN (n_2788), .A (n_3223), .B1 (n_3224), .B2 (n_3286));
NOR2_X2 i_2851 (.ZN (n_2787), .A1 (n_2789), .A2 (n_2788));
NAND2_X1 i_2850 (.ZN (n_2786), .A1 (n_2787), .A2 (n_2791));
NAND2_X1 i_2849 (.ZN (n_2785), .A1 (n_2786), .A2 (n_2792));
NAND2_X1 i_2848 (.ZN (n_2784), .A1 (n_2918), .A2 (n_2785));
NAND4_X1 i_2847 (.ZN (n_2783), .A1 (n_2919), .A2 (n_2786), .A3 (n_2921), .A4 (n_2792));
INV_X1 i_2846 (.ZN (n_2782), .A (n_2783));
NAND3_X1 i_2845 (.ZN (n_2781), .A1 (n_2950), .A2 (n_2948), .A3 (n_2943));
AOI22_X1 i_2844 (.ZN (n_2780), .A1 (n_2952), .A2 (n_3012), .B1 (n_3068), .B2 (n_3067));
INV_X1 i_2843 (.ZN (n_2779), .A (n_2948));
INV_X1 i_2842 (.ZN (n_2778), .A (n_2943));
OAI21_X1 i_2841 (.ZN (n_2777), .A (n_2778), .B1 (n_2779), .B2 (n_2780));
NAND2_X2 i_2840 (.ZN (n_2776), .A1 (n_2777), .A2 (n_2781));
OAI21_X1 i_2839 (.ZN (n_2775), .A (n_2784), .B1 (n_2776), .B2 (n_2782));
NAND2_X2 i_2838 (.ZN (n_2774), .A1 (n_2923), .A2 (n_2775));
NAND2_X1 i_2837 (.ZN (n_2773), .A1 (n_2933), .A2 (n_2940));
NAND3_X1 i_2835 (.ZN (n_2771), .A1 (n_3072), .A2 (CLOCK_opt_ipo_n337), .A3 (n_3075));
INV_X1 i_2834 (.ZN (n_2770), .A (n_2771));
OAI21_X2 i_2833 (.ZN (n_2769), .A (n_2774), .B1 (n_2770), .B2 (n_2932));
NAND3_X1 i_2832 (.ZN (n_2768), .A1 (n_2776), .A2 (n_2784), .A3 (n_2783));
INV_X1 i_2831 (.ZN (n_2767), .A (n_2776));
NAND2_X1 i_2830 (.ZN (n_2766), .A1 (n_2784), .A2 (n_2783));
NAND2_X1 i_2829 (.ZN (n_2765), .A1 (n_2766), .A2 (n_2767));
NAND3_X1 i_2828 (.ZN (n_2764), .A1 (n_3009), .A2 (n_3012), .A3 (n_2953));
INV_X1 i_2827 (.ZN (n_2763), .A (n_2764));
AOI21_X2 i_2826 (.ZN (n_2762), .A (n_2953), .B1 (n_3012), .B2 (n_3009));
NOR2_X1 i_2825 (.ZN (n_2761), .A1 (n_2763), .A2 (n_2762));
INV_X1 i_2824 (.ZN (n_2760), .A (n_3014));
NAND3_X1 i_2823 (.ZN (n_2759), .A1 (n_3022), .A2 (n_2760), .A3 (n_3020));
AOI21_X1 i_2822 (.ZN (n_2758), .A (n_3021), .B1 (n_3028), .B2 (n_3024));
OAI21_X1 i_2821 (.ZN (n_2757), .A (n_3014), .B1 (n_2758), .B2 (n_3019));
NAND2_X1 i_2820 (.ZN (n_2756), .A1 (n_2757), .A2 (n_2759));
INV_X1 i_2819 (.ZN (n_2755), .A (n_2756));
NAND3_X1 i_2818 (.ZN (n_2754), .A1 (n_2978), .A2 (n_2963), .A3 (n_2975));
INV_X1 i_2817 (.ZN (n_2753), .A (n_2963));
NAND2_X1 i_2816 (.ZN (n_2752), .A1 (n_2978), .A2 (n_2975));
NAND2_X1 i_2815 (.ZN (n_2751), .A1 (n_2752), .A2 (n_2753));
NAND2_X1 i_2814 (.ZN (n_2750), .A1 (n_3342), .A2 (n_3334));
NAND2_X1 i_2813 (.ZN (n_2749), .A1 (n_2750), .A2 (n_3335));
NAND3_X1 i_2812 (.ZN (n_2748), .A1 (n_3342), .A2 (n_3336), .A3 (n_3334));
AOI21_X1 i_2811 (.ZN (n_2747), .A (n_3052), .B1 (n_3053), .B2 (n_3051));
INV_X1 i_2810 (.ZN (n_2746), .A (n_2747));
NAND3_X1 i_2809 (.ZN (n_2745), .A1 (n_3053), .A2 (n_3052), .A3 (n_3051));
NAND4_X1 i_2808 (.ZN (n_2744), .A1 (n_2746), .A2 (n_2749), .A3 (n_2748), .A4 (n_2745));
NAND2_X1 i_2807 (.ZN (n_2743), .A1 (n_2749), .A2 (n_2748));
INV_X1 i_2806 (.ZN (n_2742), .A (n_2745));
OAI21_X1 i_2805 (.ZN (n_2741), .A (n_2743), .B1 (n_2747), .B2 (n_2742));
OAI22_X1 i_2804 (.ZN (n_2740), .A1 (n_8795), .A2 (n_8293), .B1 (n_8947), .B2 (n_8645));
NAND2_X1 i_2803 (.ZN (n_2739), .A1 (B_imm[11]), .A2 (A_imm[6]));
NAND4_X1 i_2802 (.ZN (n_2738), .A1 (B_imm[12]), .A2 (B_imm[8]), .A3 (A_imm[9]), .A4 (A_imm[5]));
NAND2_X1 i_2801 (.ZN (n_2737), .A1 (n_2738), .A2 (n_2739));
NAND2_X1 i_2800 (.ZN (n_2736), .A1 (n_2737), .A2 (n_2740));
NAND2_X1 i_2799 (.ZN (n_2735), .A1 (n_3341), .A2 (n_3338));
NAND2_X1 i_2798 (.ZN (n_2734), .A1 (n_2735), .A2 (n_3339));
NAND3_X1 i_2797 (.ZN (n_2733), .A1 (n_3341), .A2 (n_3340), .A3 (n_3338));
NAND3_X1 i_2796 (.ZN (n_2732), .A1 (n_2736), .A2 (n_2734), .A3 (n_2733));
OAI22_X1 i_2795 (.ZN (n_2731), .A1 (n_4366), .A2 (n_8858), .B1 (n_8232), .B2 (n_8926));
NAND2_X1 i_2794 (.ZN (n_2730), .A1 (A_imm[11]), .A2 (B_imm[5]));
OAI21_X1 i_2793 (.ZN (n_2729), .A (n_2730), .B1 (n_8880), .B2 (n_7691));
NAND2_X1 i_2792 (.ZN (n_2728), .A1 (A_imm[14]), .A2 (B_imm[2]));
INV_X1 i_2791 (.ZN (n_2727), .A (n_2728));
NAND4_X1 i_2790 (.ZN (n_2726), .A1 (B_imm[10]), .A2 (A_imm[11]), .A3 (B_imm[5]), .A4 (A_imm[6]));
INV_X1 i_2789 (.ZN (n_2725), .A (n_2726));
OAI21_X1 i_2788 (.ZN (n_2724), .A (n_2729), .B1 (n_2725), .B2 (n_2727));
INV_X1 i_2787 (.ZN (n_2723), .A (n_2724));
NAND4_X1 i_2786 (.ZN (n_2722), .A1 (A_imm[16]), .A2 (B_imm[6]), .A3 (B_imm[1]), .A4 (A_imm[11]));
INV_X1 i_2785 (.ZN (n_2721), .A (n_2722));
OAI21_X1 i_2784 (.ZN (n_2720), .A (n_2731), .B1 (n_2723), .B2 (n_2721));
NAND2_X1 i_2783 (.ZN (n_2719), .A1 (n_2734), .A2 (n_2733));
NAND3_X1 i_2782 (.ZN (n_2718), .A1 (n_2737), .A2 (n_2719), .A3 (n_2740));
NAND2_X1 i_2781 (.ZN (n_2717), .A1 (n_2718), .A2 (n_2720));
NAND2_X1 i_2780 (.ZN (n_2716), .A1 (n_2717), .A2 (n_2732));
NAND2_X1 i_2779 (.ZN (n_2715), .A1 (n_2716), .A2 (n_2741));
NAND2_X1 i_2778 (.ZN (n_2714), .A1 (n_3031), .A2 (n_3045));
NAND2_X1 i_2777 (.ZN (n_2713), .A1 (n_2714), .A2 (n_3034));
NAND3_X1 i_2776 (.ZN (n_2712), .A1 (n_3031), .A2 (n_3033), .A3 (n_3045));
NAND4_X1 i_2775 (.ZN (n_2711), .A1 (n_2715), .A2 (n_2713), .A3 (n_2744), .A4 (n_2712));
INV_X1 i_2774 (.ZN (n_2710), .A (n_2711));
NAND2_X1 i_2773 (.ZN (n_2709), .A1 (n_2715), .A2 (n_2744));
NAND2_X1 i_2772 (.ZN (n_2708), .A1 (n_2713), .A2 (n_2712));
NAND2_X1 i_2771 (.ZN (n_2707), .A1 (n_2709), .A2 (n_2708));
AOI21_X1 i_2770 (.ZN (n_2706), .A (n_2987), .B1 (n_2988), .B2 (n_2986));
NAND3_X1 i_2769 (.ZN (n_2705), .A1 (n_2988), .A2 (n_2987), .A3 (n_2986));
INV_X1 i_2768 (.ZN (n_2704), .A (n_2705));
INV_X1 i_2767 (.ZN (n_2703), .A (n_3039));
OAI21_X1 i_2766 (.ZN (n_2702), .A (n_3037), .B1 (n_2703), .B2 (n_3035));
NAND3_X1 i_2765 (.ZN (n_2701), .A1 (n_3039), .A2 (n_3038), .A3 (n_3036));
NAND2_X1 i_2764 (.ZN (n_2700), .A1 (n_2702), .A2 (n_2701));
OAI21_X1 i_2763 (.ZN (n_2699), .A (n_2700), .B1 (n_2706), .B2 (n_2704));
INV_X1 i_2762 (.ZN (n_2698), .A (n_2706));
NAND4_X1 i_2761 (.ZN (n_2697), .A1 (n_2698), .A2 (n_2702), .A3 (n_2705), .A4 (n_2701));
OAI22_X1 i_2760 (.ZN (n_2696), .A1 (n_6817), .A2 (n_8927), .B1 (n_8645), .B2 (n_8573));
NAND2_X1 i_2759 (.ZN (n_2695), .A1 (A_imm[15]), .A2 (B_imm[1]));
NAND4_X1 i_2758 (.ZN (n_2694), .A1 (A_imm[13]), .A2 (A_imm[9]), .A3 (B_imm[7]), .A4 (B_imm[3]));
NAND2_X1 i_2757 (.ZN (n_2693), .A1 (n_2694), .A2 (n_2695));
NAND2_X1 i_2756 (.ZN (n_2692), .A1 (n_2693), .A2 (n_2696));
OAI21_X1 i_2755 (.ZN (n_2691), .A (n_2692), .B1 (n_8347), .B2 (n_8511));
NAND2_X1 i_2754 (.ZN (n_2690), .A1 (B_imm[15]), .A2 (A_imm[2]));
NAND4_X1 i_2753 (.ZN (n_2689), .A1 (n_2693), .A2 (n_2696), .A3 (B_imm[9]), .A4 (A_imm[8]));
NAND2_X1 i_2752 (.ZN (n_2688), .A1 (n_2689), .A2 (n_2690));
NAND2_X1 i_2751 (.ZN (n_2687), .A1 (n_3044), .A2 (n_3042));
NAND3_X1 i_2750 (.ZN (n_2686), .A1 (n_2687), .A2 (B_imm[3]), .A3 (A_imm[15]));
NAND3_X1 i_2749 (.ZN (n_2685), .A1 (n_3044), .A2 (n_3043), .A3 (n_3042));
NAND2_X1 i_2748 (.ZN (n_2684), .A1 (n_2686), .A2 (n_2685));
NAND3_X1 i_2747 (.ZN (n_2683), .A1 (n_2688), .A2 (n_2691), .A3 (n_2684));
AOI21_X1 i_2746 (.ZN (n_2682), .A (n_2684), .B1 (n_2691), .B2 (n_2688));
NAND2_X1 i_2745 (.ZN (n_2681), .A1 (n_2993), .A2 (n_2991));
XNOR2_X1 i_2744 (.ZN (n_2680), .A (n_2681), .B (n_2992));
OAI21_X1 i_2743 (.ZN (n_2679), .A (n_2683), .B1 (n_2682), .B2 (n_2680));
NAND2_X1 i_2742 (.ZN (n_2678), .A1 (n_2679), .A2 (n_2697));
NAND2_X1 i_2741 (.ZN (n_2677), .A1 (n_2678), .A2 (n_2699));
AOI21_X1 i_2740 (.ZN (n_2676), .A (n_2710), .B1 (n_2677), .B2 (n_2707));
INV_X1 i_2739 (.ZN (n_2675), .A (n_2676));
NAND3_X1 i_2738 (.ZN (n_2674), .A1 (n_2675), .A2 (n_2754), .A3 (n_2751));
NAND2_X1 i_2737 (.ZN (n_2673), .A1 (n_2751), .A2 (n_2754));
NAND2_X1 i_2736 (.ZN (n_2672), .A1 (n_2676), .A2 (n_2673));
AOI21_X1 i_2735 (.ZN (n_2671), .A (n_2965), .B1 (n_2969), .B2 (n_2971));
INV_X1 i_2734 (.ZN (n_2670), .A (n_2671));
NAND3_X1 i_2733 (.ZN (n_2669), .A1 (n_2969), .A2 (n_2971), .A3 (n_2965));
NAND3_X1 i_2732 (.ZN (n_2668), .A1 (n_2984), .A2 (n_2995), .A3 (n_2998));
INV_X1 i_2731 (.ZN (n_2667), .A (n_2998));
OAI21_X1 i_2730 (.ZN (n_2666), .A (n_2977), .B1 (n_2667), .B2 (n_2994));
NAND2_X1 i_2729 (.ZN (n_2665), .A1 (n_2666), .A2 (n_2668));
NAND3_X1 i_2728 (.ZN (n_2664), .A1 (n_2670), .A2 (n_2669), .A3 (n_2665));
INV_X1 i_2727 (.ZN (n_2663), .A (n_2669));
OAI211_X1 i_2726 (.ZN (n_2662), .A (n_2668), .B (n_2666), .C1 (n_2663), .C2 (n_2671));
NAND3_X1 i_2725 (.ZN (n_2661), .A1 (n_2884), .A2 (n_2879), .A3 (n_2878));
NAND2_X1 i_2724 (.ZN (n_2660), .A1 (n_2884), .A2 (n_2878));
NAND3_X1 i_2723 (.ZN (n_2659), .A1 (n_2660), .A2 (n_2881), .A3 (n_2880));
NAND3_X1 i_2722 (.ZN (n_2658), .A1 (n_2662), .A2 (n_2661), .A3 (n_2659));
NAND2_X1 i_2721 (.ZN (n_2657), .A1 (n_2658), .A2 (n_2664));
NAND2_X1 i_2720 (.ZN (n_2656), .A1 (n_2657), .A2 (n_2672));
NAND2_X1 i_2719 (.ZN (n_2655), .A1 (n_2656), .A2 (n_2674));
NAND2_X1 i_2718 (.ZN (n_2654), .A1 (n_2655), .A2 (n_2755));
NAND3_X1 i_2717 (.ZN (n_2653), .A1 (n_2656), .A2 (n_2756), .A3 (n_2674));
NAND3_X1 i_2716 (.ZN (n_2652), .A1 (n_2960), .A2 (n_2955), .A3 (n_2959));
INV_X1 i_2715 (.ZN (n_2651), .A (n_2652));
AOI21_X1 i_2714 (.ZN (n_2650), .A (n_2955), .B1 (n_2960), .B2 (n_2959));
NOR2_X1 i_2713 (.ZN (n_2649), .A1 (n_2651), .A2 (n_2650));
NAND2_X1 i_2712 (.ZN (n_2648), .A1 (n_2653), .A2 (n_2649));
NAND2_X1 i_2711 (.ZN (n_2647), .A1 (n_2648), .A2 (n_2654));
NAND2_X1 i_2710 (.ZN (n_2646), .A1 (n_2647), .A2 (n_2761));
INV_X1 i_2709 (.ZN (n_2645), .A (n_2646));
OAI211_X2 i_2708 (.ZN (n_2644), .A (n_2648), .B (n_2654), .C1 (n_2763), .C2 (n_2762));
INV_X1 i_2707 (.ZN (n_2643), .A (n_2787));
NAND3_X1 i_2706 (.ZN (n_2642), .A1 (n_2792), .A2 (n_2791), .A3 (n_2643));
AOI21_X1 i_2705 (.ZN (n_2641), .A (n_2912), .B1 (n_2814), .B2 (n_2794));
INV_X1 i_2704 (.ZN (n_2640), .A (n_2791));
OAI21_X2 i_2703 (.ZN (n_2639), .A (n_2787), .B1 (n_2640), .B2 (n_2641));
NAND2_X2 i_2702 (.ZN (n_2638), .A1 (n_2639), .A2 (n_2642));
AOI21_X2 i_2701 (.ZN (n_2637), .A (n_2645), .B1 (n_2638), .B2 (n_2644));
AOI21_X2 i_2700 (.ZN (n_2636), .A (n_2637), .B1 (n_2765), .B2 (n_2768));
INV_X1 i_2699 (.ZN (n_2635), .A (n_2636));
INV_X1 i_2698 (.ZN (n_2634), .A (n_2775));
NAND3_X1 i_2697 (.ZN (n_2633), .A1 (n_2926), .A2 (n_2634), .A3 (n_2924));
NAND2_X2 i_2696 (.ZN (n_2632), .A1 (n_2774), .A2 (n_2633));
NAND2_X2 i_2695 (.ZN (n_2631), .A1 (n_2632), .A2 (n_2635));
NAND3_X2 i_2694 (.ZN (n_2630), .A1 (n_2928), .A2 (n_2769), .A3 (n_2631));
NAND3_X1 i_2692 (.ZN (n_2628), .A1 (n_2814), .A2 (n_2813), .A3 (n_2795));
INV_X1 i_2691 (.ZN (n_2627), .A (n_2628));
AOI21_X1 i_2690 (.ZN (n_2626), .A (n_2795), .B1 (n_2814), .B2 (n_2813));
NOR2_X1 i_2689 (.ZN (n_2625), .A1 (n_2627), .A2 (n_2626));
INV_X1 i_2688 (.ZN (n_2624), .A (n_2844));
NAND3_X1 i_2687 (.ZN (n_2623), .A1 (n_2624), .A2 (n_2841), .A3 (n_2840));
INV_X1 i_2686 (.ZN (n_2622), .A (n_2837));
INV_X1 i_2685 (.ZN (n_2621), .A (n_2818));
OAI21_X1 i_2684 (.ZN (n_2620), .A (n_2623), .B1 (n_2622), .B2 (n_2621));
NAND3_X1 i_2683 (.ZN (n_2619), .A1 (n_2875), .A2 (n_2874), .A3 (n_2620));
NAND2_X1 i_2682 (.ZN (n_2618), .A1 (n_2875), .A2 (n_2874));
NAND2_X1 i_2681 (.ZN (n_2617), .A1 (n_2618), .A2 (n_2817));
NAND2_X1 i_2680 (.ZN (n_2616), .A1 (n_2617), .A2 (n_2619));
NAND3_X1 i_2679 (.ZN (n_2615), .A1 (n_2623), .A2 (n_2837), .A3 (n_2818));
OAI21_X1 i_2678 (.ZN (n_2614), .A (n_2621), .B1 (n_2622), .B2 (n_2838));
NAND2_X1 i_2677 (.ZN (n_2613), .A1 (n_2614), .A2 (n_2615));
INV_X1 i_2676 (.ZN (n_2612), .A (n_2887));
NAND2_X1 i_2675 (.ZN (n_2611), .A1 (n_2892), .A2 (n_2891));
NAND2_X1 i_2674 (.ZN (n_2610), .A1 (n_2611), .A2 (n_2612));
NAND3_X1 i_2673 (.ZN (n_2609), .A1 (n_2892), .A2 (n_2887), .A3 (n_2891));
NAND2_X1 i_2672 (.ZN (n_2608), .A1 (n_2610), .A2 (n_2609));
INV_X1 i_2671 (.ZN (n_2607), .A (n_2608));
AOI21_X1 i_2670 (.ZN (n_2606), .A (n_2857), .B1 (n_2863), .B2 (n_2856));
NAND3_X1 i_2669 (.ZN (n_2605), .A1 (n_2863), .A2 (n_2857), .A3 (n_2856));
INV_X1 i_2668 (.ZN (n_2604), .A (n_2605));
OAI211_X1 i_2667 (.ZN (n_2603), .A (B_imm[14]), .B (A_imm[4]), .C1 (n_2606), .C2 (n_2604));
NOR2_X1 i_2666 (.ZN (n_2602), .A1 (n_2604), .A2 (n_2606));
OAI21_X1 i_2665 (.ZN (n_2601), .A (n_2602), .B1 (n_7913), .B2 (n_6678));
OAI22_X1 i_2664 (.ZN (n_2600), .A1 (n_8752), .A2 (n_6577), .B1 (n_8908), .B2 (n_3554));
NAND2_X1 i_2663 (.ZN (n_2599), .A1 (B_imm[6]), .A2 (A_imm[10]));
NAND4_X1 i_2662 (.ZN (n_2598), .A1 (A_imm[12]), .A2 (B_imm[16]), .A3 (B_imm[4]), .A4 (A_imm[0]));
NAND2_X1 i_2661 (.ZN (n_2597), .A1 (n_2598), .A2 (n_2599));
AOI22_X1 i_2660 (.ZN (n_2596), .A1 (n_2597), .A2 (n_2600), .B1 (B_imm[13]), .B2 (A_imm[4]));
INV_X1 i_2659 (.ZN (n_2595), .A (n_2596));
NAND4_X1 i_2658 (.ZN (n_2594), .A1 (n_2597), .A2 (n_2600), .A3 (B_imm[13]), .A4 (A_imm[4]));
INV_X1 i_2657 (.ZN (n_2593), .A (n_2594));
INV_X1 i_2656 (.ZN (n_2592), .A (n_2862));
OAI21_X1 i_2655 (.ZN (n_2591), .A (n_2860), .B1 (n_2592), .B2 (n_2858));
NAND3_X1 i_2654 (.ZN (n_2590), .A1 (n_2862), .A2 (n_2861), .A3 (n_2859));
NAND2_X1 i_2653 (.ZN (n_2589), .A1 (n_2591), .A2 (n_2590));
OAI21_X1 i_2652 (.ZN (n_2588), .A (n_2595), .B1 (n_2593), .B2 (n_2589));
INV_X1 i_2651 (.ZN (n_2587), .A (n_2588));
NAND2_X1 i_2650 (.ZN (n_2586), .A1 (n_2601), .A2 (n_2587));
NAND2_X1 i_2649 (.ZN (n_2585), .A1 (n_2586), .A2 (n_2603));
NAND2_X1 i_2648 (.ZN (n_2584), .A1 (n_2585), .A2 (n_2607));
NAND3_X1 i_2647 (.ZN (n_2583), .A1 (n_2586), .A2 (n_2608), .A3 (n_2603));
INV_X1 i_2646 (.ZN (n_2582), .A (n_2852));
OAI21_X1 i_2645 (.ZN (n_2581), .A (n_2845), .B1 (n_2582), .B2 (n_2851));
INV_X1 i_2644 (.ZN (n_2580), .A (n_2851));
OAI211_X1 i_2643 (.ZN (n_2579), .A (n_2580), .B (n_2852), .C1 (n_2848), .C2 (n_2846));
NAND2_X1 i_2642 (.ZN (n_2578), .A1 (n_2579), .A2 (n_2581));
INV_X1 i_2641 (.ZN (n_2577), .A (n_2578));
NAND2_X1 i_2640 (.ZN (n_2576), .A1 (n_2577), .A2 (n_2583));
NAND2_X1 i_2639 (.ZN (n_2575), .A1 (n_2576), .A2 (n_2584));
NAND2_X1 i_2638 (.ZN (n_2574), .A1 (n_2613), .A2 (n_2575));
NAND4_X1 i_2637 (.ZN (n_2573), .A1 (n_2614), .A2 (n_2576), .A3 (n_2615), .A4 (n_2584));
AOI21_X1 i_2636 (.ZN (n_2572), .A (n_2867), .B1 (n_2868), .B2 (n_2866));
NAND3_X1 i_2635 (.ZN (n_2571), .A1 (n_2868), .A2 (n_2867), .A3 (n_2866));
INV_X1 i_2634 (.ZN (n_2570), .A (n_2571));
INV_X1 i_2633 (.ZN (n_2569), .A (n_2889));
INV_X1 i_2632 (.ZN (n_2568), .A (n_2888));
OAI21_X1 i_2631 (.ZN (n_2567), .A (n_2569), .B1 (n_2568), .B2 (n_2890));
INV_X1 i_2630 (.ZN (n_2566), .A (n_2890));
NAND3_X1 i_2629 (.ZN (n_2565), .A1 (n_2566), .A2 (n_2889), .A3 (n_2888));
NAND2_X1 i_2628 (.ZN (n_2564), .A1 (n_2565), .A2 (n_2567));
OAI21_X1 i_2627 (.ZN (n_2563), .A (n_2564), .B1 (n_2570), .B2 (n_2572));
INV_X1 i_2626 (.ZN (n_2562), .A (n_2572));
INV_X1 i_2625 (.ZN (n_2561), .A (n_2564));
NAND3_X1 i_2624 (.ZN (n_2560), .A1 (n_2561), .A2 (n_2562), .A3 (n_2571));
INV_X1 i_2623 (.ZN (n_2559), .A (n_2560));
NAND2_X1 i_2622 (.ZN (n_2558), .A1 (B_imm[12]), .A2 (A_imm[4]));
OAI21_X1 i_2621 (.ZN (n_2557), .A (n_2558), .B1 (n_8849), .B2 (n_8293));
OAI22_X1 i_2620 (.ZN (n_2556), .A1 (n_8927), .A2 (n_6584), .B1 (n_8971), .B2 (n_4366));
NAND2_X1 i_2619 (.ZN (n_2555), .A1 (A_imm[15]), .A2 (B_imm[0]));
NAND4_X1 i_2618 (.ZN (n_2554), .A1 (A_imm[13]), .A2 (B_imm[2]), .A3 (B_imm[1]), .A4 (A_imm[14]));
NAND2_X1 i_2617 (.ZN (n_2553), .A1 (n_2554), .A2 (n_2555));
NAND2_X1 i_2616 (.ZN (n_2552), .A1 (n_2553), .A2 (n_2556));
NAND4_X1 i_2615 (.ZN (n_2551), .A1 (B_imm[11]), .A2 (B_imm[12]), .A3 (A_imm[5]), .A4 (A_imm[4]));
NAND2_X1 i_2614 (.ZN (n_2550), .A1 (n_2551), .A2 (n_2552));
NAND2_X1 i_2613 (.ZN (n_2549), .A1 (A_imm[16]), .A2 (B_imm[0]));
NAND2_X1 i_2612 (.ZN (n_2548), .A1 (A_imm[11]), .A2 (B_imm[4]));
OAI21_X1 i_2611 (.ZN (n_2547), .A (n_2548), .B1 (n_8880), .B2 (n_8293));
NAND2_X1 i_2610 (.ZN (n_2546), .A1 (B_imm[7]), .A2 (A_imm[8]));
INV_X1 i_2609 (.ZN (n_2545), .A (n_2546));
NAND4_X1 i_2608 (.ZN (n_2544), .A1 (B_imm[10]), .A2 (A_imm[11]), .A3 (B_imm[4]), .A4 (A_imm[5]));
INV_X1 i_2607 (.ZN (n_2543), .A (n_2544));
OAI21_X1 i_2606 (.ZN (n_2542), .A (n_2547), .B1 (n_2543), .B2 (n_2545));
NAND2_X1 i_2605 (.ZN (n_2541), .A1 (n_2542), .A2 (n_2549));
NAND2_X1 i_2604 (.ZN (n_2540), .A1 (B_imm[8]), .A2 (A_imm[8]));
OAI21_X1 i_2603 (.ZN (n_2539), .A (n_2540), .B1 (n_2542), .B2 (n_2549));
AOI22_X1 i_2602 (.ZN (n_2538), .A1 (n_2550), .A2 (n_2557), .B1 (n_2539), .B2 (n_2541));
INV_X1 i_2601 (.ZN (n_2537), .A (n_2538));
NAND4_X1 i_2600 (.ZN (n_2536), .A1 (n_2550), .A2 (n_2539), .A3 (n_2557), .A4 (n_2541));
OAI22_X1 i_2599 (.ZN (n_2535), .A1 (n_8829), .A2 (n_6836), .B1 (n_8347), .B2 (n_8644));
NAND2_X1 i_2598 (.ZN (n_2534), .A1 (B_imm[13]), .A2 (A_imm[3]));
INV_X1 i_2597 (.ZN (n_2533), .A (n_2534));
NAND4_X1 i_2596 (.ZN (n_2532), .A1 (B_imm[15]), .A2 (B_imm[9]), .A3 (A_imm[7]), .A4 (A_imm[1]));
INV_X1 i_2595 (.ZN (n_2531), .A (n_2532));
OAI21_X1 i_2594 (.ZN (n_2530), .A (n_2535), .B1 (n_2531), .B2 (n_2533));
NAND2_X1 i_2593 (.ZN (n_2529), .A1 (n_2536), .A2 (n_2530));
NAND2_X1 i_2592 (.ZN (n_2528), .A1 (n_2529), .A2 (n_2537));
OAI21_X1 i_2591 (.ZN (n_2527), .A (n_2563), .B1 (n_2559), .B2 (n_2528));
NAND3_X1 i_2590 (.ZN (n_2526), .A1 (n_2833), .A2 (n_2831), .A3 (n_2820));
INV_X1 i_2589 (.ZN (n_2525), .A (n_2820));
NAND2_X1 i_2588 (.ZN (n_2524), .A1 (n_2833), .A2 (n_2831));
NAND2_X1 i_2587 (.ZN (n_2523), .A1 (n_2524), .A2 (n_2525));
NAND2_X1 i_2586 (.ZN (n_2522), .A1 (n_2523), .A2 (n_2526));
NAND2_X1 i_2585 (.ZN (n_2521), .A1 (n_2522), .A2 (n_2527));
INV_X1 i_2584 (.ZN (n_2520), .A (n_2528));
NAND2_X1 i_2583 (.ZN (n_2519), .A1 (n_2520), .A2 (n_2560));
NAND4_X1 i_2582 (.ZN (n_2518), .A1 (n_2523), .A2 (n_2519), .A3 (n_2563), .A4 (n_2526));
INV_X1 i_2581 (.ZN (n_2517), .A (n_2825));
OAI21_X1 i_2580 (.ZN (n_2516), .A (n_2823), .B1 (n_2517), .B2 (n_2821));
NAND3_X1 i_2579 (.ZN (n_2515), .A1 (n_2825), .A2 (n_2824), .A3 (n_2822));
NAND2_X1 i_2578 (.ZN (n_2514), .A1 (n_2516), .A2 (n_2515));
INV_X1 i_2577 (.ZN (n_2513), .A (n_2829));
NAND2_X1 i_2576 (.ZN (n_2512), .A1 (n_2830), .A2 (n_2828));
NAND2_X1 i_2575 (.ZN (n_2511), .A1 (n_2512), .A2 (n_2513));
NAND3_X1 i_2574 (.ZN (n_2510), .A1 (n_2830), .A2 (n_2829), .A3 (n_2828));
NAND2_X1 i_2573 (.ZN (n_2509), .A1 (n_2511), .A2 (n_2510));
NAND2_X1 i_2572 (.ZN (n_2508), .A1 (n_2873), .A2 (n_2871));
NAND3_X1 i_2571 (.ZN (n_2507), .A1 (n_2508), .A2 (B_imm[7]), .A3 (A_imm[10]));
NAND3_X1 i_2570 (.ZN (n_2506), .A1 (n_2873), .A2 (n_2872), .A3 (n_2871));
NAND2_X1 i_2569 (.ZN (n_2505), .A1 (n_2507), .A2 (n_2506));
NAND2_X1 i_2568 (.ZN (n_2504), .A1 (n_2509), .A2 (n_2505));
NAND4_X1 i_2567 (.ZN (n_2503), .A1 (n_2511), .A2 (n_2507), .A3 (n_2510), .A4 (n_2506));
NAND3_X1 i_2566 (.ZN (n_2502), .A1 (n_2503), .A2 (B_imm[14]), .A3 (A_imm[3]));
NAND2_X1 i_2565 (.ZN (n_2501), .A1 (n_2502), .A2 (n_2504));
NAND2_X1 i_2564 (.ZN (n_2500), .A1 (n_2501), .A2 (n_2514));
NAND4_X1 i_2563 (.ZN (n_2499), .A1 (n_2502), .A2 (n_2516), .A3 (n_2515), .A4 (n_2504));
INV_X1 i_2562 (.ZN (n_2498), .A (n_2499));
NAND2_X1 i_2561 (.ZN (n_2497), .A1 (n_2732), .A2 (n_2718));
NAND2_X1 i_2560 (.ZN (n_2496), .A1 (n_2497), .A2 (n_2720));
INV_X1 i_2559 (.ZN (n_2495), .A (n_2720));
NAND3_X1 i_2558 (.ZN (n_2494), .A1 (n_2732), .A2 (n_2495), .A3 (n_2718));
NAND2_X1 i_2557 (.ZN (n_2493), .A1 (n_2496), .A2 (n_2494));
OAI21_X1 i_2556 (.ZN (n_2492), .A (n_2500), .B1 (n_2493), .B2 (n_2498));
NAND2_X1 i_2555 (.ZN (n_2491), .A1 (n_2518), .A2 (n_2492));
NAND2_X1 i_2554 (.ZN (n_2490), .A1 (n_2491), .A2 (n_2521));
NAND2_X1 i_2553 (.ZN (n_2489), .A1 (n_2573), .A2 (n_2490));
NAND2_X1 i_2552 (.ZN (n_2488), .A1 (n_2489), .A2 (n_2574));
NAND2_X1 i_2551 (.ZN (n_2487), .A1 (n_2488), .A2 (n_2616));
NAND4_X1 i_2550 (.ZN (n_2486), .A1 (n_2489), .A2 (n_2619), .A3 (n_2617), .A4 (n_2574));
OAI211_X1 i_2549 (.ZN (n_2485), .A (n_2805), .B (n_2803), .C1 (n_2798), .C2 (n_2797));
NAND2_X1 i_2548 (.ZN (n_2484), .A1 (n_2805), .A2 (n_2803));
NAND2_X1 i_2547 (.ZN (n_2483), .A1 (n_2484), .A2 (n_2796));
NAND2_X1 i_2546 (.ZN (n_2482), .A1 (n_2485), .A2 (n_2483));
INV_X1 i_2545 (.ZN (n_2481), .A (n_2482));
NAND2_X1 i_2544 (.ZN (n_2480), .A1 (n_2486), .A2 (n_2481));
NAND2_X1 i_2543 (.ZN (n_2479), .A1 (n_2480), .A2 (n_2487));
NAND2_X1 i_2542 (.ZN (n_2478), .A1 (n_2479), .A2 (n_2625));
OAI211_X1 i_2541 (.ZN (n_2477), .A (n_2480), .B (n_2487), .C1 (n_2627), .C2 (n_2626));
OAI211_X1 i_2540 (.ZN (n_2476), .A (n_2654), .B (n_2653), .C1 (n_2651), .C2 (n_2650));
NAND2_X1 i_2539 (.ZN (n_2475), .A1 (n_2654), .A2 (n_2653));
NAND2_X1 i_2538 (.ZN (n_2474), .A1 (n_2475), .A2 (n_2649));
NAND4_X1 i_2537 (.ZN (n_2473), .A1 (n_2478), .A2 (n_2477), .A3 (n_2474), .A4 (n_2476));
NAND2_X1 i_2536 (.ZN (n_2472), .A1 (n_2478), .A2 (n_2477));
NAND2_X1 i_2535 (.ZN (n_2471), .A1 (n_2476), .A2 (n_2474));
NAND2_X1 i_2534 (.ZN (n_2470), .A1 (n_2472), .A2 (n_2471));
NAND2_X1 i_2533 (.ZN (n_2469), .A1 (n_2470), .A2 (n_2473));
NAND3_X1 i_2532 (.ZN (n_2468), .A1 (n_2674), .A2 (n_2672), .A3 (n_2657));
NAND2_X1 i_2531 (.ZN (n_2467), .A1 (n_2674), .A2 (n_2672));
NAND3_X1 i_2530 (.ZN (n_2466), .A1 (n_2467), .A2 (n_2664), .A3 (n_2658));
NAND3_X1 i_2529 (.ZN (n_2465), .A1 (n_2716), .A2 (n_2741), .A3 (n_2744));
NAND2_X1 i_2528 (.ZN (n_2464), .A1 (n_2741), .A2 (n_2744));
NAND3_X1 i_2527 (.ZN (n_2463), .A1 (n_2464), .A2 (n_2732), .A3 (n_2717));
NAND2_X1 i_2526 (.ZN (n_2462), .A1 (n_2463), .A2 (n_2465));
INV_X1 i_2525 (.ZN (n_2461), .A (n_2462));
INV_X1 i_2524 (.ZN (n_2460), .A (n_2683));
OAI21_X1 i_2523 (.ZN (n_2459), .A (n_2680), .B1 (n_2460), .B2 (n_2682));
NAND2_X1 i_2522 (.ZN (n_2458), .A1 (n_2688), .A2 (n_2691));
NAND3_X1 i_2521 (.ZN (n_2457), .A1 (n_2458), .A2 (n_2686), .A3 (n_2685));
INV_X1 i_2520 (.ZN (n_2456), .A (n_2680));
NAND3_X1 i_2519 (.ZN (n_2455), .A1 (n_2457), .A2 (n_2683), .A3 (n_2456));
NAND2_X1 i_2518 (.ZN (n_2454), .A1 (n_2731), .A2 (n_2722));
NAND2_X1 i_2517 (.ZN (n_2453), .A1 (n_2454), .A2 (n_2723));
NAND3_X1 i_2516 (.ZN (n_2452), .A1 (n_2731), .A2 (n_2724), .A3 (n_2722));
NAND2_X1 i_2515 (.ZN (n_2451), .A1 (n_2453), .A2 (n_2452));
INV_X1 i_2514 (.ZN (n_2450), .A (n_2739));
NAND2_X1 i_2513 (.ZN (n_2449), .A1 (n_2740), .A2 (n_2738));
NAND2_X1 i_2512 (.ZN (n_2448), .A1 (n_2449), .A2 (n_2450));
NAND3_X1 i_2511 (.ZN (n_2447), .A1 (n_2740), .A2 (n_2739), .A3 (n_2738));
NAND2_X1 i_2510 (.ZN (n_2446), .A1 (n_2448), .A2 (n_2447));
NAND2_X1 i_2509 (.ZN (n_2445), .A1 (n_2446), .A2 (n_2451));
NAND4_X1 i_2508 (.ZN (n_2444), .A1 (n_2448), .A2 (n_2453), .A3 (n_2452), .A4 (n_2447));
INV_X1 i_2507 (.ZN (n_2443), .A (n_2444));
OAI22_X1 i_2506 (.ZN (n_2442), .A1 (n_8752), .A2 (n_6817), .B1 (n_8751), .B2 (n_8429));
NAND2_X1 i_2505 (.ZN (n_2441), .A1 (B_imm[6]), .A2 (A_imm[9]));
NAND4_X1 i_2504 (.ZN (n_2440), .A1 (A_imm[12]), .A2 (B_imm[5]), .A3 (B_imm[3]), .A4 (A_imm[10]));
NAND2_X1 i_2503 (.ZN (n_2439), .A1 (n_2440), .A2 (n_2441));
AOI21_X1 i_2502 (.ZN (n_2438), .A (n_2728), .B1 (n_2729), .B2 (n_2726));
INV_X1 i_2501 (.ZN (n_2437), .A (n_2438));
NAND3_X1 i_2500 (.ZN (n_2436), .A1 (n_2729), .A2 (n_2728), .A3 (n_2726));
NAND2_X1 i_2499 (.ZN (n_2435), .A1 (n_2437), .A2 (n_2436));
NAND3_X1 i_2498 (.ZN (n_2434), .A1 (n_2435), .A2 (n_2442), .A3 (n_2439));
INV_X1 i_2497 (.ZN (n_2433), .A (n_2434));
NAND2_X1 i_2496 (.ZN (n_2432), .A1 (n_2439), .A2 (n_2442));
NAND3_X1 i_2495 (.ZN (n_2431), .A1 (n_2432), .A2 (n_2437), .A3 (n_2436));
OAI22_X1 i_2494 (.ZN (n_2430), .A1 (n_8849), .A2 (n_6678), .B1 (n_8795), .B2 (n_3718));
NAND2_X1 i_2493 (.ZN (n_2429), .A1 (B_imm[9]), .A2 (A_imm[6]));
INV_X1 i_2492 (.ZN (n_2428), .A (n_2429));
NAND4_X1 i_2491 (.ZN (n_2427), .A1 (B_imm[11]), .A2 (B_imm[12]), .A3 (A_imm[4]), .A4 (A_imm[3]));
INV_X1 i_2490 (.ZN (n_2426), .A (n_2427));
OAI21_X1 i_2489 (.ZN (n_2425), .A (n_2430), .B1 (n_2428), .B2 (n_2426));
INV_X1 i_2488 (.ZN (n_2424), .A (n_2425));
AOI21_X1 i_2487 (.ZN (n_2423), .A (n_2433), .B1 (n_2424), .B2 (n_2431));
OAI21_X1 i_2486 (.ZN (n_2422), .A (n_2445), .B1 (n_2423), .B2 (n_2443));
NAND3_X1 i_2485 (.ZN (n_2421), .A1 (n_2422), .A2 (n_2459), .A3 (n_2455));
NAND2_X1 i_2484 (.ZN (n_2420), .A1 (n_2459), .A2 (n_2455));
INV_X1 i_2483 (.ZN (n_2419), .A (n_2422));
NAND2_X1 i_2482 (.ZN (n_2418), .A1 (n_2420), .A2 (n_2419));
NAND4_X1 i_2481 (.ZN (n_2417), .A1 (n_2595), .A2 (n_2594), .A3 (n_2591), .A4 (n_2590));
OAI21_X1 i_2480 (.ZN (n_2416), .A (n_2589), .B1 (n_2593), .B2 (n_2596));
NAND2_X1 i_2479 (.ZN (n_2415), .A1 (n_2417), .A2 (n_2416));
NAND2_X1 i_2478 (.ZN (n_2414), .A1 (n_2691), .A2 (n_2689));
NAND3_X1 i_2477 (.ZN (n_2413), .A1 (n_2414), .A2 (B_imm[15]), .A3 (A_imm[2]));
NAND3_X1 i_2476 (.ZN (n_2412), .A1 (n_2691), .A2 (n_2690), .A3 (n_2689));
NAND2_X1 i_2475 (.ZN (n_2411), .A1 (n_2413), .A2 (n_2412));
NAND2_X1 i_2474 (.ZN (n_2410), .A1 (n_2415), .A2 (n_2411));
NAND4_X2 i_2473 (.ZN (n_2409), .A1 (n_2413), .A2 (n_2416), .A3 (n_2417), .A4 (n_2412));
INV_X1 i_2472 (.ZN (n_2408), .A (n_2409));
OAI22_X1 i_2471 (.ZN (n_2407), .A1 (n_8880), .A2 (n_6678), .B1 (n_8926), .B2 (n_6817));
NAND2_X1 i_2470 (.ZN (n_2406), .A1 (B_imm[7]), .A2 (A_imm[7]));
NAND4_X1 i_2469 (.ZN (n_2405), .A1 (B_imm[10]), .A2 (A_imm[11]), .A3 (B_imm[3]), .A4 (A_imm[4]));
NAND2_X1 i_2468 (.ZN (n_2404), .A1 (n_2405), .A2 (n_2406));
NAND2_X1 i_2467 (.ZN (n_2403), .A1 (n_2404), .A2 (n_2407));
OAI21_X2 i_2466 (.ZN (n_2402), .A (n_2403), .B1 (n_8947), .B2 (n_8644));
NAND4_X1 i_2465 (.ZN (n_2401), .A1 (n_2404), .A2 (n_2407), .A3 (B_imm[8]), .A4 (A_imm[7]));
INV_X1 i_2464 (.ZN (n_2400), .A (n_2401));
OAI22_X1 i_2463 (.ZN (n_2399), .A1 (n_8645), .A2 (n_8429), .B1 (n_8971), .B2 (n_6740));
NAND2_X1 i_2462 (.ZN (n_2398), .A1 (A_imm[13]), .A2 (B_imm[1]));
INV_X1 i_2461 (.ZN (n_2397), .A (n_2398));
NAND4_X1 i_2460 (.ZN (n_2396), .A1 (A_imm[9]), .A2 (A_imm[14]), .A3 (B_imm[5]), .A4 (B_imm[0]));
INV_X1 i_2459 (.ZN (n_2395), .A (n_2396));
OAI21_X1 i_2458 (.ZN (n_2394), .A (n_2399), .B1 (n_2395), .B2 (n_2397));
INV_X1 i_2457 (.ZN (n_2393), .A (n_2394));
OAI21_X1 i_2456 (.ZN (n_2392), .A (n_2402), .B1 (n_2393), .B2 (n_2400));
INV_X1 i_2455 (.ZN (n_2391), .A (n_2392));
AOI21_X1 i_2454 (.ZN (n_2390), .A (n_2695), .B1 (n_2696), .B2 (n_2694));
NAND3_X1 i_2453 (.ZN (n_2389), .A1 (n_2696), .A2 (n_2695), .A3 (n_2694));
INV_X1 i_2452 (.ZN (n_2388), .A (n_2389));
NOR2_X1 i_2451 (.ZN (n_2387), .A1 (n_2390), .A2 (n_2388));
INV_X1 i_2450 (.ZN (n_2386), .A (n_2387));
NAND2_X1 i_2449 (.ZN (n_2385), .A1 (n_2391), .A2 (n_2386));
NAND2_X1 i_2448 (.ZN (n_2384), .A1 (n_2392), .A2 (n_2387));
INV_X1 i_2447 (.ZN (n_2383), .A (n_2599));
NAND2_X1 i_2446 (.ZN (n_2382), .A1 (n_2600), .A2 (n_2598));
NAND2_X1 i_2445 (.ZN (n_2381), .A1 (n_2382), .A2 (n_2383));
NAND3_X1 i_2444 (.ZN (n_2380), .A1 (n_2600), .A2 (n_2599), .A3 (n_2598));
NAND2_X1 i_2443 (.ZN (n_2379), .A1 (n_2381), .A2 (n_2380));
NAND2_X1 i_2442 (.ZN (n_2378), .A1 (n_2384), .A2 (n_2379));
NAND2_X1 i_2441 (.ZN (n_2377), .A1 (n_2378), .A2 (n_2385));
INV_X1 i_2440 (.ZN (n_2376), .A (n_2377));
OAI21_X1 i_2439 (.ZN (n_2375), .A (n_2410), .B1 (n_2408), .B2 (n_2376));
NAND2_X2 i_2438 (.ZN (n_2374), .A1 (n_2418), .A2 (n_2375));
AOI21_X2 i_2437 (.ZN (n_2373), .A (n_2461), .B1 (n_2374), .B2 (n_2421));
INV_X2 i_2436 (.ZN (n_2372), .A (n_2373));
NAND3_X2 i_2435 (.ZN (n_2371), .A1 (n_2374), .A2 (n_2461), .A3 (n_2421));
NAND3_X1 i_2434 (.ZN (n_2370), .A1 (n_2699), .A2 (n_2697), .A3 (n_2679));
INV_X1 i_2433 (.ZN (n_2369), .A (n_2679));
NAND2_X1 i_2432 (.ZN (n_2368), .A1 (n_2699), .A2 (n_2697));
NAND2_X1 i_2431 (.ZN (n_2367), .A1 (n_2368), .A2 (n_2369));
NAND2_X1 i_2430 (.ZN (n_2366), .A1 (n_2367), .A2 (n_2370));
INV_X1 i_2429 (.ZN (n_2365), .A (n_2366));
NAND2_X1 i_2428 (.ZN (n_2364), .A1 (n_2371), .A2 (n_2365));
NAND2_X1 i_2427 (.ZN (n_2363), .A1 (n_2364), .A2 (n_2372));
NAND3_X1 i_2426 (.ZN (n_2362), .A1 (n_2677), .A2 (n_2711), .A3 (n_2707));
NAND2_X1 i_2425 (.ZN (n_2361), .A1 (n_2711), .A2 (n_2707));
NAND3_X1 i_2424 (.ZN (n_2360), .A1 (n_2361), .A2 (n_2699), .A3 (n_2678));
NAND2_X1 i_2423 (.ZN (n_2359), .A1 (n_2360), .A2 (n_2362));
INV_X1 i_2422 (.ZN (n_2358), .A (n_2359));
NAND2_X1 i_2421 (.ZN (n_2357), .A1 (n_2363), .A2 (n_2358));
NAND3_X1 i_2420 (.ZN (n_2356), .A1 (n_2364), .A2 (n_2372), .A3 (n_2359));
NAND2_X1 i_2419 (.ZN (n_2355), .A1 (n_2659), .A2 (n_2661));
NAND3_X1 i_2418 (.ZN (n_2354), .A1 (n_2355), .A2 (n_2662), .A3 (n_2664));
NAND2_X1 i_2417 (.ZN (n_2353), .A1 (n_2662), .A2 (n_2664));
NAND3_X1 i_2416 (.ZN (n_2352), .A1 (n_2353), .A2 (n_2661), .A3 (n_2659));
NAND2_X1 i_2415 (.ZN (n_2351), .A1 (n_2352), .A2 (n_2354));
NAND2_X1 i_2414 (.ZN (n_2350), .A1 (n_2356), .A2 (n_2351));
NAND2_X1 i_2413 (.ZN (n_2349), .A1 (n_2350), .A2 (n_2357));
NAND3_X1 i_2412 (.ZN (n_2348), .A1 (n_2349), .A2 (n_2468), .A3 (n_2466));
NAND2_X1 i_2411 (.ZN (n_2347), .A1 (n_2466), .A2 (n_2468));
NAND3_X1 i_2410 (.ZN (n_2346), .A1 (n_2347), .A2 (n_2357), .A3 (n_2350));
NAND3_X1 i_2409 (.ZN (n_2345), .A1 (n_2487), .A2 (n_2486), .A3 (n_2482));
NAND2_X1 i_2408 (.ZN (n_2344), .A1 (n_2487), .A2 (n_2486));
NAND2_X1 i_2407 (.ZN (n_2343), .A1 (n_2344), .A2 (n_2481));
NAND2_X1 i_2406 (.ZN (n_2342), .A1 (n_2343), .A2 (n_2345));
NAND2_X1 i_2405 (.ZN (n_2341), .A1 (n_2342), .A2 (n_2346));
NAND2_X1 i_2404 (.ZN (n_2340), .A1 (n_2341), .A2 (n_2348));
NAND2_X1 i_2403 (.ZN (n_2339), .A1 (n_2469), .A2 (n_2340));
NAND3_X1 i_2402 (.ZN (n_2338), .A1 (n_2638), .A2 (n_2646), .A3 (n_2644));
NAND2_X1 i_2401 (.ZN (n_2337), .A1 (n_2644), .A2 (n_2646));
NAND3_X2 i_2400 (.ZN (n_2336), .A1 (n_2337), .A2 (n_2642), .A3 (n_2639));
NAND2_X1 i_2399 (.ZN (n_2335), .A1 (n_2471), .A2 (n_2477));
NAND2_X1 i_2398 (.ZN (n_2334), .A1 (n_2335), .A2 (n_2478));
NAND3_X2 i_2397 (.ZN (n_2333), .A1 (n_2334), .A2 (n_2336), .A3 (n_2338));
NAND2_X1 i_2396 (.ZN (n_2332), .A1 (n_2336), .A2 (n_2338));
INV_X1 i_2395 (.ZN (n_2331), .A (n_2334));
NAND2_X1 i_2394 (.ZN (n_2330), .A1 (n_2332), .A2 (n_2331));
NAND2_X2 i_2393 (.ZN (n_2329), .A1 (n_2330), .A2 (n_2333));
NAND2_X2 i_2392 (.ZN (n_2328), .A1 (n_2329), .A2 (n_2339));
NAND3_X1 i_2391 (.ZN (n_2327), .A1 (n_2765), .A2 (n_2637), .A3 (n_2768));
OAI21_X2 i_2389 (.ZN (n_2325), .A (n_2333), .B1 (CLOCK_opt_ipo_n423), .B2 (n_2636));
NAND2_X1 i_2388 (.ZN (n_2324), .A1 (n_2325), .A2 (n_2328));
INV_X1 i_2387 (.ZN (n_2323), .A (n_2324));
NAND3_X1 i_2386 (.ZN (n_2322), .A1 (n_2342), .A2 (n_2348), .A3 (n_2346));
INV_X1 i_2385 (.ZN (n_2321), .A (n_2342));
NAND2_X1 i_2384 (.ZN (n_2320), .A1 (n_2348), .A2 (n_2346));
NAND2_X1 i_2383 (.ZN (n_2319), .A1 (n_2320), .A2 (n_2321));
NAND3_X1 i_2382 (.ZN (n_2318), .A1 (n_2601), .A2 (n_2603), .A3 (n_2588));
INV_X1 i_2381 (.ZN (n_2317), .A (n_2318));
AOI21_X1 i_2380 (.ZN (n_2316), .A (n_2588), .B1 (n_2601), .B2 (n_2603));
NOR2_X1 i_2379 (.ZN (n_2315), .A1 (n_2317), .A2 (n_2316));
INV_X1 i_2378 (.ZN (n_2314), .A (n_2536));
INV_X1 i_2377 (.ZN (n_2313), .A (n_2530));
OAI21_X1 i_2376 (.ZN (n_2312), .A (n_2313), .B1 (n_2314), .B2 (n_2538));
NAND3_X1 i_2375 (.ZN (n_2311), .A1 (n_2537), .A2 (n_2536), .A3 (n_2530));
NAND2_X1 i_2374 (.ZN (n_2310), .A1 (n_2312), .A2 (n_2311));
INV_X1 i_2373 (.ZN (n_2309), .A (n_2540));
INV_X1 i_2372 (.ZN (n_2308), .A (n_2542));
NAND3_X1 i_2371 (.ZN (n_2307), .A1 (n_2308), .A2 (B_imm[0]), .A3 (A_imm[16]));
NAND2_X1 i_2370 (.ZN (n_2306), .A1 (n_2307), .A2 (n_2541));
NAND2_X1 i_2369 (.ZN (n_2305), .A1 (n_2306), .A2 (n_2309));
NAND3_X1 i_2368 (.ZN (n_2304), .A1 (n_2307), .A2 (n_2541), .A3 (n_2540));
NAND2_X1 i_2367 (.ZN (n_2303), .A1 (n_2305), .A2 (n_2304));
NAND3_X1 i_2366 (.ZN (n_2302), .A1 (n_2303), .A2 (B_imm[14]), .A3 (A_imm[2]));
NAND2_X1 i_2365 (.ZN (n_2301), .A1 (B_imm[14]), .A2 (A_imm[2]));
NAND3_X1 i_2364 (.ZN (n_2300), .A1 (n_2301), .A2 (n_2305), .A3 (n_2304));
NAND4_X1 i_2363 (.ZN (n_2299), .A1 (B_imm[13]), .A2 (B_imm[15]), .A3 (A_imm[2]), .A4 (A_imm[0]));
NAND2_X1 i_2362 (.ZN (n_2298), .A1 (B_imm[15]), .A2 (A_imm[0]));
OAI21_X1 i_2361 (.ZN (n_2297), .A (n_2298), .B1 (n_8973), .B2 (n_6677));
INV_X1 i_2360 (.ZN (n_2296), .A (n_2297));
NAND2_X1 i_2359 (.ZN (n_2295), .A1 (n_2547), .A2 (n_2544));
XNOR2_X1 i_2358 (.ZN (n_2294), .A (n_2295), .B (n_2546));
OAI21_X1 i_2357 (.ZN (n_2293), .A (n_2299), .B1 (n_2296), .B2 (n_2294));
NAND2_X1 i_2356 (.ZN (n_2292), .A1 (n_2300), .A2 (n_2293));
NAND2_X1 i_2355 (.ZN (n_2291), .A1 (n_2302), .A2 (n_2292));
NAND2_X1 i_2354 (.ZN (n_2290), .A1 (n_2291), .A2 (n_2310));
NAND4_X1 i_2353 (.ZN (n_2289), .A1 (n_2292), .A2 (n_2312), .A3 (n_2311), .A4 (n_2302));
INV_X1 i_2352 (.ZN (n_2288), .A (n_2552));
NAND2_X1 i_2351 (.ZN (n_2287), .A1 (n_2557), .A2 (n_2551));
NAND2_X1 i_2350 (.ZN (n_2286), .A1 (n_2287), .A2 (n_2288));
NAND3_X1 i_2349 (.ZN (n_2285), .A1 (n_2557), .A2 (n_2552), .A3 (n_2551));
NAND2_X1 i_2348 (.ZN (n_2284), .A1 (n_2286), .A2 (n_2285));
OAI22_X1 i_2347 (.ZN (n_2283), .A1 (n_8849), .A2 (n_3718), .B1 (n_8795), .B2 (n_6677));
NAND2_X1 i_2346 (.ZN (n_2282), .A1 (B_imm[9]), .A2 (A_imm[5]));
NAND4_X1 i_2345 (.ZN (n_2281), .A1 (B_imm[11]), .A2 (B_imm[12]), .A3 (A_imm[3]), .A4 (A_imm[2]));
NAND2_X1 i_2344 (.ZN (n_2280), .A1 (n_2281), .A2 (n_2282));
AOI22_X1 i_2343 (.ZN (n_2279), .A1 (A_imm[12]), .A2 (B_imm[2]), .B1 (A_imm[10]), .B2 (B_imm[4]));
OAI22_X1 i_2342 (.ZN (n_2278), .A1 (n_6584), .A2 (n_8926), .B1 (n_8429), .B2 (n_8511));
NAND2_X1 i_2341 (.ZN (n_2277), .A1 (B_imm[10]), .A2 (A_imm[3]));
INV_X1 i_2340 (.ZN (n_2276), .A (n_2277));
NAND4_X1 i_2339 (.ZN (n_2275), .A1 (A_imm[11]), .A2 (B_imm[5]), .A3 (B_imm[2]), .A4 (A_imm[8]));
INV_X1 i_2338 (.ZN (n_2274), .A (n_2275));
OAI21_X1 i_2337 (.ZN (n_2273), .A (n_2278), .B1 (n_2276), .B2 (n_2274));
NAND4_X1 i_2336 (.ZN (n_2272), .A1 (A_imm[12]), .A2 (B_imm[4]), .A3 (B_imm[2]), .A4 (A_imm[10]));
AOI21_X1 i_2335 (.ZN (n_2271), .A (n_2279), .B1 (n_2273), .B2 (n_2272));
AOI21_X1 i_2334 (.ZN (n_2270), .A (n_2271), .B1 (n_2283), .B2 (n_2280));
INV_X1 i_2333 (.ZN (n_2269), .A (n_2270));
NAND3_X1 i_2332 (.ZN (n_2268), .A1 (n_2271), .A2 (n_2280), .A3 (n_2283));
NAND2_X1 i_2331 (.ZN (n_2267), .A1 (n_2556), .A2 (n_2554));
NAND3_X1 i_2330 (.ZN (n_2266), .A1 (n_2267), .A2 (B_imm[0]), .A3 (A_imm[15]));
NAND3_X1 i_2329 (.ZN (n_2265), .A1 (n_2556), .A2 (n_2555), .A3 (n_2554));
NAND2_X1 i_2328 (.ZN (n_2264), .A1 (n_2266), .A2 (n_2265));
INV_X1 i_2327 (.ZN (n_2263), .A (n_2264));
NAND2_X1 i_2326 (.ZN (n_2262), .A1 (n_2268), .A2 (n_2263));
NAND3_X1 i_2325 (.ZN (n_2261), .A1 (n_2262), .A2 (n_2284), .A3 (n_2269));
AOI21_X1 i_2324 (.ZN (n_2260), .A (n_2284), .B1 (n_2269), .B2 (n_2262));
AOI21_X1 i_2323 (.ZN (n_2259), .A (n_2534), .B1 (n_2535), .B2 (n_2532));
NAND3_X1 i_2322 (.ZN (n_2258), .A1 (n_2535), .A2 (n_2534), .A3 (n_2532));
INV_X1 i_2321 (.ZN (n_2257), .A (n_2258));
NOR2_X1 i_2320 (.ZN (n_2256), .A1 (n_2259), .A2 (n_2257));
OAI21_X2 i_2319 (.ZN (n_2255), .A (n_2261), .B1 (n_2260), .B2 (n_2256));
NAND2_X2 i_2318 (.ZN (n_2254), .A1 (n_2255), .A2 (n_2289));
AOI21_X2 i_2317 (.ZN (n_2253), .A (n_2315), .B1 (n_2254), .B2 (n_2290));
INV_X1 i_2316 (.ZN (n_2252), .A (n_2253));
NAND3_X1 i_2315 (.ZN (n_2251), .A1 (n_2254), .A2 (n_2315), .A3 (n_2290));
NAND2_X1 i_2314 (.ZN (n_2250), .A1 (n_2560), .A2 (n_2563));
XNOR2_X1 i_2313 (.ZN (n_2249), .A (n_2250), .B (n_2520));
NAND2_X1 i_2312 (.ZN (n_2248), .A1 (n_2251), .A2 (n_2249));
NAND3_X1 i_2311 (.ZN (n_2247), .A1 (n_2584), .A2 (n_2577), .A3 (n_2583));
NAND2_X1 i_2310 (.ZN (n_2246), .A1 (n_2584), .A2 (n_2583));
NAND2_X1 i_2309 (.ZN (n_2245), .A1 (n_2246), .A2 (n_2578));
NAND2_X1 i_2308 (.ZN (n_2244), .A1 (n_2245), .A2 (n_2247));
AOI21_X1 i_2307 (.ZN (n_2243), .A (n_2244), .B1 (n_2252), .B2 (n_2248));
INV_X1 i_2306 (.ZN (n_2242), .A (n_2243));
NAND3_X1 i_2305 (.ZN (n_2241), .A1 (n_2248), .A2 (n_2252), .A3 (n_2244));
NAND3_X1 i_2304 (.ZN (n_2240), .A1 (n_2521), .A2 (n_2518), .A3 (n_2492));
INV_X1 i_2303 (.ZN (n_2239), .A (n_2492));
NAND2_X1 i_2302 (.ZN (n_2238), .A1 (n_2521), .A2 (n_2518));
NAND2_X1 i_2301 (.ZN (n_2237), .A1 (n_2238), .A2 (n_2239));
NAND2_X1 i_2300 (.ZN (n_2236), .A1 (n_2237), .A2 (n_2240));
INV_X1 i_2299 (.ZN (n_2235), .A (n_2236));
NAND2_X1 i_2298 (.ZN (n_2234), .A1 (n_2241), .A2 (n_2235));
NAND2_X1 i_2297 (.ZN (n_2233), .A1 (n_2242), .A2 (n_2234));
NAND3_X1 i_2296 (.ZN (n_2232), .A1 (n_2574), .A2 (n_2573), .A3 (n_2490));
NAND2_X1 i_2295 (.ZN (n_2231), .A1 (n_2574), .A2 (n_2573));
NAND3_X1 i_2294 (.ZN (n_2230), .A1 (n_2231), .A2 (n_2521), .A3 (n_2491));
NAND2_X1 i_2293 (.ZN (n_2229), .A1 (n_2230), .A2 (n_2232));
INV_X1 i_2292 (.ZN (n_2228), .A (n_2229));
NAND2_X1 i_2291 (.ZN (n_2227), .A1 (n_2233), .A2 (n_2228));
NAND3_X1 i_2290 (.ZN (n_2226), .A1 (n_2229), .A2 (n_2234), .A3 (n_2242));
NAND3_X1 i_2289 (.ZN (n_2225), .A1 (n_2357), .A2 (n_2356), .A3 (n_2351));
AOI21_X1 i_2288 (.ZN (n_2224), .A (n_2359), .B1 (n_2372), .B2 (n_2364));
INV_X1 i_2287 (.ZN (n_2223), .A (n_2356));
INV_X1 i_2286 (.ZN (n_2222), .A (n_2351));
OAI21_X1 i_2285 (.ZN (n_2221), .A (n_2222), .B1 (n_2223), .B2 (n_2224));
NAND3_X1 i_2284 (.ZN (n_2220), .A1 (n_2226), .A2 (n_2225), .A3 (n_2221));
NAND2_X1 i_2283 (.ZN (n_2219), .A1 (n_2220), .A2 (n_2227));
NAND3_X1 i_2282 (.ZN (n_2218), .A1 (n_2319), .A2 (n_2322), .A3 (n_2219));
INV_X1 i_2281 (.ZN (n_2217), .A (n_2218));
NAND4_X1 i_2280 (.ZN (n_2216), .A1 (n_2470), .A2 (n_2473), .A3 (n_2348), .A4 (n_2341));
AOI21_X2 i_2279 (.ZN (n_2215), .A (n_2217), .B1 (n_2339), .B2 (n_2216));
NAND2_X1 i_2278 (.ZN (n_2214), .A1 (n_2319), .A2 (n_2322));
INV_X1 i_2277 (.ZN (n_2213), .A (n_2219));
NAND2_X1 i_2276 (.ZN (n_2212), .A1 (n_2214), .A2 (n_2213));
NAND2_X1 i_2275 (.ZN (n_2211), .A1 (n_2221), .A2 (n_2225));
NAND3_X1 i_2274 (.ZN (n_2210), .A1 (n_2211), .A2 (n_2227), .A3 (n_2226));
INV_X1 i_2273 (.ZN (n_2209), .A (n_2211));
NAND2_X1 i_2272 (.ZN (n_2208), .A1 (n_2227), .A2 (n_2226));
NAND2_X2 i_2271 (.ZN (n_2207), .A1 (n_2208), .A2 (n_2209));
NAND2_X1 i_2270 (.ZN (n_2206), .A1 (n_2504), .A2 (n_2503));
NAND3_X1 i_2269 (.ZN (n_2205), .A1 (n_2206), .A2 (B_imm[14]), .A3 (A_imm[3]));
OAI211_X1 i_2268 (.ZN (n_2204), .A (n_2504), .B (n_2503), .C1 (n_7913), .C2 (n_3718));
NAND2_X1 i_2267 (.ZN (n_2203), .A1 (n_2205), .A2 (n_2204));
NAND2_X1 i_2266 (.ZN (n_2202), .A1 (n_2434), .A2 (n_2431));
NAND2_X1 i_2265 (.ZN (n_2201), .A1 (n_2202), .A2 (n_2425));
NAND3_X1 i_2264 (.ZN (n_2200), .A1 (n_2424), .A2 (n_2434), .A3 (n_2431));
OAI22_X1 i_2263 (.ZN (n_2199), .A1 (n_8947), .A2 (n_7691), .B1 (n_8232), .B2 (n_8511));
OAI22_X1 i_2262 (.ZN (n_2198), .A1 (n_8645), .A2 (n_6577), .B1 (n_8573), .B2 (n_7691));
NAND2_X1 i_2261 (.ZN (n_2197), .A1 (A_imm[13]), .A2 (B_imm[0]));
INV_X1 i_2260 (.ZN (n_2196), .A (n_2197));
NAND4_X1 i_2259 (.ZN (n_2195), .A1 (A_imm[9]), .A2 (B_imm[7]), .A3 (B_imm[4]), .A4 (A_imm[6]));
INV_X1 i_2258 (.ZN (n_2194), .A (n_2195));
OAI21_X1 i_2257 (.ZN (n_2193), .A (n_2198), .B1 (n_2194), .B2 (n_2196));
INV_X1 i_2256 (.ZN (n_2192), .A (n_2193));
NAND4_X1 i_2255 (.ZN (n_2191), .A1 (B_imm[8]), .A2 (B_imm[6]), .A3 (A_imm[8]), .A4 (A_imm[6]));
INV_X1 i_2254 (.ZN (n_2190), .A (n_2191));
OAI21_X1 i_2253 (.ZN (n_2189), .A (n_2199), .B1 (n_2192), .B2 (n_2190));
INV_X1 i_2252 (.ZN (n_2188), .A (n_2189));
INV_X1 i_2251 (.ZN (n_2187), .A (n_2441));
NAND2_X1 i_2250 (.ZN (n_2186), .A1 (n_2442), .A2 (n_2440));
NAND2_X1 i_2249 (.ZN (n_2185), .A1 (n_2186), .A2 (n_2187));
NAND3_X1 i_2248 (.ZN (n_2184), .A1 (n_2442), .A2 (n_2441), .A3 (n_2440));
NAND2_X1 i_2247 (.ZN (n_2183), .A1 (n_2185), .A2 (n_2184));
NAND2_X1 i_2246 (.ZN (n_2182), .A1 (n_2188), .A2 (n_2183));
NAND3_X1 i_2245 (.ZN (n_2181), .A1 (n_2189), .A2 (n_2185), .A3 (n_2184));
NAND2_X1 i_2244 (.ZN (n_2180), .A1 (B_imm[14]), .A2 (A_imm[1]));
INV_X1 i_2243 (.ZN (n_2179), .A (n_2180));
NAND2_X1 i_2242 (.ZN (n_2178), .A1 (n_2181), .A2 (n_2179));
NAND2_X1 i_2241 (.ZN (n_2177), .A1 (n_2178), .A2 (n_2182));
NAND3_X1 i_2240 (.ZN (n_2176), .A1 (n_2177), .A2 (n_2201), .A3 (n_2200));
NAND2_X1 i_2239 (.ZN (n_2175), .A1 (n_2200), .A2 (n_2201));
NAND3_X1 i_2238 (.ZN (n_2174), .A1 (n_2175), .A2 (n_2182), .A3 (n_2178));
NAND2_X1 i_2237 (.ZN (n_2173), .A1 (B_imm[13]), .A2 (A_imm[1]));
INV_X1 i_2236 (.ZN (n_2172), .A (n_2173));
AOI22_X1 i_2235 (.ZN (n_2171), .A1 (A_imm[12]), .A2 (B_imm[1]), .B1 (A_imm[10]), .B2 (B_imm[3]));
OAI22_X1 i_2234 (.ZN (n_2170), .A1 (n_8429), .A2 (n_8644), .B1 (n_6577), .B2 (n_8511));
NAND2_X1 i_2233 (.ZN (n_2169), .A1 (A_imm[11]), .A2 (B_imm[1]));
INV_X1 i_2232 (.ZN (n_2168), .A (n_2169));
NAND4_X1 i_2231 (.ZN (n_2167), .A1 (B_imm[5]), .A2 (B_imm[4]), .A3 (A_imm[8]), .A4 (A_imm[7]));
INV_X1 i_2230 (.ZN (n_2166), .A (n_2167));
OAI21_X1 i_2229 (.ZN (n_2165), .A (n_2170), .B1 (n_2168), .B2 (n_2166));
NAND4_X1 i_2228 (.ZN (n_2164), .A1 (A_imm[12]), .A2 (B_imm[3]), .A3 (B_imm[1]), .A4 (A_imm[10]));
AOI21_X1 i_2227 (.ZN (n_2163), .A (n_2171), .B1 (n_2165), .B2 (n_2164));
NAND2_X1 i_2226 (.ZN (n_2162), .A1 (n_2163), .A2 (n_2172));
NAND2_X1 i_2225 (.ZN (n_2161), .A1 (n_2407), .A2 (n_2405));
NAND3_X1 i_2224 (.ZN (n_2160), .A1 (n_2161), .A2 (B_imm[7]), .A3 (A_imm[7]));
NAND3_X1 i_2223 (.ZN (n_2159), .A1 (n_2407), .A2 (n_2406), .A3 (n_2405));
NAND2_X1 i_2222 (.ZN (n_2158), .A1 (n_2160), .A2 (n_2159));
OAI21_X1 i_2221 (.ZN (n_2157), .A (n_2158), .B1 (n_2163), .B2 (n_2172));
NAND2_X1 i_2220 (.ZN (n_2156), .A1 (n_2157), .A2 (n_2162));
INV_X1 i_2219 (.ZN (n_2155), .A (n_2402));
OAI21_X1 i_2218 (.ZN (n_2154), .A (n_2393), .B1 (n_2155), .B2 (n_2400));
NAND3_X1 i_2217 (.ZN (n_2153), .A1 (n_2402), .A2 (n_2401), .A3 (n_2394));
NAND2_X1 i_2216 (.ZN (n_2152), .A1 (n_2154), .A2 (n_2153));
NAND2_X1 i_2215 (.ZN (n_2151), .A1 (n_2152), .A2 (n_2156));
NAND4_X1 i_2214 (.ZN (n_2150), .A1 (n_2157), .A2 (n_2154), .A3 (n_2162), .A4 (n_2153));
INV_X1 i_2213 (.ZN (n_2149), .A (n_2150));
AOI21_X1 i_2212 (.ZN (n_2148), .A (n_2429), .B1 (n_2430), .B2 (n_2427));
NAND3_X1 i_2211 (.ZN (n_2147), .A1 (n_2430), .A2 (n_2429), .A3 (n_2427));
INV_X1 i_2210 (.ZN (n_2146), .A (n_2147));
NOR2_X1 i_2209 (.ZN (n_2145), .A1 (n_2148), .A2 (n_2146));
OAI21_X1 i_2208 (.ZN (n_2144), .A (n_2151), .B1 (n_2149), .B2 (n_2145));
NAND2_X2 i_2207 (.ZN (n_2143), .A1 (n_2174), .A2 (n_2144));
NAND2_X1 i_2206 (.ZN (n_2142), .A1 (n_2143), .A2 (n_2176));
NAND2_X1 i_2205 (.ZN (n_2141), .A1 (n_2142), .A2 (n_2203));
INV_X1 i_2204 (.ZN (n_2140), .A (n_2203));
NAND3_X2 i_2203 (.ZN (n_2139), .A1 (n_2143), .A2 (n_2140), .A3 (n_2176));
INV_X1 i_2202 (.ZN (n_2138), .A (n_2423));
NAND3_X1 i_2201 (.ZN (n_2137), .A1 (n_2138), .A2 (n_2445), .A3 (n_2444));
INV_X1 i_2200 (.ZN (n_2136), .A (n_2445));
OAI21_X1 i_2199 (.ZN (n_2135), .A (n_2423), .B1 (n_2136), .B2 (n_2443));
NAND2_X1 i_2198 (.ZN (n_2134), .A1 (n_2135), .A2 (n_2137));
INV_X1 i_2197 (.ZN (n_2133), .A (n_2134));
NAND2_X1 i_2196 (.ZN (n_2132), .A1 (n_2139), .A2 (n_2133));
NAND2_X1 i_2195 (.ZN (n_2131), .A1 (n_2132), .A2 (n_2141));
NAND4_X1 i_2194 (.ZN (n_2130), .A1 (n_2500), .A2 (n_2499), .A3 (n_2496), .A4 (n_2494));
INV_X1 i_2193 (.ZN (n_2129), .A (n_2500));
OAI21_X1 i_2192 (.ZN (n_2128), .A (n_2493), .B1 (n_2129), .B2 (n_2498));
NAND3_X1 i_2191 (.ZN (n_2127), .A1 (n_2131), .A2 (n_2130), .A3 (n_2128));
NAND2_X1 i_2190 (.ZN (n_2126), .A1 (n_2128), .A2 (n_2130));
NAND3_X1 i_2189 (.ZN (n_2125), .A1 (n_2132), .A2 (n_2141), .A3 (n_2126));
NAND3_X1 i_2188 (.ZN (n_2124), .A1 (n_2418), .A2 (n_2421), .A3 (n_2375));
INV_X1 i_2187 (.ZN (n_2123), .A (n_2124));
AOI21_X1 i_2186 (.ZN (n_2122), .A (n_2375), .B1 (n_2421), .B2 (n_2418));
NOR2_X1 i_2185 (.ZN (n_2121), .A1 (n_2123), .A2 (n_2122));
NAND2_X1 i_2184 (.ZN (n_2120), .A1 (n_2125), .A2 (n_2121));
NAND2_X1 i_2183 (.ZN (n_2119), .A1 (n_2120), .A2 (n_2127));
NAND3_X1 i_2182 (.ZN (n_2118), .A1 (n_2372), .A2 (n_2371), .A3 (n_2366));
INV_X1 i_2181 (.ZN (n_2117), .A (n_2371));
OAI21_X1 i_2180 (.ZN (n_2116), .A (n_2365), .B1 (n_2117), .B2 (n_2373));
NAND2_X1 i_2179 (.ZN (n_2115), .A1 (n_2116), .A2 (n_2118));
NAND2_X1 i_2178 (.ZN (n_2114), .A1 (n_2119), .A2 (n_2115));
INV_X1 i_2177 (.ZN (n_2113), .A (n_2114));
NAND4_X1 i_2176 (.ZN (n_2112), .A1 (n_2120), .A2 (n_2116), .A3 (n_2127), .A4 (n_2118));
NAND3_X1 i_2175 (.ZN (n_2111), .A1 (n_2242), .A2 (n_2241), .A3 (n_2236));
INV_X1 i_2174 (.ZN (n_2110), .A (n_2241));
OAI21_X1 i_2173 (.ZN (n_2109), .A (n_2235), .B1 (n_2243), .B2 (n_2110));
NAND2_X1 i_2172 (.ZN (n_2108), .A1 (n_2111), .A2 (n_2109));
AOI21_X1 i_2171 (.ZN (n_2107), .A (n_2113), .B1 (n_2108), .B2 (n_2112));
AOI21_X1 i_2170 (.ZN (n_2106), .A (n_2107), .B1 (n_2210), .B2 (n_2207));
AOI21_X1 i_2169 (.ZN (n_2105), .A (n_2106), .B1 (n_2212), .B2 (n_2218));
NOR2_X4 i_2168 (.ZN (n_2104), .A1 (n_2215), .A2 (CLOCK_opt_ipo_n425));
NAND3_X1 i_2167 (.ZN (n_2103), .A1 (n_2176), .A2 (n_2174), .A3 (n_2144));
INV_X1 i_2166 (.ZN (n_2102), .A (n_2144));
NAND2_X1 i_2165 (.ZN (n_2101), .A1 (n_2174), .A2 (n_2176));
NAND2_X1 i_2164 (.ZN (n_2100), .A1 (n_2101), .A2 (n_2102));
NAND2_X1 i_2163 (.ZN (n_2099), .A1 (n_2100), .A2 (n_2103));
NAND3_X1 i_2162 (.ZN (n_2098), .A1 (n_2269), .A2 (n_2268), .A3 (n_2263));
INV_X1 i_2161 (.ZN (n_2097), .A (n_2268));
OAI21_X1 i_2160 (.ZN (n_2096), .A (n_2264), .B1 (n_2270), .B2 (n_2097));
NAND2_X1 i_2159 (.ZN (n_2095), .A1 (n_2098), .A2 (n_2096));
NAND2_X1 i_2158 (.ZN (n_2094), .A1 (n_2283), .A2 (n_2281));
NAND3_X1 i_2157 (.ZN (n_2093), .A1 (n_2094), .A2 (B_imm[9]), .A3 (A_imm[5]));
NAND3_X1 i_2156 (.ZN (n_2092), .A1 (n_2283), .A2 (n_2282), .A3 (n_2281));
NAND2_X1 i_2155 (.ZN (n_2091), .A1 (n_2093), .A2 (n_2092));
NAND2_X1 i_2154 (.ZN (n_2090), .A1 (A_imm[10]), .A2 (B_imm[2]));
OAI22_X1 i_2153 (.ZN (n_2089), .A1 (n_6577), .A2 (n_8644), .B1 (n_6817), .B2 (n_8511));
NAND2_X1 i_2152 (.ZN (n_2088), .A1 (B_imm[5]), .A2 (A_imm[6]));
NAND4_X1 i_2151 (.ZN (n_2087), .A1 (B_imm[4]), .A2 (B_imm[3]), .A3 (A_imm[8]), .A4 (A_imm[7]));
NAND2_X1 i_2150 (.ZN (n_2086), .A1 (n_2087), .A2 (n_2088));
NAND2_X1 i_2149 (.ZN (n_2085), .A1 (n_2086), .A2 (n_2089));
NAND2_X1 i_2148 (.ZN (n_2084), .A1 (n_2085), .A2 (n_2090));
NAND4_X1 i_2147 (.ZN (n_2083), .A1 (n_2086), .A2 (n_2089), .A3 (B_imm[2]), .A4 (A_imm[10]));
NAND2_X1 i_2146 (.ZN (n_2082), .A1 (A_imm[12]), .A2 (B_imm[0]));
NAND2_X1 i_2145 (.ZN (n_2081), .A1 (n_2083), .A2 (n_2082));
NAND4_X1 i_2144 (.ZN (n_2080), .A1 (n_2081), .A2 (B_imm[13]), .A3 (A_imm[0]), .A4 (n_2084));
AOI22_X1 i_2143 (.ZN (n_2079), .A1 (n_2081), .A2 (n_2084), .B1 (B_imm[13]), .B2 (A_imm[0]));
NAND2_X1 i_2142 (.ZN (n_2078), .A1 (n_2278), .A2 (n_2275));
XNOR2_X1 i_2141 (.ZN (n_2077), .A (n_2078), .B (n_2277));
OAI21_X1 i_2140 (.ZN (n_2076), .A (n_2080), .B1 (n_2077), .B2 (n_2079));
NAND2_X1 i_2139 (.ZN (n_2075), .A1 (n_2091), .A2 (n_2076));
INV_X1 i_2138 (.ZN (n_2074), .A (n_2076));
NAND3_X1 i_2137 (.ZN (n_2073), .A1 (n_2074), .A2 (n_2093), .A3 (n_2092));
NAND2_X1 i_2136 (.ZN (n_2072), .A1 (B_imm[6]), .A2 (A_imm[6]));
OAI22_X1 i_2135 (.ZN (n_2071), .A1 (n_8880), .A2 (n_6836), .B1 (n_8926), .B2 (n_6740));
NAND2_X1 i_2134 (.ZN (n_2070), .A1 (B_imm[7]), .A2 (A_imm[4]));
NAND4_X1 i_2133 (.ZN (n_2069), .A1 (B_imm[10]), .A2 (A_imm[11]), .A3 (B_imm[0]), .A4 (A_imm[1]));
NAND2_X1 i_2132 (.ZN (n_2068), .A1 (n_2069), .A2 (n_2070));
NAND2_X1 i_2131 (.ZN (n_2067), .A1 (n_2068), .A2 (n_2071));
NAND2_X1 i_2130 (.ZN (n_2066), .A1 (n_2067), .A2 (n_2072));
INV_X1 i_2129 (.ZN (n_2065), .A (n_2072));
NAND3_X1 i_2128 (.ZN (n_2064), .A1 (n_2065), .A2 (n_2071), .A3 (n_2068));
INV_X1 i_2127 (.ZN (n_2063), .A (n_2064));
NAND2_X1 i_2126 (.ZN (n_2062), .A1 (B_imm[8]), .A2 (A_imm[4]));
INV_X1 i_2125 (.ZN (n_2061), .A (n_2062));
OAI21_X1 i_2124 (.ZN (n_2060), .A (n_2066), .B1 (n_2063), .B2 (n_2061));
INV_X1 i_2123 (.ZN (n_2059), .A (n_2060));
AOI21_X1 i_2122 (.ZN (n_2058), .A (n_2197), .B1 (n_2198), .B2 (n_2195));
NAND3_X1 i_2121 (.ZN (n_2057), .A1 (n_2198), .A2 (n_2197), .A3 (n_2195));
INV_X1 i_2120 (.ZN (n_2056), .A (n_2057));
OAI21_X1 i_2119 (.ZN (n_2055), .A (n_2059), .B1 (n_2058), .B2 (n_2056));
INV_X1 i_2118 (.ZN (n_2054), .A (n_2058));
NAND3_X1 i_2117 (.ZN (n_2053), .A1 (n_2060), .A2 (n_2054), .A3 (n_2057));
NAND2_X1 i_2116 (.ZN (n_2052), .A1 (B_imm[12]), .A2 (A_imm[0]));
OAI21_X1 i_2115 (.ZN (n_2051), .A (n_2052), .B1 (n_8849), .B2 (n_6836));
NAND2_X1 i_2114 (.ZN (n_2050), .A1 (B_imm[9]), .A2 (A_imm[3]));
INV_X1 i_2113 (.ZN (n_2049), .A (n_2050));
NAND4_X1 i_2112 (.ZN (n_2048), .A1 (B_imm[11]), .A2 (B_imm[12]), .A3 (A_imm[1]), .A4 (A_imm[0]));
INV_X1 i_2111 (.ZN (n_2047), .A (n_2048));
OAI21_X1 i_2110 (.ZN (n_2046), .A (n_2051), .B1 (n_2047), .B2 (n_2049));
INV_X1 i_2109 (.ZN (n_2045), .A (n_2046));
NAND2_X1 i_2108 (.ZN (n_2044), .A1 (n_2053), .A2 (n_2045));
NAND2_X1 i_2107 (.ZN (n_2043), .A1 (n_2044), .A2 (n_2055));
NAND2_X2 i_2106 (.ZN (n_2042), .A1 (n_2043), .A2 (n_2073));
NAND2_X1 i_2105 (.ZN (n_2041), .A1 (n_2042), .A2 (n_2075));
NAND2_X1 i_2104 (.ZN (n_2040), .A1 (n_2041), .A2 (n_2095));
INV_X1 i_2103 (.ZN (n_2039), .A (n_2095));
NAND3_X1 i_2102 (.ZN (n_2038), .A1 (n_2042), .A2 (n_2039), .A3 (n_2075));
INV_X1 i_2101 (.ZN (n_2037), .A (n_2038));
AOI21_X1 i_2100 (.ZN (n_2036), .A (n_2179), .B1 (n_2181), .B2 (n_2182));
NAND3_X1 i_2099 (.ZN (n_2035), .A1 (n_2182), .A2 (n_2181), .A3 (n_2179));
INV_X1 i_2098 (.ZN (n_2034), .A (n_2035));
NOR2_X1 i_2097 (.ZN (n_2033), .A1 (n_2034), .A2 (n_2036));
INV_X1 i_2096 (.ZN (n_2032), .A (n_2033));
OAI21_X1 i_2095 (.ZN (n_2031), .A (n_2040), .B1 (n_2037), .B2 (n_2032));
INV_X1 i_2094 (.ZN (n_2030), .A (n_2261));
OAI21_X1 i_2093 (.ZN (n_2029), .A (n_2256), .B1 (n_2030), .B2 (n_2260));
NAND2_X1 i_2092 (.ZN (n_2028), .A1 (n_2262), .A2 (n_2269));
NAND3_X1 i_2091 (.ZN (n_2027), .A1 (n_2028), .A2 (n_2286), .A3 (n_2285));
INV_X1 i_2090 (.ZN (n_2026), .A (n_2256));
NAND3_X1 i_2089 (.ZN (n_2025), .A1 (n_2027), .A2 (n_2026), .A3 (n_2261));
NAND2_X1 i_2088 (.ZN (n_2024), .A1 (n_2029), .A2 (n_2025));
INV_X1 i_2087 (.ZN (n_2023), .A (n_2024));
NAND2_X1 i_2086 (.ZN (n_2022), .A1 (n_2031), .A2 (n_2023));
OAI211_X1 i_2085 (.ZN (n_2021), .A (n_2024), .B (n_2040), .C1 (n_2037), .C2 (n_2032));
NAND3_X1 i_2084 (.ZN (n_2020), .A1 (n_2022), .A2 (n_2099), .A3 (n_2021));
INV_X1 i_2083 (.ZN (n_2019), .A (n_2099));
NAND2_X1 i_2082 (.ZN (n_2018), .A1 (n_2022), .A2 (n_2021));
NAND2_X1 i_2081 (.ZN (n_2017), .A1 (n_2018), .A2 (n_2019));
NAND2_X1 i_2080 (.ZN (n_2016), .A1 (n_2017), .A2 (n_2020));
INV_X1 i_2079 (.ZN (n_2015), .A (n_2293));
NAND2_X1 i_2078 (.ZN (n_2014), .A1 (n_2302), .A2 (n_2300));
NAND2_X1 i_2077 (.ZN (n_2013), .A1 (n_2014), .A2 (n_2015));
NAND3_X1 i_2076 (.ZN (n_2012), .A1 (n_2302), .A2 (n_2300), .A3 (n_2293));
NAND3_X1 i_2075 (.ZN (n_2011), .A1 (n_2294), .A2 (n_2299), .A3 (n_2297));
INV_X1 i_2074 (.ZN (n_2010), .A (n_2294));
NAND2_X1 i_2073 (.ZN (n_2009), .A1 (n_2297), .A2 (n_2299));
NAND2_X1 i_2072 (.ZN (n_2008), .A1 (n_2009), .A2 (n_2010));
NAND2_X1 i_2071 (.ZN (n_2007), .A1 (n_2008), .A2 (n_2011));
INV_X1 i_2070 (.ZN (n_2006), .A (n_2007));
OAI22_X1 i_2069 (.ZN (n_2005), .A1 (n_8849), .A2 (n_6677), .B1 (n_8795), .B2 (n_6836));
NAND2_X1 i_2068 (.ZN (n_2004), .A1 (B_imm[9]), .A2 (A_imm[4]));
INV_X1 i_2067 (.ZN (n_2003), .A (n_2004));
NAND4_X1 i_2066 (.ZN (n_2002), .A1 (B_imm[11]), .A2 (B_imm[12]), .A3 (A_imm[2]), .A4 (A_imm[1]));
INV_X1 i_2065 (.ZN (n_2001), .A (n_2002));
OAI21_X1 i_2064 (.ZN (n_2000), .A (n_2005), .B1 (n_2003), .B2 (n_2001));
NAND2_X1 i_2063 (.ZN (n_1999), .A1 (n_2399), .A2 (n_2396));
NAND2_X1 i_2062 (.ZN (n_1998), .A1 (n_1999), .A2 (n_2397));
NAND3_X1 i_2061 (.ZN (n_1997), .A1 (n_2399), .A2 (n_2398), .A3 (n_2396));
NAND3_X1 i_2060 (.ZN (n_1996), .A1 (n_2000), .A2 (n_1998), .A3 (n_1997));
NAND2_X1 i_2059 (.ZN (n_1995), .A1 (n_1998), .A2 (n_1997));
OAI211_X1 i_2058 (.ZN (n_1994), .A (n_1995), .B (n_2005), .C1 (n_2003), .C2 (n_2001));
OAI22_X1 i_2057 (.ZN (n_1993), .A1 (n_8947), .A2 (n_8293), .B1 (n_8232), .B2 (n_8644));
OAI22_X1 i_2056 (.ZN (n_1992), .A1 (n_8573), .A2 (n_8293), .B1 (n_8880), .B2 (n_6677));
NAND2_X1 i_2055 (.ZN (n_1991), .A1 (A_imm[9]), .A2 (B_imm[3]));
INV_X1 i_2054 (.ZN (n_1990), .A (n_1991));
NAND4_X1 i_2053 (.ZN (n_1989), .A1 (B_imm[7]), .A2 (B_imm[10]), .A3 (A_imm[5]), .A4 (A_imm[2]));
INV_X1 i_2052 (.ZN (n_1988), .A (n_1989));
OAI21_X1 i_2051 (.ZN (n_1987), .A (n_1992), .B1 (n_1990), .B2 (n_1988));
INV_X1 i_2050 (.ZN (n_1986), .A (n_1987));
NAND4_X1 i_2049 (.ZN (n_1985), .A1 (B_imm[8]), .A2 (B_imm[6]), .A3 (A_imm[7]), .A4 (A_imm[5]));
INV_X1 i_2048 (.ZN (n_1984), .A (n_1985));
OAI21_X1 i_2047 (.ZN (n_1983), .A (n_1993), .B1 (n_1986), .B2 (n_1984));
NAND2_X1 i_2046 (.ZN (n_1982), .A1 (n_1994), .A2 (n_1983));
NAND2_X1 i_2045 (.ZN (n_1981), .A1 (n_1982), .A2 (n_1996));
NAND2_X1 i_2044 (.ZN (n_1980), .A1 (n_1981), .A2 (n_2006));
NAND3_X1 i_2043 (.ZN (n_1979), .A1 (n_2007), .A2 (n_1996), .A3 (n_1982));
INV_X1 i_2042 (.ZN (n_1978), .A (n_2273));
INV_X1 i_2041 (.ZN (n_1977), .A (n_2272));
OAI21_X1 i_2040 (.ZN (n_1976), .A (n_1978), .B1 (n_2279), .B2 (n_1977));
INV_X1 i_2039 (.ZN (n_1975), .A (n_2279));
NAND3_X1 i_2038 (.ZN (n_1974), .A1 (n_1975), .A2 (n_2273), .A3 (n_2272));
OAI211_X1 i_2037 (.ZN (n_1973), .A (n_1976), .B (n_1974), .C1 (n_7913), .C2 (n_3554));
NAND2_X1 i_2036 (.ZN (n_1972), .A1 (n_1976), .A2 (n_1974));
NAND3_X1 i_2035 (.ZN (n_1971), .A1 (n_1972), .A2 (B_imm[14]), .A3 (A_imm[0]));
NAND2_X1 i_2034 (.ZN (n_1970), .A1 (n_2199), .A2 (n_2191));
NAND2_X1 i_2033 (.ZN (n_1969), .A1 (n_1970), .A2 (n_2192));
NAND3_X1 i_2032 (.ZN (n_1968), .A1 (n_2199), .A2 (n_2193), .A3 (n_2191));
NAND2_X1 i_2031 (.ZN (n_1967), .A1 (n_1969), .A2 (n_1968));
INV_X1 i_2030 (.ZN (n_1966), .A (n_1967));
NAND2_X1 i_2029 (.ZN (n_1965), .A1 (n_1971), .A2 (n_1966));
NAND2_X1 i_2028 (.ZN (n_1964), .A1 (n_1965), .A2 (n_1973));
NAND2_X1 i_2027 (.ZN (n_1963), .A1 (n_1979), .A2 (n_1964));
NAND2_X1 i_2026 (.ZN (n_1962), .A1 (n_1963), .A2 (n_1980));
AOI21_X1 i_2025 (.ZN (n_1961), .A (n_2379), .B1 (n_2384), .B2 (n_2385));
NAND3_X1 i_2024 (.ZN (n_1960), .A1 (n_2385), .A2 (n_2384), .A3 (n_2379));
INV_X1 i_2023 (.ZN (n_1959), .A (n_1960));
OAI21_X1 i_2022 (.ZN (n_1958), .A (n_1962), .B1 (n_1961), .B2 (n_1959));
NOR2_X1 i_2021 (.ZN (n_1957), .A1 (n_1959), .A2 (n_1961));
NAND3_X1 i_2020 (.ZN (n_1956), .A1 (n_1963), .A2 (n_1957), .A3 (n_1980));
NAND4_X1 i_2019 (.ZN (n_1955), .A1 (n_1958), .A2 (n_2013), .A3 (n_2012), .A4 (n_1956));
NAND2_X1 i_2018 (.ZN (n_1954), .A1 (n_2013), .A2 (n_2012));
AOI21_X1 i_2017 (.ZN (n_1953), .A (n_1957), .B1 (n_1963), .B2 (n_1980));
INV_X1 i_2016 (.ZN (n_1952), .A (n_1956));
OAI21_X1 i_2015 (.ZN (n_1951), .A (n_1954), .B1 (n_1952), .B2 (n_1953));
NAND2_X1 i_2014 (.ZN (n_1950), .A1 (n_1955), .A2 (n_1951));
INV_X1 i_2013 (.ZN (n_1949), .A (n_1950));
NAND2_X1 i_2012 (.ZN (n_1948), .A1 (n_2150), .A2 (n_2151));
NAND2_X1 i_2011 (.ZN (n_1947), .A1 (n_1948), .A2 (n_2145));
OAI211_X1 i_2010 (.ZN (n_1946), .A (n_2151), .B (n_2150), .C1 (n_2148), .C2 (n_2146));
NAND2_X1 i_2009 (.ZN (n_1945), .A1 (n_1947), .A2 (n_1946));
INV_X1 i_2008 (.ZN (n_1944), .A (n_1945));
NAND2_X1 i_2007 (.ZN (n_1943), .A1 (n_2165), .A2 (n_2164));
INV_X1 i_2006 (.ZN (n_1942), .A (n_1943));
OAI21_X1 i_2005 (.ZN (n_1941), .A (n_2173), .B1 (n_1942), .B2 (n_2171));
NAND2_X1 i_2004 (.ZN (n_1940), .A1 (n_1941), .A2 (n_2162));
NAND3_X1 i_2003 (.ZN (n_1939), .A1 (n_1940), .A2 (n_2160), .A3 (n_2159));
NAND3_X1 i_2002 (.ZN (n_1938), .A1 (n_1941), .A2 (n_2162), .A3 (n_2158));
NAND2_X1 i_2001 (.ZN (n_1937), .A1 (n_1939), .A2 (n_1938));
INV_X1 i_2000 (.ZN (n_1936), .A (n_1937));
NAND2_X1 i_1999 (.ZN (n_1935), .A1 (n_1993), .A2 (n_1985));
NAND2_X1 i_1998 (.ZN (n_1934), .A1 (n_1935), .A2 (n_1986));
NAND3_X1 i_1997 (.ZN (n_1933), .A1 (n_1993), .A2 (n_1987), .A3 (n_1985));
NAND2_X1 i_1996 (.ZN (n_1932), .A1 (n_1934), .A2 (n_1933));
INV_X1 i_1995 (.ZN (n_1931), .A (n_2165));
INV_X1 i_1994 (.ZN (n_1930), .A (n_2164));
OAI21_X1 i_1993 (.ZN (n_1929), .A (n_1931), .B1 (n_1930), .B2 (n_2171));
INV_X1 i_1992 (.ZN (n_1928), .A (n_2171));
NAND3_X1 i_1991 (.ZN (n_1927), .A1 (n_1928), .A2 (n_2165), .A3 (n_2164));
NAND2_X1 i_1990 (.ZN (n_1926), .A1 (n_1929), .A2 (n_1927));
NAND2_X1 i_1989 (.ZN (n_1925), .A1 (n_1932), .A2 (n_1926));
NAND4_X1 i_1988 (.ZN (n_1924), .A1 (n_1934), .A2 (n_1933), .A3 (n_1929), .A4 (n_1927));
INV_X1 i_1987 (.ZN (n_1923), .A (n_2005));
OAI21_X1 i_1986 (.ZN (n_1922), .A (n_2003), .B1 (n_1923), .B2 (n_2001));
NAND3_X1 i_1985 (.ZN (n_1921), .A1 (n_2005), .A2 (n_2004), .A3 (n_2002));
NAND2_X1 i_1984 (.ZN (n_1920), .A1 (n_1922), .A2 (n_1921));
NAND2_X1 i_1983 (.ZN (n_1919), .A1 (n_1920), .A2 (n_1924));
NAND2_X1 i_1982 (.ZN (n_1918), .A1 (n_1919), .A2 (n_1925));
NAND2_X1 i_1981 (.ZN (n_1917), .A1 (n_1918), .A2 (n_1936));
NAND3_X1 i_1980 (.ZN (n_1916), .A1 (n_1937), .A2 (n_1925), .A3 (n_1919));
NAND3_X1 i_1979 (.ZN (n_1915), .A1 (n_1996), .A2 (n_1994), .A3 (n_1983));
INV_X1 i_1978 (.ZN (n_1914), .A (n_1983));
NAND2_X1 i_1977 (.ZN (n_1913), .A1 (n_1996), .A2 (n_1994));
NAND2_X1 i_1976 (.ZN (n_1912), .A1 (n_1913), .A2 (n_1914));
NAND2_X1 i_1975 (.ZN (n_1911), .A1 (n_1912), .A2 (n_1915));
NAND2_X1 i_1974 (.ZN (n_1910), .A1 (n_1916), .A2 (n_1911));
NAND2_X1 i_1973 (.ZN (n_1909), .A1 (n_1910), .A2 (n_1917));
NAND2_X1 i_1972 (.ZN (n_1908), .A1 (n_1909), .A2 (n_1944));
NAND3_X1 i_1971 (.ZN (n_1907), .A1 (n_1910), .A2 (n_1945), .A3 (n_1917));
NAND3_X1 i_1970 (.ZN (n_1906), .A1 (n_1980), .A2 (n_1979), .A3 (n_1964));
NAND2_X1 i_1969 (.ZN (n_1905), .A1 (n_1980), .A2 (n_1979));
NAND3_X1 i_1968 (.ZN (n_1904), .A1 (n_1905), .A2 (n_1973), .A3 (n_1965));
NAND2_X1 i_1967 (.ZN (n_1903), .A1 (n_1904), .A2 (n_1906));
NAND2_X1 i_1966 (.ZN (n_1902), .A1 (n_1903), .A2 (n_1907));
NAND2_X1 i_1965 (.ZN (n_1901), .A1 (n_1902), .A2 (n_1908));
NAND2_X1 i_1964 (.ZN (n_1900), .A1 (n_1949), .A2 (n_1901));
INV_X1 i_1963 (.ZN (n_1899), .A (n_1901));
NAND2_X1 i_1962 (.ZN (n_1898), .A1 (n_1899), .A2 (n_1950));
NAND3_X1 i_1961 (.ZN (n_1897), .A1 (n_2016), .A2 (n_1900), .A3 (n_1898));
INV_X1 i_1960 (.ZN (n_1896), .A (n_2020));
AOI21_X1 i_1959 (.ZN (n_1895), .A (n_2099), .B1 (n_2022), .B2 (n_2021));
NOR2_X2 i_1958 (.ZN (n_1894), .A1 (n_1896), .A2 (n_1895));
NAND2_X1 i_1957 (.ZN (n_1893), .A1 (n_1900), .A2 (n_1898));
NAND2_X1 i_1956 (.ZN (n_1892), .A1 (n_1893), .A2 (n_1894));
NAND3_X1 i_1955 (.ZN (n_1891), .A1 (n_1973), .A2 (n_1971), .A3 (n_1966));
NAND2_X1 i_1954 (.ZN (n_1890), .A1 (n_1973), .A2 (n_1971));
NAND2_X1 i_1953 (.ZN (n_1889), .A1 (n_1890), .A2 (n_1967));
NAND2_X1 i_1952 (.ZN (n_1888), .A1 (n_1889), .A2 (n_1891));
INV_X1 i_1951 (.ZN (n_1887), .A (n_2079));
XNOR2_X1 i_1950 (.ZN (n_1886), .A (n_2078), .B (n_2276));
AOI21_X1 i_1949 (.ZN (n_1885), .A (n_1886), .B1 (n_1887), .B2 (n_2080));
NAND3_X1 i_1948 (.ZN (n_1884), .A1 (n_1887), .A2 (n_2080), .A3 (n_1886));
INV_X1 i_1947 (.ZN (n_1883), .A (n_1884));
NOR2_X1 i_1946 (.ZN (n_1882), .A1 (n_1883), .A2 (n_1885));
OAI22_X1 i_1945 (.ZN (n_1881), .A1 (n_8751), .A2 (n_4366), .B1 (n_8645), .B2 (n_6584));
OAI22_X1 i_1944 (.ZN (n_1880), .A1 (n_8511), .A2 (n_6584), .B1 (n_6817), .B2 (n_8644));
NAND2_X1 i_1943 (.ZN (n_1879), .A1 (B_imm[4]), .A2 (A_imm[6]));
INV_X1 i_1942 (.ZN (n_1878), .A (n_1879));
NAND4_X1 i_1941 (.ZN (n_1877), .A1 (A_imm[8]), .A2 (B_imm[3]), .A3 (B_imm[2]), .A4 (A_imm[7]));
INV_X1 i_1940 (.ZN (n_1876), .A (n_1877));
OAI21_X1 i_1939 (.ZN (n_1875), .A (n_1880), .B1 (n_1878), .B2 (n_1876));
NAND4_X1 i_1938 (.ZN (n_1874), .A1 (A_imm[10]), .A2 (B_imm[2]), .A3 (B_imm[1]), .A4 (A_imm[9]));
NAND2_X1 i_1937 (.ZN (n_1873), .A1 (n_1874), .A2 (n_1875));
NAND2_X1 i_1936 (.ZN (n_1872), .A1 (n_1873), .A2 (n_1881));
INV_X1 i_1935 (.ZN (n_1871), .A (n_1872));
AOI21_X1 i_1934 (.ZN (n_1870), .A (n_2169), .B1 (n_2170), .B2 (n_2167));
NAND3_X1 i_1933 (.ZN (n_1869), .A1 (n_2170), .A2 (n_2169), .A3 (n_2167));
INV_X1 i_1932 (.ZN (n_1868), .A (n_1869));
OAI21_X1 i_1931 (.ZN (n_1867), .A (n_1871), .B1 (n_1870), .B2 (n_1868));
INV_X1 i_1930 (.ZN (n_1866), .A (n_1867));
NOR2_X1 i_1929 (.ZN (n_1865), .A1 (n_1870), .A2 (n_1868));
NAND2_X1 i_1928 (.ZN (n_1864), .A1 (n_1865), .A2 (n_1872));
NAND2_X1 i_1927 (.ZN (n_1863), .A1 (n_1992), .A2 (n_1989));
XNOR2_X1 i_1926 (.ZN (n_1862), .A (n_1863), .B (n_1991));
INV_X1 i_1925 (.ZN (n_1861), .A (n_1862));
AOI21_X1 i_1924 (.ZN (n_1860), .A (n_1866), .B1 (n_1861), .B2 (n_1864));
INV_X1 i_1923 (.ZN (n_1859), .A (n_1860));
NAND2_X1 i_1922 (.ZN (n_1858), .A1 (n_1882), .A2 (n_1859));
OAI21_X1 i_1921 (.ZN (n_1857), .A (n_1860), .B1 (n_1885), .B2 (n_1883));
NAND2_X1 i_1919 (.ZN (n_1855), .A1 (A_imm[8]), .A2 (B_imm[1]));
NAND4_X1 i_1918 (.ZN (n_1854), .A1 (B_imm[2]), .A2 (A_imm[6]), .A3 (B_imm[3]), .A4 (A_imm[7]));
NAND2_X1 i_1917 (.ZN (n_1853), .A1 (n_1854), .A2 (n_1855));
NAND2_X1 i_1916 (.ZN (n_1852), .A1 (n_1853), .A2 (n_1856));
OAI21_X1 i_1915 (.ZN (n_1851), .A (n_1852), .B1 (n_8645), .B2 (n_4366));
NAND2_X1 i_1914 (.ZN (n_1850), .A1 (A_imm[10]), .A2 (B_imm[0]));
NAND4_X1 i_1913 (.ZN (n_1849), .A1 (A_imm[9]), .A2 (n_1853), .A3 (n_1856), .A4 (B_imm[1]));
NAND2_X1 i_1912 (.ZN (n_1848), .A1 (n_1849), .A2 (n_1850));
NAND2_X1 i_1911 (.ZN (n_1847), .A1 (n_1848), .A2 (n_1851));
OAI21_X1 i_1910 (.ZN (n_1846), .A (n_1847), .B1 (n_8849), .B2 (n_3554));
NAND2_X1 i_1909 (.ZN (n_1845), .A1 (B_imm[9]), .A2 (A_imm[2]));
NAND4_X1 i_1908 (.ZN (n_1844), .A1 (n_1848), .A2 (B_imm[11]), .A3 (n_1851), .A4 (A_imm[0]));
NAND2_X1 i_1907 (.ZN (n_1843), .A1 (n_1844), .A2 (n_1845));
OAI22_X1 i_1906 (.ZN (n_1842), .A1 (n_8880), .A2 (n_3554), .B1 (n_8429), .B2 (n_8293));
NAND2_X1 i_1905 (.ZN (n_1841), .A1 (B_imm[7]), .A2 (A_imm[3]));
NAND4_X1 i_1904 (.ZN (n_1840), .A1 (B_imm[10]), .A2 (B_imm[5]), .A3 (A_imm[5]), .A4 (A_imm[0]));
NAND2_X1 i_1903 (.ZN (n_1839), .A1 (n_1840), .A2 (n_1841));
NAND2_X1 i_1902 (.ZN (n_1838), .A1 (n_1839), .A2 (n_1842));
OAI21_X1 i_1901 (.ZN (n_1837), .A (n_1838), .B1 (n_8232), .B2 (n_8293));
NAND4_X1 i_1900 (.ZN (n_1836), .A1 (n_1839), .A2 (n_1842), .A3 (B_imm[6]), .A4 (A_imm[5]));
NAND2_X1 i_1899 (.ZN (n_1835), .A1 (B_imm[8]), .A2 (A_imm[3]));
NAND2_X1 i_1898 (.ZN (n_1834), .A1 (n_1836), .A2 (n_1835));
NAND4_X1 i_1897 (.ZN (n_1833), .A1 (n_1843), .A2 (n_1834), .A3 (n_1846), .A4 (n_1837));
NAND2_X1 i_1896 (.ZN (n_1832), .A1 (n_1843), .A2 (n_1846));
AOI22_X1 i_1895 (.ZN (n_1831), .A1 (n_1839), .A2 (n_1842), .B1 (B_imm[6]), .B2 (A_imm[5]));
INV_X1 i_1894 (.ZN (n_1830), .A (n_1834));
OAI21_X1 i_1893 (.ZN (n_1829), .A (n_1832), .B1 (n_1831), .B2 (n_1830));
NAND2_X1 i_1892 (.ZN (n_1828), .A1 (n_2084), .A2 (n_2083));
NAND3_X1 i_1891 (.ZN (n_1827), .A1 (n_1828), .A2 (B_imm[0]), .A3 (A_imm[12]));
NAND3_X1 i_1890 (.ZN (n_1826), .A1 (n_2084), .A2 (n_2083), .A3 (n_2082));
NAND2_X1 i_1889 (.ZN (n_1825), .A1 (n_1827), .A2 (n_1826));
NAND2_X1 i_1888 (.ZN (n_1824), .A1 (n_1829), .A2 (n_1825));
NAND2_X1 i_1887 (.ZN (n_1823), .A1 (n_1824), .A2 (n_1833));
NAND2_X1 i_1886 (.ZN (n_1822), .A1 (n_1857), .A2 (n_1823));
NAND2_X1 i_1885 (.ZN (n_1821), .A1 (n_1822), .A2 (n_1858));
NAND2_X1 i_1884 (.ZN (n_1820), .A1 (n_1821), .A2 (n_1888));
NAND4_X1 i_1883 (.ZN (n_1819), .A1 (n_1822), .A2 (n_1891), .A3 (n_1889), .A4 (n_1858));
NAND3_X1 i_1882 (.ZN (n_1818), .A1 (n_2073), .A2 (n_2043), .A3 (n_2075));
INV_X1 i_1881 (.ZN (n_1817), .A (n_2043));
NAND2_X1 i_1880 (.ZN (n_1816), .A1 (n_2073), .A2 (n_2075));
NAND2_X1 i_1879 (.ZN (n_1815), .A1 (n_1816), .A2 (n_1817));
NAND2_X1 i_1878 (.ZN (n_1814), .A1 (n_1815), .A2 (n_1818));
INV_X1 i_1877 (.ZN (n_1813), .A (n_1814));
NAND2_X1 i_1876 (.ZN (n_1812), .A1 (n_1819), .A2 (n_1813));
NAND2_X1 i_1875 (.ZN (n_1811), .A1 (n_1812), .A2 (n_1820));
NAND3_X1 i_1874 (.ZN (n_1810), .A1 (n_2040), .A2 (n_2038), .A3 (n_2033));
AOI22_X1 i_1873 (.ZN (n_1809), .A1 (n_2042), .A2 (n_2075), .B1 (n_2098), .B2 (n_2096));
OAI21_X1 i_1872 (.ZN (n_1808), .A (n_2032), .B1 (n_2037), .B2 (n_1809));
NAND3_X1 i_1871 (.ZN (n_1807), .A1 (n_1811), .A2 (n_1810), .A3 (n_1808));
INV_X1 i_1870 (.ZN (n_1806), .A (n_1811));
NAND2_X1 i_1869 (.ZN (n_1805), .A1 (n_1808), .A2 (n_1810));
NAND2_X1 i_1868 (.ZN (n_1804), .A1 (n_1806), .A2 (n_1805));
INV_X1 i_1867 (.ZN (n_1803), .A (n_1804));
NAND3_X1 i_1866 (.ZN (n_1802), .A1 (n_1908), .A2 (n_1907), .A3 (n_1903));
INV_X1 i_1865 (.ZN (n_1801), .A (n_1903));
NAND2_X1 i_1864 (.ZN (n_1800), .A1 (n_1908), .A2 (n_1907));
NAND2_X1 i_1863 (.ZN (n_1799), .A1 (n_1800), .A2 (n_1801));
NAND2_X1 i_1862 (.ZN (n_1798), .A1 (n_1799), .A2 (n_1802));
OAI21_X1 i_1861 (.ZN (n_1797), .A (n_1807), .B1 (n_1798), .B2 (n_1803));
NAND3_X2 i_1860 (.ZN (n_1796), .A1 (n_1897), .A2 (n_1892), .A3 (n_1797));
INV_X2 i_1859 (.ZN (n_1795), .A (n_1796));
AOI21_X1 i_1858 (.ZN (n_1794), .A (n_1797), .B1 (n_1892), .B2 (n_1897));
NAND3_X1 i_1857 (.ZN (n_1793), .A1 (n_1798), .A2 (n_1807), .A3 (n_1804));
INV_X1 i_1856 (.ZN (n_1792), .A (n_1802));
AOI21_X1 i_1855 (.ZN (n_1791), .A (n_1903), .B1 (n_1908), .B2 (n_1907));
NOR2_X1 i_1854 (.ZN (n_1790), .A1 (n_1792), .A2 (n_1791));
NAND2_X1 i_1853 (.ZN (n_1789), .A1 (n_1804), .A2 (n_1807));
NAND2_X1 i_1852 (.ZN (n_1788), .A1 (n_1789), .A2 (n_1790));
NAND3_X1 i_1851 (.ZN (n_1787), .A1 (n_1917), .A2 (n_1916), .A3 (n_1911));
INV_X1 i_1850 (.ZN (n_1786), .A (n_1911));
NAND2_X1 i_1849 (.ZN (n_1785), .A1 (n_1917), .A2 (n_1916));
NAND2_X1 i_1848 (.ZN (n_1784), .A1 (n_1785), .A2 (n_1786));
NAND2_X1 i_1847 (.ZN (n_1783), .A1 (n_2051), .A2 (n_2048));
NAND2_X1 i_1846 (.ZN (n_1782), .A1 (n_1783), .A2 (n_2049));
NAND3_X1 i_1845 (.ZN (n_1781), .A1 (n_2051), .A2 (n_2050), .A3 (n_2048));
NAND2_X1 i_1844 (.ZN (n_1780), .A1 (n_1782), .A2 (n_1781));
NAND2_X1 i_1843 (.ZN (n_1779), .A1 (n_2066), .A2 (n_2064));
NAND2_X1 i_1842 (.ZN (n_1778), .A1 (n_1779), .A2 (n_2061));
NAND3_X1 i_1841 (.ZN (n_1777), .A1 (n_2066), .A2 (n_2064), .A3 (n_2062));
NAND2_X1 i_1840 (.ZN (n_1776), .A1 (n_1778), .A2 (n_1777));
NAND2_X1 i_1839 (.ZN (n_1775), .A1 (n_1780), .A2 (n_1776));
NAND4_X1 i_1838 (.ZN (n_1774), .A1 (n_1782), .A2 (n_1778), .A3 (n_1781), .A4 (n_1777));
AOI21_X1 i_1837 (.ZN (n_1773), .A (n_2070), .B1 (n_2071), .B2 (n_2069));
NAND3_X1 i_1836 (.ZN (n_1772), .A1 (n_2071), .A2 (n_2070), .A3 (n_2069));
INV_X1 i_1835 (.ZN (n_1771), .A (n_1772));
NAND2_X1 i_1834 (.ZN (n_1770), .A1 (n_2089), .A2 (n_2087));
NAND3_X1 i_1833 (.ZN (n_1769), .A1 (n_1770), .A2 (B_imm[5]), .A3 (A_imm[6]));
NAND3_X1 i_1832 (.ZN (n_1768), .A1 (n_2089), .A2 (n_2088), .A3 (n_2087));
NAND2_X1 i_1831 (.ZN (n_1767), .A1 (n_1769), .A2 (n_1768));
OAI21_X1 i_1830 (.ZN (n_1766), .A (n_1767), .B1 (n_1773), .B2 (n_1771));
NOR2_X1 i_1829 (.ZN (n_1765), .A1 (n_1773), .A2 (n_1771));
INV_X1 i_1828 (.ZN (n_1764), .A (n_1767));
NAND2_X1 i_1827 (.ZN (n_1763), .A1 (n_1765), .A2 (n_1764));
OAI22_X1 i_1826 (.ZN (n_1762), .A1 (n_8947), .A2 (n_6677), .B1 (n_8232), .B2 (n_6678));
OAI22_X1 i_1825 (.ZN (n_1761), .A1 (n_6584), .A2 (n_7691), .B1 (n_8644), .B2 (n_4366));
NAND2_X1 i_1824 (.ZN (n_1760), .A1 (A_imm[5]), .A2 (B_imm[3]));
NAND4_X1 i_1823 (.ZN (n_1759), .A1 (B_imm[2]), .A2 (A_imm[6]), .A3 (B_imm[1]), .A4 (A_imm[7]));
NAND2_X1 i_1822 (.ZN (n_1758), .A1 (n_1759), .A2 (n_1760));
AOI22_X1 i_1821 (.ZN (n_1757), .A1 (n_1758), .A2 (n_1761), .B1 (B_imm[4]), .B2 (A_imm[5]));
INV_X1 i_1820 (.ZN (n_1756), .A (n_1757));
NAND4_X1 i_1819 (.ZN (n_1755), .A1 (n_1758), .A2 (n_1761), .A3 (B_imm[4]), .A4 (A_imm[5]));
INV_X1 i_1818 (.ZN (n_1754), .A (n_1755));
NAND2_X1 i_1817 (.ZN (n_1753), .A1 (B_imm[5]), .A2 (A_imm[4]));
INV_X1 i_1816 (.ZN (n_1752), .A (n_1753));
OAI21_X1 i_1815 (.ZN (n_1751), .A (n_1756), .B1 (n_1754), .B2 (n_1752));
NAND4_X1 i_1814 (.ZN (n_1750), .A1 (B_imm[8]), .A2 (B_imm[6]), .A3 (A_imm[4]), .A4 (A_imm[2]));
NAND2_X1 i_1813 (.ZN (n_1749), .A1 (n_1751), .A2 (n_1750));
NAND2_X1 i_1812 (.ZN (n_1748), .A1 (n_1749), .A2 (n_1762));
INV_X1 i_1811 (.ZN (n_1747), .A (n_1748));
NAND2_X1 i_1810 (.ZN (n_1746), .A1 (n_1763), .A2 (n_1747));
NAND2_X1 i_1809 (.ZN (n_1745), .A1 (n_1746), .A2 (n_1766));
NAND2_X1 i_1808 (.ZN (n_1744), .A1 (n_1774), .A2 (n_1745));
NAND2_X1 i_1807 (.ZN (n_1743), .A1 (n_1744), .A2 (n_1775));
NAND2_X1 i_1806 (.ZN (n_1742), .A1 (n_2055), .A2 (n_2053));
NAND2_X1 i_1805 (.ZN (n_1741), .A1 (n_1742), .A2 (n_2046));
NAND3_X1 i_1804 (.ZN (n_1740), .A1 (n_2055), .A2 (n_2053), .A3 (n_2045));
NAND3_X1 i_1803 (.ZN (n_1739), .A1 (n_1743), .A2 (n_1741), .A3 (n_1740));
NAND2_X1 i_1802 (.ZN (n_1738), .A1 (n_1741), .A2 (n_1740));
NAND3_X1 i_1801 (.ZN (n_1737), .A1 (n_1738), .A2 (n_1775), .A3 (n_1744));
NAND2_X1 i_1800 (.ZN (n_1736), .A1 (n_1925), .A2 (n_1924));
NAND3_X1 i_1799 (.ZN (n_1735), .A1 (n_1736), .A2 (n_1922), .A3 (n_1921));
NAND3_X1 i_1798 (.ZN (n_1734), .A1 (n_1920), .A2 (n_1925), .A3 (n_1924));
NAND2_X1 i_1797 (.ZN (n_1733), .A1 (n_1735), .A2 (n_1734));
INV_X1 i_1796 (.ZN (n_1732), .A (n_1733));
NAND2_X1 i_1795 (.ZN (n_1731), .A1 (n_1737), .A2 (n_1732));
NAND2_X1 i_1794 (.ZN (n_1730), .A1 (n_1731), .A2 (n_1739));
NAND3_X1 i_1793 (.ZN (n_1729), .A1 (n_1730), .A2 (n_1787), .A3 (n_1784));
INV_X1 i_1792 (.ZN (n_1728), .A (n_1729));
NAND2_X1 i_1791 (.ZN (n_1727), .A1 (n_1784), .A2 (n_1787));
NAND3_X1 i_1790 (.ZN (n_1726), .A1 (n_1727), .A2 (n_1739), .A3 (n_1731));
NAND3_X1 i_1789 (.ZN (n_1725), .A1 (n_1820), .A2 (n_1819), .A3 (n_1814));
NAND2_X1 i_1788 (.ZN (n_1724), .A1 (n_1820), .A2 (n_1819));
NAND2_X1 i_1787 (.ZN (n_1723), .A1 (n_1724), .A2 (n_1813));
NAND2_X1 i_1786 (.ZN (n_1722), .A1 (n_1723), .A2 (n_1725));
AOI21_X1 i_1785 (.ZN (n_1721), .A (n_1728), .B1 (n_1722), .B2 (n_1726));
AOI21_X1 i_1784 (.ZN (n_1720), .A (n_1721), .B1 (n_1788), .B2 (n_1793));
INV_X1 i_1783 (.ZN (n_1719), .A (n_1720));
OAI21_X1 i_1782 (.ZN (n_1718), .A (n_1719), .B1 (n_1795), .B2 (n_1794));
INV_X1 i_1781 (.ZN (n_1717), .A (n_1718));
AOI21_X1 i_1780 (.ZN (n_1716), .A (n_1875), .B1 (n_1881), .B2 (n_1874));
NAND3_X1 i_1779 (.ZN (n_1715), .A1 (n_1881), .A2 (n_1875), .A3 (n_1874));
INV_X1 i_1778 (.ZN (n_1714), .A (n_1715));
NOR2_X1 i_1777 (.ZN (n_1713), .A1 (n_1716), .A2 (n_1714));
INV_X1 i_1776 (.ZN (n_1712), .A (n_1836));
INV_X1 i_1775 (.ZN (n_1711), .A (n_1835));
OAI21_X1 i_1774 (.ZN (n_1710), .A (n_1711), .B1 (n_1712), .B2 (n_1831));
NAND3_X1 i_1773 (.ZN (n_1709), .A1 (n_1837), .A2 (n_1836), .A3 (n_1835));
NAND3_X1 i_1772 (.ZN (n_1708), .A1 (n_1713), .A2 (n_1709), .A3 (n_1710));
AOI21_X1 i_1771 (.ZN (n_1707), .A (n_1713), .B1 (n_1710), .B2 (n_1709));
NAND2_X1 i_1770 (.ZN (n_1706), .A1 (B_imm[9]), .A2 (A_imm[1]));
NAND2_X1 i_1769 (.ZN (n_1705), .A1 (n_1880), .A2 (n_1877));
XNOR2_X1 i_1768 (.ZN (n_1704), .A (n_1705), .B (n_1878));
INV_X1 i_1767 (.ZN (n_1703), .A (n_1704));
NAND2_X1 i_1766 (.ZN (n_1702), .A1 (n_1703), .A2 (n_1706));
NAND3_X1 i_1765 (.ZN (n_1701), .A1 (n_1704), .A2 (B_imm[9]), .A3 (A_imm[1]));
INV_X1 i_1764 (.ZN (n_1700), .A (n_1701));
NAND2_X1 i_1763 (.ZN (n_1699), .A1 (n_1842), .A2 (n_1840));
NAND3_X1 i_1762 (.ZN (n_1698), .A1 (n_1699), .A2 (B_imm[7]), .A3 (A_imm[3]));
NAND3_X1 i_1761 (.ZN (n_1697), .A1 (n_1842), .A2 (n_1841), .A3 (n_1840));
NAND2_X1 i_1760 (.ZN (n_1696), .A1 (n_1698), .A2 (n_1697));
OAI21_X1 i_1759 (.ZN (n_1695), .A (n_1702), .B1 (n_1700), .B2 (n_1696));
INV_X1 i_1758 (.ZN (n_1694), .A (n_1695));
OAI21_X1 i_1757 (.ZN (n_1693), .A (n_1708), .B1 (n_1694), .B2 (n_1707));
INV_X1 i_1756 (.ZN (n_1692), .A (n_1864));
OAI21_X1 i_1755 (.ZN (n_1691), .A (n_1862), .B1 (n_1866), .B2 (n_1692));
NAND3_X1 i_1754 (.ZN (n_1690), .A1 (n_1861), .A2 (n_1867), .A3 (n_1864));
NAND2_X1 i_1753 (.ZN (n_1689), .A1 (n_1691), .A2 (n_1690));
NAND2_X1 i_1752 (.ZN (n_1688), .A1 (n_1693), .A2 (n_1689));
INV_X1 i_1751 (.ZN (n_1687), .A (n_1710));
INV_X1 i_1750 (.ZN (n_1686), .A (n_1709));
OAI22_X1 i_1749 (.ZN (n_1685), .A1 (n_1687), .A2 (n_1686), .B1 (n_1716), .B2 (n_1714));
NAND2_X1 i_1748 (.ZN (n_1684), .A1 (n_1685), .A2 (n_1695));
NAND4_X1 i_1747 (.ZN (n_1683), .A1 (n_1684), .A2 (n_1708), .A3 (n_1691), .A4 (n_1690));
NAND2_X1 i_1746 (.ZN (n_1682), .A1 (n_1829), .A2 (n_1833));
NAND3_X1 i_1745 (.ZN (n_1681), .A1 (n_1682), .A2 (n_1827), .A3 (n_1826));
NAND3_X1 i_1744 (.ZN (n_1680), .A1 (n_1829), .A2 (n_1833), .A3 (n_1825));
NAND2_X1 i_1743 (.ZN (n_1679), .A1 (n_1681), .A2 (n_1680));
NAND2_X1 i_1742 (.ZN (n_1678), .A1 (n_1679), .A2 (n_1683));
NAND2_X1 i_1741 (.ZN (n_1677), .A1 (n_1678), .A2 (n_1688));
NAND3_X1 i_1740 (.ZN (n_1676), .A1 (n_1858), .A2 (n_1857), .A3 (n_1823));
INV_X1 i_1739 (.ZN (n_1675), .A (n_1823));
NAND2_X1 i_1738 (.ZN (n_1674), .A1 (n_1858), .A2 (n_1857));
NAND2_X1 i_1737 (.ZN (n_1673), .A1 (n_1674), .A2 (n_1675));
NAND2_X1 i_1736 (.ZN (n_1672), .A1 (n_1673), .A2 (n_1676));
NAND2_X1 i_1735 (.ZN (n_1671), .A1 (n_1672), .A2 (n_1677));
NAND4_X1 i_1734 (.ZN (n_1670), .A1 (n_1673), .A2 (n_1678), .A3 (n_1688), .A4 (n_1676));
NAND3_X1 i_1733 (.ZN (n_1669), .A1 (n_1737), .A2 (n_1732), .A3 (n_1739));
NAND2_X1 i_1732 (.ZN (n_1668), .A1 (n_1737), .A2 (n_1739));
NAND2_X1 i_1731 (.ZN (n_1667), .A1 (n_1668), .A2 (n_1733));
NAND2_X1 i_1730 (.ZN (n_1666), .A1 (n_1667), .A2 (n_1669));
NAND3_X1 i_1729 (.ZN (n_1665), .A1 (n_1666), .A2 (n_1671), .A3 (n_1670));
NAND2_X1 i_1728 (.ZN (n_1664), .A1 (n_1671), .A2 (n_1670));
INV_X1 i_1727 (.ZN (n_1663), .A (n_1666));
NAND2_X1 i_1726 (.ZN (n_1662), .A1 (n_1664), .A2 (n_1663));
INV_X1 i_1725 (.ZN (n_1661), .A (n_1745));
NAND3_X1 i_1724 (.ZN (n_1660), .A1 (n_1775), .A2 (n_1661), .A3 (n_1774));
NAND2_X1 i_1723 (.ZN (n_1659), .A1 (n_1775), .A2 (n_1774));
NAND2_X1 i_1722 (.ZN (n_1658), .A1 (n_1659), .A2 (n_1745));
NAND2_X1 i_1721 (.ZN (n_1657), .A1 (n_1658), .A2 (n_1660));
OAI22_X1 i_1720 (.ZN (n_1656), .A1 (n_8947), .A2 (n_6836), .B1 (n_8232), .B2 (n_3718));
OAI22_X1 i_1719 (.ZN (n_1655), .A1 (n_4366), .A2 (n_7691), .B1 (n_8644), .B2 (n_6740));
NAND2_X1 i_1718 (.ZN (n_1654), .A1 (A_imm[4]), .A2 (B_imm[3]));
NAND4_X1 i_1717 (.ZN (n_1653), .A1 (A_imm[6]), .A2 (A_imm[7]), .A3 (B_imm[1]), .A4 (B_imm[0]));
NAND2_X1 i_1716 (.ZN (n_1652), .A1 (n_1653), .A2 (n_1654));
NAND2_X1 i_1715 (.ZN (n_1651), .A1 (n_1652), .A2 (n_1655));
OAI21_X1 i_1714 (.ZN (n_1650), .A (n_1651), .B1 (n_6740), .B2 (n_8511));
NAND4_X1 i_1713 (.ZN (n_1649), .A1 (n_1652), .A2 (n_1655), .A3 (B_imm[0]), .A4 (A_imm[8]));
INV_X1 i_1712 (.ZN (n_1648), .A (n_1649));
NAND2_X1 i_1711 (.ZN (n_1647), .A1 (B_imm[4]), .A2 (A_imm[4]));
INV_X1 i_1710 (.ZN (n_1646), .A (n_1647));
OAI21_X1 i_1709 (.ZN (n_1645), .A (n_1650), .B1 (n_1648), .B2 (n_1646));
NAND4_X1 i_1708 (.ZN (n_1644), .A1 (B_imm[8]), .A2 (B_imm[6]), .A3 (A_imm[3]), .A4 (A_imm[1]));
NAND2_X1 i_1707 (.ZN (n_1643), .A1 (n_1644), .A2 (n_1645));
NAND4_X1 i_1706 (.ZN (n_1642), .A1 (A_imm[9]), .A2 (B_imm[7]), .A3 (B_imm[0]), .A4 (A_imm[2]));
OAI22_X1 i_1705 (.ZN (n_1641), .A1 (n_8645), .A2 (n_6740), .B1 (n_8573), .B2 (n_6677));
NAND2_X1 i_1704 (.ZN (n_1640), .A1 (n_1856), .A2 (n_1854));
NAND3_X1 i_1703 (.ZN (n_1639), .A1 (n_1640), .A2 (B_imm[1]), .A3 (A_imm[8]));
NAND3_X1 i_1702 (.ZN (n_1638), .A1 (n_1856), .A2 (n_1855), .A3 (n_1854));
NAND2_X1 i_1701 (.ZN (n_1637), .A1 (n_1639), .A2 (n_1638));
NAND2_X1 i_1700 (.ZN (n_1636), .A1 (n_1637), .A2 (n_1641));
NAND2_X1 i_1699 (.ZN (n_1635), .A1 (n_1636), .A2 (n_1642));
NAND3_X1 i_1698 (.ZN (n_1634), .A1 (n_1635), .A2 (n_1656), .A3 (n_1643));
NAND2_X1 i_1697 (.ZN (n_1633), .A1 (n_1643), .A2 (n_1656));
NAND3_X1 i_1696 (.ZN (n_1632), .A1 (n_1633), .A2 (n_1642), .A3 (n_1636));
NAND2_X1 i_1695 (.ZN (n_1631), .A1 (n_1851), .A2 (n_1849));
NAND3_X1 i_1694 (.ZN (n_1630), .A1 (n_1631), .A2 (B_imm[0]), .A3 (A_imm[10]));
NAND3_X1 i_1693 (.ZN (n_1629), .A1 (n_1851), .A2 (n_1850), .A3 (n_1849));
NAND2_X1 i_1692 (.ZN (n_1628), .A1 (n_1630), .A2 (n_1629));
NAND2_X1 i_1691 (.ZN (n_1627), .A1 (n_1632), .A2 (n_1628));
NAND2_X1 i_1690 (.ZN (n_1626), .A1 (n_1627), .A2 (n_1634));
NAND2_X1 i_1689 (.ZN (n_1625), .A1 (n_1846), .A2 (n_1844));
NAND3_X1 i_1688 (.ZN (n_1624), .A1 (n_1625), .A2 (B_imm[9]), .A3 (A_imm[2]));
NAND3_X1 i_1687 (.ZN (n_1623), .A1 (n_1846), .A2 (n_1844), .A3 (n_1845));
NAND2_X1 i_1686 (.ZN (n_1622), .A1 (n_1624), .A2 (n_1623));
NAND2_X1 i_1685 (.ZN (n_1621), .A1 (n_1626), .A2 (n_1622));
NAND4_X1 i_1684 (.ZN (n_1620), .A1 (n_1627), .A2 (n_1624), .A3 (n_1634), .A4 (n_1623));
NAND3_X1 i_1683 (.ZN (n_1619), .A1 (n_1763), .A2 (n_1766), .A3 (n_1748));
NAND2_X1 i_1682 (.ZN (n_1618), .A1 (n_1763), .A2 (n_1766));
NAND2_X1 i_1681 (.ZN (n_1617), .A1 (n_1618), .A2 (n_1747));
NAND2_X1 i_1680 (.ZN (n_1616), .A1 (n_1617), .A2 (n_1619));
NAND2_X1 i_1679 (.ZN (n_1615), .A1 (n_1620), .A2 (n_1616));
NAND2_X1 i_1678 (.ZN (n_1614), .A1 (n_1615), .A2 (n_1621));
NAND2_X1 i_1677 (.ZN (n_1613), .A1 (n_1657), .A2 (n_1614));
NAND4_X1 i_1676 (.ZN (n_1612), .A1 (n_1658), .A2 (n_1615), .A3 (n_1660), .A4 (n_1621));
INV_X1 i_1675 (.ZN (n_1611), .A (n_1679));
NAND2_X1 i_1674 (.ZN (n_1610), .A1 (n_1683), .A2 (n_1688));
NAND2_X1 i_1673 (.ZN (n_1609), .A1 (n_1610), .A2 (n_1611));
NAND3_X1 i_1672 (.ZN (n_1608), .A1 (n_1679), .A2 (n_1683), .A3 (n_1688));
NAND2_X1 i_1671 (.ZN (n_1607), .A1 (n_1609), .A2 (n_1608));
NAND2_X1 i_1670 (.ZN (n_1606), .A1 (n_1607), .A2 (n_1612));
AND2_X1 i_1669 (.ZN (n_1605), .A1 (n_1606), .A2 (n_1613));
AOI21_X1 i_1668 (.ZN (n_1604), .A (n_1605), .B1 (n_1662), .B2 (n_1665));
NAND3_X1 i_1667 (.ZN (n_1603), .A1 (n_1722), .A2 (n_1729), .A3 (n_1726));
NAND2_X1 i_1666 (.ZN (n_1602), .A1 (n_1726), .A2 (n_1729));
NAND3_X1 i_1665 (.ZN (n_1601), .A1 (n_1602), .A2 (n_1725), .A3 (n_1723));
NAND2_X1 i_1664 (.ZN (n_1600), .A1 (n_1663), .A2 (n_1671));
NAND2_X1 i_1663 (.ZN (n_1599), .A1 (n_1600), .A2 (n_1670));
NAND3_X1 i_1662 (.ZN (n_1598), .A1 (n_1601), .A2 (n_1603), .A3 (n_1599));
NAND2_X1 i_1661 (.ZN (n_1597), .A1 (n_1601), .A2 (n_1603));
INV_X1 i_1660 (.ZN (n_1596), .A (n_1599));
NAND2_X1 i_1659 (.ZN (n_1595), .A1 (n_1597), .A2 (n_1596));
NAND3_X1 i_1658 (.ZN (n_1594), .A1 (n_1595), .A2 (n_1604), .A3 (n_1598));
INV_X1 i_1657 (.ZN (n_1593), .A (n_1604));
NAND3_X1 i_1656 (.ZN (n_1592), .A1 (n_1605), .A2 (n_1662), .A3 (n_1665));
NAND2_X1 i_1655 (.ZN (n_1591), .A1 (n_1613), .A2 (n_1612));
NAND3_X1 i_1654 (.ZN (n_1590), .A1 (n_1591), .A2 (n_1609), .A3 (n_1608));
INV_X1 i_1653 (.ZN (n_1589), .A (n_1591));
NAND2_X1 i_1652 (.ZN (n_1588), .A1 (n_1589), .A2 (n_1607));
NAND3_X1 i_1651 (.ZN (n_1587), .A1 (n_1685), .A2 (n_1708), .A3 (n_1695));
INV_X1 i_1650 (.ZN (n_1586), .A (n_1587));
AOI21_X1 i_1649 (.ZN (n_1585), .A (n_1695), .B1 (n_1685), .B2 (n_1708));
INV_X1 i_1648 (.ZN (n_1584), .A (n_1751));
NAND2_X1 i_1647 (.ZN (n_1583), .A1 (n_1762), .A2 (n_1750));
NAND2_X1 i_1646 (.ZN (n_1582), .A1 (n_1583), .A2 (n_1584));
NAND3_X1 i_1645 (.ZN (n_1581), .A1 (n_1762), .A2 (n_1751), .A3 (n_1750));
NAND2_X1 i_1644 (.ZN (n_1580), .A1 (n_1582), .A2 (n_1581));
OAI21_X1 i_1643 (.ZN (n_1579), .A (n_1752), .B1 (n_1754), .B2 (n_1757));
NAND3_X1 i_1642 (.ZN (n_1578), .A1 (n_1756), .A2 (n_1755), .A3 (n_1753));
NAND2_X1 i_1641 (.ZN (n_1577), .A1 (n_1578), .A2 (n_1579));
NAND3_X1 i_1640 (.ZN (n_1576), .A1 (n_1577), .A2 (B_imm[9]), .A3 (A_imm[0]));
OAI211_X1 i_1639 (.ZN (n_1575), .A (n_1578), .B (n_1579), .C1 (n_8347), .C2 (n_3554));
OAI22_X1 i_1638 (.ZN (n_1574), .A1 (n_8947), .A2 (n_3554), .B1 (n_8232), .B2 (n_6677));
OAI22_X1 i_1637 (.ZN (n_1573), .A1 (n_6577), .A2 (n_3718), .B1 (n_6584), .B2 (n_8293));
OAI22_X1 i_1636 (.ZN (n_1572), .A1 (n_7691), .A2 (n_6740), .B1 (n_6817), .B2 (n_3718));
NAND2_X1 i_1635 (.ZN (n_1571), .A1 (A_imm[4]), .A2 (B_imm[2]));
INV_X1 i_1634 (.ZN (n_1570), .A (n_1571));
NAND4_X1 i_1633 (.ZN (n_1569), .A1 (A_imm[6]), .A2 (B_imm[3]), .A3 (B_imm[0]), .A4 (A_imm[3]));
INV_X1 i_1632 (.ZN (n_1568), .A (n_1569));
OAI21_X1 i_1631 (.ZN (n_1567), .A (n_1572), .B1 (n_1568), .B2 (n_1570));
INV_X1 i_1630 (.ZN (n_1566), .A (n_1567));
NAND4_X1 i_1629 (.ZN (n_1565), .A1 (B_imm[4]), .A2 (B_imm[2]), .A3 (A_imm[5]), .A4 (A_imm[3]));
INV_X1 i_1628 (.ZN (n_1564), .A (n_1565));
OAI21_X1 i_1627 (.ZN (n_1563), .A (n_1573), .B1 (n_1566), .B2 (n_1564));
NAND4_X1 i_1626 (.ZN (n_1562), .A1 (B_imm[8]), .A2 (B_imm[6]), .A3 (A_imm[2]), .A4 (A_imm[0]));
NAND2_X1 i_1625 (.ZN (n_1561), .A1 (n_1562), .A2 (n_1563));
NAND2_X1 i_1624 (.ZN (n_1560), .A1 (n_1561), .A2 (n_1574));
INV_X1 i_1623 (.ZN (n_1559), .A (n_1560));
NAND2_X1 i_1622 (.ZN (n_1558), .A1 (n_1559), .A2 (n_1575));
NAND2_X1 i_1621 (.ZN (n_1557), .A1 (n_1558), .A2 (n_1576));
NAND2_X1 i_1620 (.ZN (n_1556), .A1 (n_1557), .A2 (n_1580));
NAND4_X1 i_1619 (.ZN (n_1555), .A1 (n_1558), .A2 (n_1582), .A3 (n_1581), .A4 (n_1576));
NAND4_X1 i_1618 (.ZN (n_1554), .A1 (n_1702), .A2 (n_1701), .A3 (n_1698), .A4 (n_1697));
NAND2_X1 i_1617 (.ZN (n_1553), .A1 (n_1701), .A2 (n_1702));
NAND2_X1 i_1616 (.ZN (n_1552), .A1 (n_1553), .A2 (n_1696));
NAND2_X1 i_1615 (.ZN (n_1551), .A1 (n_1552), .A2 (n_1554));
NAND2_X1 i_1614 (.ZN (n_1550), .A1 (n_1551), .A2 (n_1555));
NAND2_X1 i_1613 (.ZN (n_1549), .A1 (n_1550), .A2 (n_1556));
OAI21_X1 i_1612 (.ZN (n_1548), .A (n_1549), .B1 (n_1586), .B2 (n_1585));
INV_X1 i_1611 (.ZN (n_1547), .A (n_1585));
NAND4_X1 i_1610 (.ZN (n_1546), .A1 (n_1547), .A2 (n_1550), .A3 (n_1587), .A4 (n_1556));
NAND3_X1 i_1609 (.ZN (n_1545), .A1 (n_1621), .A2 (n_1620), .A3 (n_1616));
INV_X1 i_1608 (.ZN (n_1544), .A (n_1545));
AOI21_X1 i_1607 (.ZN (n_1543), .A (n_1616), .B1 (n_1621), .B2 (n_1620));
NOR2_X1 i_1606 (.ZN (n_1542), .A1 (n_1544), .A2 (n_1543));
NAND2_X1 i_1605 (.ZN (n_1541), .A1 (n_1542), .A2 (n_1546));
NAND2_X1 i_1604 (.ZN (n_1540), .A1 (n_1541), .A2 (n_1548));
NAND3_X2 i_1603 (.ZN (n_1539), .A1 (n_1588), .A2 (n_1590), .A3 (n_1540));
INV_X1 i_1602 (.ZN (n_1538), .A (n_1539));
NAND3_X1 i_1601 (.ZN (n_1537), .A1 (n_1593), .A2 (n_1592), .A3 (n_1538));
INV_X1 i_1600 (.ZN (n_1536), .A (n_1592));
OAI21_X2 i_1599 (.ZN (n_1535), .A (n_1539), .B1 (n_1604), .B2 (n_1536));
INV_X1 i_1598 (.ZN (n_1534), .A (n_1535));
NAND2_X1 i_1597 (.ZN (n_1533), .A1 (n_1590), .A2 (n_1588));
INV_X1 i_1596 (.ZN (n_1532), .A (n_1540));
NAND2_X1 i_1595 (.ZN (n_1531), .A1 (n_1533), .A2 (n_1532));
NAND2_X2 i_1594 (.ZN (n_1530), .A1 (n_1531), .A2 (n_1539));
INV_X1 i_1593 (.ZN (n_1529), .A (n_1530));
OAI211_X1 i_1592 (.ZN (n_1528), .A (n_1548), .B (n_1546), .C1 (n_1544), .C2 (n_1543));
NAND2_X1 i_1591 (.ZN (n_1527), .A1 (n_1548), .A2 (n_1546));
NAND2_X1 i_1590 (.ZN (n_1526), .A1 (n_1527), .A2 (n_1542));
AOI21_X1 i_1589 (.ZN (n_1525), .A (n_1628), .B1 (n_1632), .B2 (n_1634));
INV_X1 i_1588 (.ZN (n_1524), .A (n_1525));
NAND3_X1 i_1587 (.ZN (n_1523), .A1 (n_1632), .A2 (n_1634), .A3 (n_1628));
NAND4_X1 i_1586 (.ZN (n_1522), .A1 (B_imm[7]), .A2 (B_imm[5]), .A3 (A_imm[3]), .A4 (A_imm[1]));
INV_X1 i_1585 (.ZN (n_1521), .A (n_1522));
OAI22_X1 i_1584 (.ZN (n_1520), .A1 (n_8573), .A2 (n_6836), .B1 (n_8429), .B2 (n_3718));
NAND2_X1 i_1583 (.ZN (n_1519), .A1 (n_1761), .A2 (n_1759));
XNOR2_X1 i_1582 (.ZN (n_1518), .A (n_1519), .B (n_1760));
INV_X1 i_1581 (.ZN (n_1517), .A (n_1518));
AOI21_X1 i_1580 (.ZN (n_1516), .A (n_1521), .B1 (n_1517), .B2 (n_1520));
INV_X1 i_1579 (.ZN (n_1515), .A (n_1516));
NAND4_X1 i_1578 (.ZN (n_1514), .A1 (n_1641), .A2 (n_1642), .A3 (n_1639), .A4 (n_1638));
NAND2_X1 i_1577 (.ZN (n_1513), .A1 (n_1641), .A2 (n_1642));
NAND2_X1 i_1576 (.ZN (n_1512), .A1 (n_1513), .A2 (n_1637));
NAND2_X1 i_1575 (.ZN (n_1511), .A1 (n_1512), .A2 (n_1514));
NAND2_X1 i_1574 (.ZN (n_1510), .A1 (n_1515), .A2 (n_1511));
NAND3_X1 i_1573 (.ZN (n_1509), .A1 (n_1516), .A2 (n_1514), .A3 (n_1512));
INV_X1 i_1572 (.ZN (n_1508), .A (n_1645));
NAND2_X1 i_1571 (.ZN (n_1507), .A1 (n_1656), .A2 (n_1644));
NAND2_X1 i_1570 (.ZN (n_1506), .A1 (n_1507), .A2 (n_1508));
NAND3_X1 i_1569 (.ZN (n_1505), .A1 (n_1656), .A2 (n_1645), .A3 (n_1644));
NAND2_X1 i_1568 (.ZN (n_1504), .A1 (n_1506), .A2 (n_1505));
NAND2_X1 i_1567 (.ZN (n_1503), .A1 (n_1504), .A2 (n_1509));
NAND2_X1 i_1566 (.ZN (n_1502), .A1 (n_1503), .A2 (n_1510));
NAND3_X1 i_1565 (.ZN (n_1501), .A1 (n_1502), .A2 (n_1524), .A3 (n_1523));
INV_X1 i_1564 (.ZN (n_1500), .A (n_1523));
OAI211_X1 i_1563 (.ZN (n_1499), .A (n_1510), .B (n_1503), .C1 (n_1500), .C2 (n_1525));
NAND3_X1 i_1562 (.ZN (n_1498), .A1 (n_1556), .A2 (n_1555), .A3 (n_1551));
NAND2_X1 i_1561 (.ZN (n_1497), .A1 (n_1556), .A2 (n_1555));
NAND3_X1 i_1560 (.ZN (n_1496), .A1 (n_1497), .A2 (n_1554), .A3 (n_1552));
NAND3_X1 i_1559 (.ZN (n_1495), .A1 (n_1496), .A2 (n_1499), .A3 (n_1498));
NAND2_X1 i_1558 (.ZN (n_1494), .A1 (n_1495), .A2 (n_1501));
INV_X1 i_1557 (.ZN (n_1493), .A (n_1494));
AOI21_X1 i_1556 (.ZN (n_1492), .A (n_1493), .B1 (n_1528), .B2 (n_1526));
NAND2_X1 i_1555 (.ZN (n_1491), .A1 (n_1529), .A2 (n_1492));
INV_X1 i_1554 (.ZN (n_1490), .A (n_1491));
NAND2_X1 i_1553 (.ZN (n_1489), .A1 (n_1526), .A2 (n_1528));
NAND2_X2 i_1552 (.ZN (n_1488), .A1 (n_1489), .A2 (n_1494));
NAND3_X1 i_1551 (.ZN (n_1487), .A1 (n_1526), .A2 (n_1528), .A3 (n_1493));
NAND2_X1 i_1550 (.ZN (n_1486), .A1 (n_1576), .A2 (n_1575));
NAND2_X1 i_1549 (.ZN (n_1485), .A1 (n_1486), .A2 (n_1560));
NAND3_X1 i_1548 (.ZN (n_1484), .A1 (n_1559), .A2 (n_1576), .A3 (n_1575));
NAND2_X1 i_1547 (.ZN (n_1483), .A1 (n_1485), .A2 (n_1484));
NAND4_X1 i_1546 (.ZN (n_1482), .A1 (B_imm[7]), .A2 (B_imm[5]), .A3 (A_imm[2]), .A4 (A_imm[0]));
OAI22_X1 i_1545 (.ZN (n_1481), .A1 (n_8573), .A2 (n_3554), .B1 (n_8429), .B2 (n_6677));
INV_X1 i_1544 (.ZN (n_1480), .A (n_1481));
NAND2_X1 i_1543 (.ZN (n_1479), .A1 (n_1655), .A2 (n_1653));
XNOR2_X1 i_1542 (.ZN (n_1478), .A (n_1479), .B (n_1654));
NAND2_X1 i_1541 (.ZN (n_1477), .A1 (n_1650), .A2 (n_1649));
NAND2_X1 i_1540 (.ZN (n_1476), .A1 (n_1477), .A2 (n_1646));
NAND3_X1 i_1539 (.ZN (n_1475), .A1 (n_1650), .A2 (n_1649), .A3 (n_1647));
NAND2_X1 i_1538 (.ZN (n_1474), .A1 (n_1476), .A2 (n_1475));
INV_X1 i_1537 (.ZN (n_1473), .A (n_1474));
OAI211_X1 i_1536 (.ZN (n_1472), .A (n_1473), .B (n_1482), .C1 (n_1480), .C2 (n_1478));
OAI21_X1 i_1535 (.ZN (n_1471), .A (n_1482), .B1 (n_1478), .B2 (n_1480));
NAND2_X1 i_1534 (.ZN (n_1470), .A1 (n_1471), .A2 (n_1474));
NAND3_X1 i_1533 (.ZN (n_1469), .A1 (n_1518), .A2 (n_1522), .A3 (n_1520));
INV_X1 i_1532 (.ZN (n_1468), .A (n_1520));
OAI21_X1 i_1531 (.ZN (n_1467), .A (n_1517), .B1 (n_1521), .B2 (n_1468));
NAND2_X1 i_1530 (.ZN (n_1466), .A1 (n_1467), .A2 (n_1469));
INV_X1 i_1529 (.ZN (n_1465), .A (n_1466));
NAND2_X1 i_1528 (.ZN (n_1464), .A1 (n_1465), .A2 (n_1470));
NAND2_X1 i_1527 (.ZN (n_1463), .A1 (n_1464), .A2 (n_1472));
NAND2_X1 i_1526 (.ZN (n_1462), .A1 (n_1483), .A2 (n_1463));
NAND4_X1 i_1525 (.ZN (n_1461), .A1 (n_1485), .A2 (n_1464), .A3 (n_1484), .A4 (n_1472));
NAND2_X1 i_1524 (.ZN (n_1460), .A1 (n_1509), .A2 (n_1510));
NAND3_X1 i_1523 (.ZN (n_1459), .A1 (n_1460), .A2 (n_1506), .A3 (n_1505));
NAND3_X1 i_1522 (.ZN (n_1458), .A1 (n_1504), .A2 (n_1510), .A3 (n_1509));
NAND2_X1 i_1521 (.ZN (n_1457), .A1 (n_1459), .A2 (n_1458));
NAND2_X1 i_1520 (.ZN (n_1456), .A1 (n_1457), .A2 (n_1461));
NAND2_X1 i_1519 (.ZN (n_1455), .A1 (n_1456), .A2 (n_1462));
NAND2_X1 i_1518 (.ZN (n_1454), .A1 (n_1496), .A2 (n_1498));
NAND3_X1 i_1517 (.ZN (n_1453), .A1 (n_1454), .A2 (n_1501), .A3 (n_1499));
NAND2_X1 i_1516 (.ZN (n_1452), .A1 (n_1499), .A2 (n_1501));
NAND3_X1 i_1515 (.ZN (n_1451), .A1 (n_1452), .A2 (n_1498), .A3 (n_1496));
AOI21_X1 i_1514 (.ZN (n_1450), .A (n_1455), .B1 (n_1451), .B2 (n_1453));
NAND3_X1 i_1513 (.ZN (n_1449), .A1 (n_1488), .A2 (n_1487), .A3 (n_1450));
NAND3_X1 i_1512 (.ZN (n_1448), .A1 (n_1453), .A2 (n_1455), .A3 (n_1451));
INV_X1 i_1511 (.ZN (n_1447), .A (n_1448));
NAND4_X1 i_1510 (.ZN (n_1446), .A1 (A_imm[2]), .A2 (B_imm[1]), .A3 (B_imm[0]), .A4 (A_imm[1]));
INV_X1 i_1509 (.ZN (n_1445), .A (n_1446));
NAND2_X1 i_1508 (.ZN (n_1444), .A1 (n_1445), .A2 (B_imm[2]));
INV_X1 i_1507 (.ZN (n_1443), .A (n_1444));
NAND2_X1 i_1506 (.ZN (n_1442), .A1 (B_imm[2]), .A2 (A_imm[2]));
INV_X1 i_1505 (.ZN (n_1441), .A (n_1442));
AOI22_X1 i_1504 (.ZN (n_1440), .A1 (B_imm[3]), .A2 (A_imm[1]), .B1 (A_imm[3]), .B2 (B_imm[1]));
NAND4_X1 i_1503 (.ZN (n_1439), .A1 (B_imm[3]), .A2 (B_imm[1]), .A3 (A_imm[3]), .A4 (A_imm[1]));
INV_X1 i_1502 (.ZN (n_1438), .A (n_1439));
OAI21_X1 i_1501 (.ZN (n_1437), .A (n_1441), .B1 (n_1438), .B2 (n_1440));
INV_X1 i_1500 (.ZN (n_1436), .A (n_1440));
NAND3_X1 i_1499 (.ZN (n_1435), .A1 (n_1436), .A2 (n_1442), .A3 (n_1439));
NAND2_X1 i_1498 (.ZN (n_1434), .A1 (n_1437), .A2 (n_1435));
NAND2_X1 i_1497 (.ZN (n_1433), .A1 (n_1434), .A2 (n_1443));
AOI21_X1 i_1496 (.ZN (n_1432), .A (n_1440), .B1 (n_1442), .B2 (n_1439));
NAND3_X1 i_1495 (.ZN (n_1431), .A1 (n_1432), .A2 (B_imm[0]), .A3 (A_imm[5]));
INV_X1 i_1494 (.ZN (n_1430), .A (n_1432));
OAI21_X1 i_1493 (.ZN (n_1429), .A (n_1430), .B1 (n_6740), .B2 (n_8293));
NAND2_X1 i_1492 (.ZN (n_1428), .A1 (n_1429), .A2 (n_1431));
NAND2_X1 i_1491 (.ZN (n_1427), .A1 (B_imm[4]), .A2 (A_imm[1]));
INV_X1 i_1490 (.ZN (n_1426), .A (n_1427));
NAND2_X1 i_1489 (.ZN (n_1425), .A1 (n_1428), .A2 (n_1426));
NAND3_X1 i_1488 (.ZN (n_1424), .A1 (n_1429), .A2 (n_1431), .A3 (n_1427));
AOI21_X1 i_1487 (.ZN (n_1423), .A (n_1433), .B1 (n_1425), .B2 (n_1424));
NAND2_X1 i_1486 (.ZN (n_1422), .A1 (n_1572), .A2 (n_1569));
NAND2_X1 i_1485 (.ZN (n_1421), .A1 (n_1422), .A2 (n_1570));
NAND3_X1 i_1484 (.ZN (n_1420), .A1 (n_1572), .A2 (n_1571), .A3 (n_1569));
NAND2_X1 i_1483 (.ZN (n_1419), .A1 (n_1421), .A2 (n_1420));
NAND3_X1 i_1482 (.ZN (n_1418), .A1 (n_1419), .A2 (B_imm[5]), .A3 (A_imm[1]));
OAI211_X1 i_1481 (.ZN (n_1417), .A (n_1421), .B (n_1420), .C1 (n_8429), .C2 (n_6836));
NAND2_X1 i_1480 (.ZN (n_1416), .A1 (n_1418), .A2 (n_1417));
NAND3_X1 i_1479 (.ZN (n_1415), .A1 (n_1416), .A2 (B_imm[6]), .A3 (A_imm[0]));
OAI211_X1 i_1478 (.ZN (n_1414), .A (n_1418), .B (n_1417), .C1 (n_8232), .C2 (n_3554));
NAND2_X1 i_1477 (.ZN (n_1413), .A1 (n_1415), .A2 (n_1414));
AOI22_X1 i_1476 (.ZN (n_1412), .A1 (B_imm[4]), .A2 (A_imm[2]), .B1 (B_imm[1]), .B2 (A_imm[5]));
OAI22_X1 i_1475 (.ZN (n_1411), .A1 (n_6584), .A2 (n_3718), .B1 (n_6817), .B2 (n_6677));
NAND2_X1 i_1474 (.ZN (n_1410), .A1 (A_imm[4]), .A2 (B_imm[1]));
INV_X1 i_1473 (.ZN (n_1409), .A (n_1410));
NAND4_X1 i_1472 (.ZN (n_1408), .A1 (B_imm[2]), .A2 (B_imm[3]), .A3 (A_imm[3]), .A4 (A_imm[2]));
INV_X1 i_1471 (.ZN (n_1407), .A (n_1408));
OAI21_X1 i_1470 (.ZN (n_1406), .A (n_1411), .B1 (n_1407), .B2 (n_1409));
NAND4_X1 i_1469 (.ZN (n_1405), .A1 (B_imm[4]), .A2 (B_imm[1]), .A3 (A_imm[5]), .A4 (A_imm[2]));
AOI21_X1 i_1468 (.ZN (n_1404), .A (n_1412), .B1 (n_1406), .B2 (n_1405));
NAND3_X1 i_1467 (.ZN (n_1403), .A1 (n_1404), .A2 (B_imm[6]), .A3 (A_imm[1]));
INV_X1 i_1466 (.ZN (n_1402), .A (n_1404));
OAI21_X1 i_1465 (.ZN (n_1401), .A (n_1402), .B1 (n_8232), .B2 (n_6836));
NAND2_X1 i_1464 (.ZN (n_1400), .A1 (n_1401), .A2 (n_1403));
NAND2_X1 i_1463 (.ZN (n_1399), .A1 (n_1573), .A2 (n_1565));
XNOR2_X1 i_1462 (.ZN (n_1398), .A (n_1399), .B (n_1566));
INV_X1 i_1461 (.ZN (n_1397), .A (n_1398));
NAND2_X1 i_1460 (.ZN (n_1396), .A1 (n_1397), .A2 (n_1400));
NAND3_X1 i_1459 (.ZN (n_1395), .A1 (n_1398), .A2 (n_1403), .A3 (n_1401));
NAND4_X2 i_1458 (.ZN (n_1394), .A1 (n_1396), .A2 (n_1413), .A3 (n_1395), .A4 (n_1423));
INV_X1 i_1457 (.ZN (n_1393), .A (n_1394));
NAND3_X1 i_1456 (.ZN (n_1392), .A1 (n_1472), .A2 (n_1470), .A3 (n_1465));
NAND2_X1 i_1455 (.ZN (n_1391), .A1 (n_1472), .A2 (n_1470));
NAND2_X1 i_1454 (.ZN (n_1390), .A1 (n_1391), .A2 (n_1466));
NAND2_X1 i_1453 (.ZN (n_1389), .A1 (n_1390), .A2 (n_1392));
AOI21_X1 i_1452 (.ZN (n_1388), .A (n_1563), .B1 (n_1574), .B2 (n_1562));
NAND3_X1 i_1451 (.ZN (n_1387), .A1 (n_1574), .A2 (n_1563), .A3 (n_1562));
INV_X1 i_1450 (.ZN (n_1386), .A (n_1387));
NOR2_X1 i_1449 (.ZN (n_1385), .A1 (n_1388), .A2 (n_1386));
INV_X1 i_1448 (.ZN (n_1384), .A (n_1403));
OAI21_X1 i_1447 (.ZN (n_1383), .A (n_1401), .B1 (n_1398), .B2 (n_1384));
NAND2_X1 i_1446 (.ZN (n_1382), .A1 (n_1385), .A2 (n_1383));
INV_X1 i_1445 (.ZN (n_1381), .A (n_1383));
OAI21_X1 i_1444 (.ZN (n_1380), .A (n_1381), .B1 (n_1388), .B2 (n_1386));
NAND2_X1 i_1443 (.ZN (n_1379), .A1 (n_1481), .A2 (n_1482));
INV_X1 i_1442 (.ZN (n_1378), .A (n_1379));
NAND2_X1 i_1441 (.ZN (n_1377), .A1 (n_1478), .A2 (n_1378));
INV_X1 i_1440 (.ZN (n_1376), .A (n_1478));
NAND2_X1 i_1439 (.ZN (n_1375), .A1 (n_1376), .A2 (n_1379));
NAND2_X1 i_1438 (.ZN (n_1374), .A1 (n_1375), .A2 (n_1377));
NAND3_X1 i_1437 (.ZN (n_1373), .A1 (n_1417), .A2 (B_imm[6]), .A3 (A_imm[0]));
NAND2_X1 i_1436 (.ZN (n_1372), .A1 (n_1373), .A2 (n_1418));
NAND2_X1 i_1435 (.ZN (n_1371), .A1 (n_1374), .A2 (n_1372));
NAND4_X1 i_1434 (.ZN (n_1370), .A1 (n_1375), .A2 (n_1373), .A3 (n_1377), .A4 (n_1418));
INV_X1 i_1433 (.ZN (n_1369), .A (n_1406));
INV_X1 i_1432 (.ZN (n_1368), .A (n_1405));
OAI21_X1 i_1431 (.ZN (n_1367), .A (n_1369), .B1 (n_1368), .B2 (n_1412));
INV_X1 i_1430 (.ZN (n_1366), .A (n_1412));
NAND3_X1 i_1429 (.ZN (n_1365), .A1 (n_1366), .A2 (n_1406), .A3 (n_1405));
INV_X1 i_1428 (.ZN (n_1364), .A (n_1431));
OAI21_X1 i_1427 (.ZN (n_1363), .A (n_1429), .B1 (n_1364), .B2 (n_1426));
AOI21_X1 i_1426 (.ZN (n_1362), .A (n_1363), .B1 (n_1365), .B2 (n_1367));
NAND3_X1 i_1425 (.ZN (n_1361), .A1 (n_1363), .A2 (n_1365), .A3 (n_1367));
OAI22_X1 i_1424 (.ZN (n_1360), .A1 (n_6677), .A2 (n_4366), .B1 (n_3718), .B2 (n_6740));
NAND2_X1 i_1423 (.ZN (n_1359), .A1 (B_imm[3]), .A2 (A_imm[0]));
NAND4_X1 i_1422 (.ZN (n_1358), .A1 (A_imm[2]), .A2 (B_imm[1]), .A3 (B_imm[0]), .A4 (A_imm[3]));
NAND2_X1 i_1421 (.ZN (n_1357), .A1 (n_1358), .A2 (n_1359));
NAND2_X1 i_1420 (.ZN (n_1356), .A1 (n_1357), .A2 (n_1360));
OAI21_X1 i_1419 (.ZN (n_1355), .A (n_1356), .B1 (n_6740), .B2 (n_6678));
NAND2_X1 i_1418 (.ZN (n_1354), .A1 (B_imm[4]), .A2 (A_imm[0]));
NAND4_X1 i_1417 (.ZN (n_1353), .A1 (n_1357), .A2 (n_1360), .A3 (B_imm[0]), .A4 (A_imm[4]));
NAND2_X1 i_1416 (.ZN (n_1352), .A1 (n_1353), .A2 (n_1354));
NAND4_X1 i_1415 (.ZN (n_1351), .A1 (n_1352), .A2 (n_1355), .A3 (B_imm[5]), .A4 (A_imm[0]));
NAND2_X1 i_1414 (.ZN (n_1350), .A1 (n_1352), .A2 (n_1355));
OAI21_X1 i_1413 (.ZN (n_1349), .A (n_1350), .B1 (n_8429), .B2 (n_3554));
NAND2_X1 i_1412 (.ZN (n_1348), .A1 (n_1411), .A2 (n_1408));
XNOR2_X1 i_1411 (.ZN (n_1347), .A (n_1348), .B (n_1409));
NAND2_X1 i_1410 (.ZN (n_1346), .A1 (n_1349), .A2 (n_1347));
NAND2_X1 i_1409 (.ZN (n_1345), .A1 (n_1346), .A2 (n_1351));
AOI21_X1 i_1408 (.ZN (n_1344), .A (n_1362), .B1 (n_1345), .B2 (n_1361));
INV_X1 i_1407 (.ZN (n_1343), .A (n_1344));
NAND2_X1 i_1406 (.ZN (n_1342), .A1 (n_1343), .A2 (n_1370));
NAND3_X1 i_1405 (.ZN (n_1341), .A1 (n_1380), .A2 (n_1342), .A3 (n_1371));
NAND4_X1 i_1404 (.ZN (n_1340), .A1 (n_1389), .A2 (n_1341), .A3 (n_1393), .A4 (n_1382));
OAI21_X1 i_1403 (.ZN (n_1339), .A (n_1340), .B1 (n_1447), .B2 (n_1450));
INV_X1 i_1402 (.ZN (n_1338), .A (n_1455));
NAND2_X1 i_1401 (.ZN (n_1337), .A1 (n_1453), .A2 (n_1451));
NAND2_X1 i_1400 (.ZN (n_1336), .A1 (n_1337), .A2 (n_1338));
INV_X1 i_1399 (.ZN (n_1335), .A (n_1340));
NAND3_X1 i_1398 (.ZN (n_1334), .A1 (n_1336), .A2 (n_1448), .A3 (n_1335));
INV_X1 i_1397 (.ZN (n_1333), .A (n_1334));
AOI22_X1 i_1396 (.ZN (n_1332), .A1 (n_1341), .A2 (n_1382), .B1 (n_1389), .B2 (n_1393));
NAND2_X1 i_1395 (.ZN (n_1331), .A1 (n_1462), .A2 (n_1461));
NAND3_X1 i_1394 (.ZN (n_1330), .A1 (n_1331), .A2 (n_1459), .A3 (n_1458));
NAND3_X1 i_1393 (.ZN (n_1329), .A1 (n_1457), .A2 (n_1462), .A3 (n_1461));
OAI211_X1 i_1392 (.ZN (n_1328), .A (n_1330), .B (n_1329), .C1 (n_1335), .C2 (n_1332));
INV_X1 i_1391 (.ZN (n_1327), .A (n_1328));
INV_X1 i_1390 (.ZN (n_1326), .A (n_1332));
NAND2_X1 i_1389 (.ZN (n_1325), .A1 (n_1330), .A2 (n_1329));
NAND3_X1 i_1388 (.ZN (n_1324), .A1 (n_1325), .A2 (n_1340), .A3 (n_1326));
NAND2_X1 i_1387 (.ZN (n_1323), .A1 (n_1389), .A2 (n_1393));
NAND3_X1 i_1386 (.ZN (n_1322), .A1 (n_1390), .A2 (n_1394), .A3 (n_1392));
NAND2_X1 i_1385 (.ZN (n_1321), .A1 (n_1323), .A2 (n_1322));
NAND2_X1 i_1384 (.ZN (n_1320), .A1 (n_1342), .A2 (n_1371));
NAND3_X1 i_1383 (.ZN (n_1319), .A1 (n_1320), .A2 (n_1382), .A3 (n_1380));
NAND2_X1 i_1382 (.ZN (n_1318), .A1 (n_1380), .A2 (n_1382));
NAND3_X1 i_1381 (.ZN (n_1317), .A1 (n_1318), .A2 (n_1371), .A3 (n_1342));
NAND2_X1 i_1380 (.ZN (n_1316), .A1 (n_1317), .A2 (n_1319));
NAND2_X1 i_1379 (.ZN (n_1315), .A1 (n_1321), .A2 (n_1316));
NAND4_X1 i_1378 (.ZN (n_1314), .A1 (n_1317), .A2 (n_1319), .A3 (n_1323), .A4 (n_1322));
INV_X1 i_1377 (.ZN (n_1313), .A (n_1314));
NAND2_X1 i_1376 (.ZN (n_1312), .A1 (n_1413), .A2 (n_1423));
NAND2_X1 i_1375 (.ZN (n_1311), .A1 (n_1395), .A2 (n_1396));
NAND2_X1 i_1374 (.ZN (n_1310), .A1 (n_1311), .A2 (n_1312));
NAND3_X1 i_1373 (.ZN (n_1309), .A1 (n_1343), .A2 (n_1371), .A3 (n_1370));
NAND2_X1 i_1372 (.ZN (n_1308), .A1 (n_1371), .A2 (n_1370));
NAND2_X1 i_1371 (.ZN (n_1307), .A1 (n_1308), .A2 (n_1344));
NAND4_X1 i_1370 (.ZN (n_1306), .A1 (n_1310), .A2 (n_1307), .A3 (n_1309), .A4 (n_1394));
INV_X1 i_1369 (.ZN (n_1305), .A (n_1423));
NAND3_X1 i_1368 (.ZN (n_1304), .A1 (n_1305), .A2 (n_1415), .A3 (n_1414));
NAND2_X1 i_1367 (.ZN (n_1303), .A1 (n_1312), .A2 (n_1304));
INV_X1 i_1366 (.ZN (n_1302), .A (n_1362));
NAND3_X1 i_1365 (.ZN (n_1301), .A1 (n_1302), .A2 (n_1361), .A3 (n_1345));
INV_X1 i_1364 (.ZN (n_1300), .A (n_1361));
OAI211_X1 i_1363 (.ZN (n_1299), .A (n_1351), .B (n_1346), .C1 (n_1362), .C2 (n_1300));
NAND2_X1 i_1362 (.ZN (n_1298), .A1 (n_1299), .A2 (n_1301));
NAND2_X1 i_1361 (.ZN (n_1297), .A1 (n_1303), .A2 (n_1298));
NAND4_X1 i_1360 (.ZN (n_1296), .A1 (n_1312), .A2 (n_1301), .A3 (n_1299), .A4 (n_1304));
NAND3_X1 i_1359 (.ZN (n_1295), .A1 (n_1425), .A2 (n_1433), .A3 (n_1424));
INV_X1 i_1358 (.ZN (n_1294), .A (n_1295));
INV_X1 i_1357 (.ZN (n_1293), .A (n_1347));
NAND2_X1 i_1356 (.ZN (n_1292), .A1 (n_1349), .A2 (n_1351));
NAND2_X1 i_1355 (.ZN (n_1291), .A1 (n_1292), .A2 (n_1293));
NAND3_X1 i_1354 (.ZN (n_1290), .A1 (n_1349), .A2 (n_1347), .A3 (n_1351));
NAND2_X1 i_1353 (.ZN (n_1289), .A1 (n_1291), .A2 (n_1290));
OAI21_X1 i_1352 (.ZN (n_1288), .A (n_1289), .B1 (n_1423), .B2 (n_1294));
NAND4_X1 i_1351 (.ZN (n_1287), .A1 (n_1291), .A2 (n_1305), .A3 (n_1295), .A4 (n_1290));
XNOR2_X1 i_1350 (.ZN (n_1286), .A (n_1434), .B (n_1443));
INV_X1 i_1349 (.ZN (n_1285), .A (n_1286));
INV_X1 i_1348 (.ZN (n_1284), .A (n_1354));
NAND2_X1 i_1347 (.ZN (n_1283), .A1 (n_1355), .A2 (n_1353));
XNOR2_X1 i_1346 (.ZN (n_1282), .A (n_1283), .B (n_1284));
OR2_X1 i_1345 (.ZN (n_1281), .A1 (n_1282), .A2 (n_1285));
NAND2_X1 i_1344 (.ZN (n_1280), .A1 (n_1282), .A2 (n_1285));
OAI21_X1 i_1343 (.ZN (n_1279), .A (n_1446), .B1 (n_6584), .B2 (n_6836));
NAND2_X1 i_1342 (.ZN (n_1278), .A1 (n_1279), .A2 (n_1444));
INV_X1 i_1341 (.ZN (n_1277), .A (n_1278));
INV_X1 i_1340 (.ZN (n_1276), .A (n_1359));
NAND2_X1 i_1339 (.ZN (n_1275), .A1 (n_1360), .A2 (n_1358));
XNOR2_X1 i_1338 (.ZN (n_1274), .A (n_1275), .B (n_1276));
OR2_X1 i_1337 (.ZN (n_1273), .A1 (n_1274), .A2 (n_1277));
NAND2_X1 i_1336 (.ZN (n_1272), .A1 (n_1274), .A2 (n_1277));
NAND4_X1 i_1335 (.ZN (n_1271), .A1 (A_imm[1]), .A2 (B_imm[1]), .A3 (B_imm[0]), .A4 (A_imm[0]));
OAI21_X1 i_1334 (.ZN (n_1270), .A (n_1271), .B1 (n_6584), .B2 (n_3554));
INV_X1 i_1333 (.ZN (n_1269), .A (n_1271));
NAND2_X1 i_1332 (.ZN (n_1268), .A1 (B_imm[2]), .A2 (n_1269));
INV_X1 i_1331 (.ZN (n_1267), .A (n_1268));
AOI22_X1 i_1330 (.ZN (n_1266), .A1 (A_imm[2]), .A2 (B_imm[0]), .B1 (B_imm[1]), .B2 (A_imm[1]));
NOR2_X1 i_1329 (.ZN (n_1265), .A1 (n_1445), .A2 (n_1266));
OAI21_X1 i_1328 (.ZN (n_1264), .A (n_1270), .B1 (n_1265), .B2 (n_1267));
NAND2_X1 i_1327 (.ZN (n_1263), .A1 (n_1272), .A2 (n_1264));
NAND2_X1 i_1326 (.ZN (n_1262), .A1 (n_1273), .A2 (n_1263));
NAND2_X1 i_1325 (.ZN (n_1261), .A1 (n_1280), .A2 (n_1262));
NAND2_X1 i_1324 (.ZN (n_1260), .A1 (n_1281), .A2 (n_1261));
NAND2_X1 i_1323 (.ZN (n_1259), .A1 (n_1260), .A2 (n_1287));
NAND2_X1 i_1322 (.ZN (n_1258), .A1 (n_1259), .A2 (n_1288));
NAND2_X1 i_1321 (.ZN (n_1257), .A1 (n_1258), .A2 (n_1296));
NAND2_X1 i_1320 (.ZN (n_1256), .A1 (n_1257), .A2 (n_1297));
NAND2_X1 i_1319 (.ZN (n_1255), .A1 (n_1310), .A2 (n_1394));
NAND2_X1 i_1318 (.ZN (n_1254), .A1 (n_1309), .A2 (n_1307));
NAND2_X1 i_1317 (.ZN (n_1253), .A1 (n_1254), .A2 (n_1255));
INV_X1 i_1316 (.ZN (n_1252), .A (n_1253));
AOI21_X1 i_1315 (.ZN (n_1251), .A (n_1252), .B1 (n_1256), .B2 (n_1306));
OAI21_X2 i_1314 (.ZN (n_1250), .A (n_1315), .B1 (n_1251), .B2 (n_1313));
AOI21_X2 i_1313 (.ZN (n_1249), .A (n_1327), .B1 (n_1250), .B2 (n_1324));
OAI21_X2 i_1312 (.ZN (n_1248), .A (n_1339), .B1 (n_1333), .B2 (n_1249));
NAND2_X2 i_1311 (.ZN (n_1247), .A1 (n_1248), .A2 (n_1449));
AOI21_X1 i_1310 (.ZN (n_1246), .A (n_1450), .B1 (n_1488), .B2 (n_1487));
AOI21_X2 i_1309 (.ZN (n_1245), .A (n_1246), .B1 (n_1530), .B2 (n_1488));
AOI21_X4 i_1308 (.ZN (n_1244), .A (n_1490), .B1 (n_1245), .B2 (n_1247));
OAI211_X2 i_1307 (.ZN (n_1243), .A (n_1594), .B (n_1537), .C1 (n_1244), .C2 (n_1534));
NAND3_X1 i_1306 (.ZN (n_1242), .A1 (n_1788), .A2 (n_1793), .A3 (n_1721));
INV_X1 i_1305 (.ZN (n_1241), .A (n_1242));
OAI21_X1 i_1304 (.ZN (n_1240), .A (n_1598), .B1 (n_1241), .B2 (n_1720));
NAND2_X1 i_1303 (.ZN (n_1239), .A1 (n_1595), .A2 (n_1598));
NAND2_X1 i_1302 (.ZN (n_1238), .A1 (n_1239), .A2 (n_1593));
NAND2_X1 i_1301 (.ZN (n_1237), .A1 (n_1240), .A2 (n_1238));
INV_X1 i_1300 (.ZN (n_1236), .A (n_1237));
NAND2_X2 i_1299 (.ZN (n_1235), .A1 (n_1243), .A2 (n_1236));
INV_X1 i_1298 (.ZN (n_1234), .A (n_1598));
NAND3_X1 i_1297 (.ZN (n_1233), .A1 (n_1719), .A2 (n_1234), .A3 (n_1242));
NAND2_X1 i_1296 (.ZN (n_1232), .A1 (n_1897), .A2 (n_1892));
INV_X1 i_1295 (.ZN (n_1231), .A (n_1797));
NAND2_X1 i_1294 (.ZN (n_1230), .A1 (n_1232), .A2 (n_1231));
NAND3_X1 i_1293 (.ZN (n_1229), .A1 (n_1230), .A2 (n_1796), .A3 (n_1720));
NAND2_X1 i_1292 (.ZN (n_1228), .A1 (n_1229), .A2 (n_1233));
INV_X1 i_1291 (.ZN (n_1227), .A (n_1228));
AOI21_X4 i_1290 (.ZN (n_1226), .A (n_1717), .B1 (n_1235), .B2 (n_1227));
NAND2_X1 i_1289 (.ZN (n_1225), .A1 (n_2207), .A2 (n_2210));
INV_X1 i_1288 (.ZN (n_1224), .A (n_2107));
NAND2_X1 i_1287 (.ZN (n_1223), .A1 (n_1225), .A2 (n_1224));
NAND3_X1 i_1286 (.ZN (n_1222), .A1 (n_2107), .A2 (n_2210), .A3 (n_2207));
NAND3_X1 i_1285 (.ZN (n_1221), .A1 (n_2108), .A2 (n_2114), .A3 (n_2112));
NAND2_X1 i_1284 (.ZN (n_1220), .A1 (n_2112), .A2 (n_2114));
NAND3_X2 i_1283 (.ZN (n_1219), .A1 (n_1220), .A2 (n_2111), .A3 (n_2109));
NAND3_X1 i_1282 (.ZN (n_1218), .A1 (n_2252), .A2 (n_2251), .A3 (n_2249));
INV_X1 i_1281 (.ZN (n_1217), .A (n_2251));
INV_X1 i_1280 (.ZN (n_1216), .A (n_2249));
OAI21_X1 i_1279 (.ZN (n_1215), .A (n_1216), .B1 (n_2253), .B2 (n_1217));
NAND2_X1 i_1278 (.ZN (n_1214), .A1 (n_1215), .A2 (n_1218));
INV_X1 i_1277 (.ZN (n_1213), .A (n_1214));
NAND2_X1 i_1276 (.ZN (n_1212), .A1 (n_1956), .A2 (n_1954));
NAND3_X1 i_1275 (.ZN (n_1211), .A1 (n_2409), .A2 (n_2410), .A3 (n_2377));
INV_X1 i_1274 (.ZN (n_1210), .A (n_1211));
AOI21_X1 i_1273 (.ZN (n_1209), .A (n_2377), .B1 (n_2410), .B2 (n_2409));
NOR2_X1 i_1272 (.ZN (n_1208), .A1 (n_1210), .A2 (n_1209));
NAND3_X1 i_1271 (.ZN (n_1207), .A1 (n_1212), .A2 (n_1208), .A3 (n_1958));
INV_X1 i_1270 (.ZN (n_1206), .A (n_1209));
AOI22_X1 i_1269 (.ZN (n_1205), .A1 (n_1212), .A2 (n_1958), .B1 (n_1211), .B2 (n_1206));
NAND3_X1 i_1268 (.ZN (n_1204), .A1 (n_2255), .A2 (n_2290), .A3 (n_2289));
INV_X1 i_1267 (.ZN (n_1203), .A (n_2255));
NAND2_X1 i_1266 (.ZN (n_1202), .A1 (n_2290), .A2 (n_2289));
NAND2_X1 i_1265 (.ZN (n_1201), .A1 (n_1202), .A2 (n_1203));
NAND2_X1 i_1264 (.ZN (n_1200), .A1 (n_1201), .A2 (n_1204));
OAI21_X1 i_1263 (.ZN (n_1199), .A (n_1207), .B1 (n_1205), .B2 (n_1200));
NAND2_X1 i_1262 (.ZN (n_1198), .A1 (n_1213), .A2 (n_1199));
INV_X1 i_1261 (.ZN (n_1197), .A (n_1199));
NAND2_X1 i_1260 (.ZN (n_1196), .A1 (n_1214), .A2 (n_1197));
INV_X1 i_1259 (.ZN (n_1195), .A (n_1196));
INV_X1 i_1258 (.ZN (n_1194), .A (n_2121));
NAND3_X1 i_1257 (.ZN (n_1193), .A1 (n_2127), .A2 (n_1194), .A3 (n_2125));
AOI21_X1 i_1256 (.ZN (n_1192), .A (n_2126), .B1 (n_2132), .B2 (n_2141));
INV_X1 i_1255 (.ZN (n_1191), .A (n_2125));
OAI21_X1 i_1254 (.ZN (n_1190), .A (n_2121), .B1 (n_1192), .B2 (n_1191));
NAND2_X1 i_1253 (.ZN (n_1189), .A1 (n_1193), .A2 (n_1190));
INV_X1 i_1252 (.ZN (n_1188), .A (n_1189));
OAI21_X2 i_1251 (.ZN (n_1187), .A (n_1198), .B1 (n_1188), .B2 (n_1195));
NAND3_X2 i_1250 (.ZN (n_1186), .A1 (n_1187), .A2 (n_1219), .A3 (n_1221));
INV_X1 i_1249 (.ZN (n_1185), .A (n_1186));
AOI21_X1 i_1248 (.ZN (n_1184), .A (n_1185), .B1 (n_1223), .B2 (n_1222));
NAND2_X1 i_1247 (.ZN (n_1183), .A1 (n_1198), .A2 (n_1196));
NAND2_X1 i_1246 (.ZN (n_1182), .A1 (n_1183), .A2 (n_1188));
NAND3_X1 i_1245 (.ZN (n_1181), .A1 (n_1189), .A2 (n_1196), .A3 (n_1198));
NAND3_X1 i_1244 (.ZN (n_1180), .A1 (n_2141), .A2 (n_2139), .A3 (n_2134));
AOI21_X1 i_1243 (.ZN (n_1179), .A (n_2140), .B1 (n_2143), .B2 (n_2176));
INV_X1 i_1242 (.ZN (n_1178), .A (n_2139));
OAI21_X1 i_1241 (.ZN (n_1177), .A (n_2133), .B1 (n_1179), .B2 (n_1178));
NAND2_X1 i_1240 (.ZN (n_1176), .A1 (n_1177), .A2 (n_1180));
NAND2_X1 i_1239 (.ZN (n_1175), .A1 (n_2021), .A2 (n_2019));
NAND2_X1 i_1238 (.ZN (n_1174), .A1 (n_1175), .A2 (n_2022));
NAND2_X1 i_1237 (.ZN (n_1173), .A1 (n_1174), .A2 (n_1176));
NAND4_X1 i_1236 (.ZN (n_1172), .A1 (n_1175), .A2 (n_1177), .A3 (n_2022), .A4 (n_1180));
NAND2_X1 i_1235 (.ZN (n_1171), .A1 (n_1212), .A2 (n_1958));
OAI21_X1 i_1234 (.ZN (n_1170), .A (n_1171), .B1 (n_1210), .B2 (n_1209));
NAND3_X1 i_1233 (.ZN (n_1169), .A1 (n_1170), .A2 (n_1207), .A3 (n_1200));
INV_X1 i_1232 (.ZN (n_1168), .A (n_1207));
INV_X1 i_1231 (.ZN (n_1167), .A (n_1200));
OAI21_X1 i_1230 (.ZN (n_1166), .A (n_1167), .B1 (n_1168), .B2 (n_1205));
NAND2_X1 i_1229 (.ZN (n_1165), .A1 (n_1166), .A2 (n_1169));
NAND2_X1 i_1228 (.ZN (n_1164), .A1 (n_1165), .A2 (n_1172));
NAND2_X1 i_1227 (.ZN (n_1163), .A1 (n_1164), .A2 (n_1173));
NAND3_X2 i_1226 (.ZN (n_1162), .A1 (n_1182), .A2 (n_1181), .A3 (n_1163));
INV_X1 i_1225 (.ZN (n_1161), .A (n_1162));
NAND2_X1 i_1224 (.ZN (n_1160), .A1 (n_1221), .A2 (n_1219));
INV_X1 i_1223 (.ZN (n_1159), .A (n_1187));
NAND2_X1 i_1222 (.ZN (n_1158), .A1 (n_1160), .A2 (n_1159));
AOI21_X1 i_1221 (.ZN (n_1157), .A (n_1161), .B1 (n_1158), .B2 (n_1186));
NOR2_X1 i_1220 (.ZN (n_1156), .A1 (n_1184), .A2 (n_1157));
NAND2_X1 i_1219 (.ZN (n_1155), .A1 (n_1182), .A2 (n_1181));
INV_X1 i_1218 (.ZN (n_1154), .A (n_1163));
NAND2_X1 i_1217 (.ZN (n_1153), .A1 (n_1155), .A2 (n_1154));
NAND3_X1 i_1216 (.ZN (n_1152), .A1 (n_1165), .A2 (n_1173), .A3 (n_1172));
INV_X1 i_1215 (.ZN (n_1151), .A (n_1165));
NAND2_X1 i_1214 (.ZN (n_1150), .A1 (n_1173), .A2 (n_1172));
NAND2_X1 i_1213 (.ZN (n_1149), .A1 (n_1150), .A2 (n_1151));
INV_X1 i_1212 (.ZN (n_1148), .A (n_1898));
OAI21_X1 i_1211 (.ZN (n_1147), .A (n_1900), .B1 (n_1894), .B2 (n_1148));
NAND3_X2 i_1210 (.ZN (n_1146), .A1 (n_1147), .A2 (n_1149), .A3 (n_1152));
INV_X2 i_1209 (.ZN (n_1145), .A (n_1146));
AOI21_X1 i_1208 (.ZN (n_1144), .A (n_1145), .B1 (n_1153), .B2 (n_1162));
NAND2_X1 i_1207 (.ZN (n_1143), .A1 (n_1149), .A2 (n_1152));
INV_X1 i_1206 (.ZN (n_1142), .A (n_1147));
NAND2_X1 i_1205 (.ZN (n_1141), .A1 (n_1143), .A2 (n_1142));
AOI21_X1 i_1204 (.ZN (n_1140), .A (n_1795), .B1 (n_1141), .B2 (n_1146));
NOR2_X1 i_1203 (.ZN (n_1139), .A1 (n_1144), .A2 (n_1140));
NAND3_X2 i_1202 (.ZN (n_1138), .A1 (n_1226), .A2 (n_1156), .A3 (n_1139));
INV_X2 i_1201 (.ZN (n_1137), .A (n_1138));
NAND3_X4 i_1200 (.ZN (n_1136), .A1 (n_2323), .A2 (n_2104), .A3 (n_1137));
NAND3_X4 i_1198 (.ZN (n_1134), .A1 (CLOCK_opt_ipo_n333), .A2 (n_3077), .A3 (CLOCK_opt_ipo_n418));
AOI21_X1 i_1197 (.ZN (n_1133), .A (n_1187), .B1 (n_1221), .B2 (n_1219));
OAI21_X1 i_1196 (.ZN (n_1132), .A (n_1186), .B1 (n_1133), .B2 (n_1162));
NAND3_X1 i_1195 (.ZN (n_1131), .A1 (n_1132), .A2 (n_1223), .A3 (n_1222));
INV_X1 i_1194 (.ZN (n_1130), .A (n_1222));
OAI21_X1 i_1193 (.ZN (n_1129), .A (n_1186), .B1 (n_1130), .B2 (n_2106));
OAI21_X2 i_1192 (.ZN (n_1128), .A (n_1162), .B1 (n_1185), .B2 (n_1133));
NAND2_X1 i_1191 (.ZN (n_1127), .A1 (n_1153), .A2 (n_1162));
AOI21_X1 i_1190 (.ZN (n_1126), .A (n_1145), .B1 (n_1795), .B2 (n_1141));
NOR2_X1 i_1189 (.ZN (n_1125), .A1 (n_1127), .A2 (n_1126));
NAND3_X2 i_1188 (.ZN (n_1124), .A1 (n_1129), .A2 (n_1125), .A3 (n_1128));
NAND2_X2 i_1187 (.ZN (n_1123), .A1 (n_1124), .A2 (n_1131));
NAND4_X2 i_1186 (.ZN (n_1122), .A1 (n_1123), .A2 (n_2104), .A3 (n_2328), .A4 (n_2325));
NOR2_X1 i_1185 (.ZN (n_1121), .A1 (CLOCK_opt_ipo_n423), .A2 (n_2636));
OAI21_X1 i_1184 (.ZN (n_1120), .A (n_2333), .B1 (n_2329), .B2 (n_2339));
NAND2_X1 i_1183 (.ZN (n_1119), .A1 (n_1120), .A2 (n_1121));
NAND2_X1 i_1182 (.ZN (n_1118), .A1 (n_2339), .A2 (n_2216));
INV_X1 i_1181 (.ZN (n_1117), .A (n_1118));
NAND3_X1 i_1180 (.ZN (n_1116), .A1 (n_2212), .A2 (n_2218), .A3 (n_2106));
NAND2_X1 i_1179 (.ZN (n_1115), .A1 (n_1116), .A2 (n_2218));
NAND4_X2 i_1178 (.ZN (n_1114), .A1 (n_2325), .A2 (n_2328), .A3 (n_1117), .A4 (n_1115));
NAND3_X2 i_1177 (.ZN (n_1113), .A1 (n_1122), .A2 (n_1119), .A3 (n_1114));
NAND3_X1 i_1176 (.ZN (n_1112), .A1 (n_1113), .A2 (CLOCK_opt_ipo_n333), .A3 (n_3077));
INV_X1 i_1175 (.ZN (n_1111), .A (n_2929));
INV_X1 i_1174 (.ZN (n_1110), .A (n_2633));
OAI21_X1 i_1173 (.ZN (n_1109), .A (n_2774), .B1 (n_2635), .B2 (n_1110));
NAND4_X1 i_1172 (.ZN (n_1108), .A1 (n_1111), .A2 (n_1109), .A3 (n_2931), .A4 (n_2771));
INV_X2 i_1171 (.ZN (n_1107), .A (n_1108));
INV_X1 i_1170 (.ZN (n_1106), .A (n_3135));
NAND3_X1 i_1169 (.ZN (n_1105), .A1 (n_3082), .A2 (n_1106), .A3 (n_3079));
NAND3_X1 i_1168 (.ZN (n_1104), .A1 (n_2932), .A2 (n_3135), .A3 (n_2930));
NAND2_X1 i_1167 (.ZN (n_1103), .A1 (n_1105), .A2 (n_1104));
OAI21_X4 i_1166 (.ZN (n_1102), .A (n_3077), .B1 (n_1107), .B2 (n_1103));
NAND3_X4 i_1165 (.ZN (n_1101), .A1 (n_1112), .A2 (n_1102), .A3 (n_1134));
NAND4_X1 i_1164 (.ZN (n_1100), .A1 (n_4097), .A2 (n_4025), .A3 (n_4034), .A4 (n_4026));
NAND2_X1 i_1163 (.ZN (n_1099), .A1 (n_4026), .A2 (n_4034));
NAND2_X1 i_1162 (.ZN (n_1098), .A1 (n_4097), .A2 (n_4025));
NAND2_X1 i_1161 (.ZN (n_1097), .A1 (n_1098), .A2 (n_1099));
NAND2_X1 i_1160 (.ZN (n_1096), .A1 (n_1097), .A2 (n_1100));
NAND2_X1 i_1159 (.ZN (n_1095), .A1 (n_3106), .A2 (n_3098));
NAND3_X1 i_1158 (.ZN (n_1094), .A1 (n_1096), .A2 (n_3103), .A3 (n_1095));
NAND2_X1 i_1157 (.ZN (n_1093), .A1 (n_1095), .A2 (n_3103));
NAND3_X1 i_1156 (.ZN (n_1092), .A1 (n_1093), .A2 (n_1100), .A3 (n_1097));
NAND3_X1 i_1155 (.ZN (n_1091), .A1 (n_4730), .A2 (n_4728), .A3 (n_4669));
NAND2_X1 i_1154 (.ZN (n_1090), .A1 (n_4730), .A2 (n_4728));
NAND2_X1 i_1153 (.ZN (n_1089), .A1 (n_1090), .A2 (n_4670));
NAND2_X1 i_1152 (.ZN (n_1088), .A1 (n_1089), .A2 (n_1091));
NAND2_X1 i_1151 (.ZN (n_1087), .A1 (n_3128), .A2 (n_3122));
NAND3_X1 i_1150 (.ZN (n_1086), .A1 (n_1087), .A2 (n_3124), .A3 (n_1088));
INV_X1 i_1149 (.ZN (n_1085), .A (n_1088));
NAND2_X1 i_1148 (.ZN (n_1084), .A1 (n_1087), .A2 (n_3124));
NAND2_X1 i_1147 (.ZN (n_1083), .A1 (n_1084), .A2 (n_1085));
AOI21_X1 i_1146 (.ZN (n_1082), .A (n_4432), .B1 (n_4474), .B2 (n_4473));
INV_X1 i_1145 (.ZN (n_1081), .A (n_4315));
NOR2_X1 i_1144 (.ZN (n_1080), .A1 (n_1081), .A2 (n_1082));
NAND3_X1 i_1143 (.ZN (n_1079), .A1 (n_4320), .A2 (n_1080), .A3 (n_4319));
INV_X1 i_1142 (.ZN (n_1078), .A (n_1079));
AOI22_X1 i_1141 (.ZN (n_1077), .A1 (n_4320), .A2 (n_4319), .B1 (n_4316), .B2 (n_4315));
NOR2_X1 i_1140 (.ZN (n_1076), .A1 (n_1078), .A2 (n_1077));
INV_X1 i_1139 (.ZN (n_1075), .A (n_1076));
NAND3_X1 i_1138 (.ZN (n_1074), .A1 (n_1083), .A2 (n_1075), .A3 (n_1086));
INV_X1 i_1137 (.ZN (n_1073), .A (n_1086));
AOI21_X1 i_1136 (.ZN (n_1072), .A (n_1088), .B1 (n_1087), .B2 (n_3124));
OAI21_X1 i_1135 (.ZN (n_1071), .A (n_1076), .B1 (n_1073), .B2 (n_1072));
NAND2_X1 i_1134 (.ZN (n_1070), .A1 (n_1071), .A2 (n_1074));
NAND3_X1 i_1133 (.ZN (n_1069), .A1 (n_1070), .A2 (n_1094), .A3 (n_1092));
NAND2_X1 i_1132 (.ZN (n_1068), .A1 (n_1092), .A2 (n_1094));
INV_X1 i_1131 (.ZN (n_1067), .A (n_1070));
NAND2_X1 i_1130 (.ZN (n_1066), .A1 (n_1068), .A2 (n_1067));
INV_X1 i_1129 (.ZN (n_1065), .A (n_3115));
OAI21_X1 i_1128 (.ZN (n_1064), .A (n_3112), .B1 (n_3088), .B2 (n_1065));
NAND3_X1 i_1127 (.ZN (n_1063), .A1 (n_1066), .A2 (n_1064), .A3 (n_1069));
INV_X2 i_1126 (.ZN (n_1062), .A (n_1063));
AOI21_X1 i_1125 (.ZN (n_1061), .A (n_1064), .B1 (n_1066), .B2 (n_1069));
OAI21_X1 i_1124 (.ZN (n_1060), .A (n_3082), .B1 (n_1062), .B2 (n_1061));
NAND4_X1 i_1123 (.ZN (n_1059), .A1 (n_4214), .A2 (n_4216), .A3 (n_4007), .A4 (n_4000));
NAND2_X2 i_1122 (.ZN (n_1058), .A1 (n_3998), .A2 (n_1059));
NAND3_X1 i_1121 (.ZN (n_1057), .A1 (n_4001), .A2 (n_4007), .A3 (n_4006));
INV_X1 i_1120 (.ZN (n_1056), .A (n_4001));
NAND2_X1 i_1119 (.ZN (n_1055), .A1 (n_4006), .A2 (n_4007));
NAND2_X1 i_1118 (.ZN (n_1054), .A1 (n_1055), .A2 (n_1056));
NAND3_X1 i_1117 (.ZN (n_1053), .A1 (n_4313), .A2 (n_4394), .A3 (n_4392));
INV_X1 i_1116 (.ZN (n_1052), .A (n_4313));
NAND2_X1 i_1115 (.ZN (n_1051), .A1 (n_4394), .A2 (n_4392));
NAND2_X1 i_1114 (.ZN (n_1050), .A1 (n_1051), .A2 (n_1052));
NAND2_X2 i_1113 (.ZN (n_1049), .A1 (n_1050), .A2 (n_1053));
INV_X1 i_1112 (.ZN (n_1048), .A (n_1049));
NAND2_X1 i_1111 (.ZN (n_1047), .A1 (n_1086), .A2 (n_1076));
NAND2_X1 i_1110 (.ZN (n_1046), .A1 (n_1047), .A2 (n_1083));
NAND2_X2 i_1109 (.ZN (n_1045), .A1 (n_1046), .A2 (n_1048));
NAND3_X1 i_1108 (.ZN (n_1044), .A1 (n_1049), .A2 (n_1047), .A3 (n_1083));
NAND3_X1 i_1107 (.ZN (n_1043), .A1 (n_4022), .A2 (n_4021), .A3 (n_4016));
INV_X1 i_1106 (.ZN (n_1042), .A (n_1043));
AOI21_X1 i_1105 (.ZN (n_1041), .A (n_4016), .B1 (n_4022), .B2 (n_4021));
OAI21_X1 i_1104 (.ZN (n_1040), .A (n_1044), .B1 (n_1042), .B2 (n_1041));
NAND2_X1 i_1103 (.ZN (n_1039), .A1 (n_1040), .A2 (n_1045));
NAND3_X2 i_1102 (.ZN (n_1038), .A1 (n_1054), .A2 (n_1039), .A3 (n_1057));
NAND2_X1 i_1101 (.ZN (n_1037), .A1 (n_1058), .A2 (n_1038));
OAI211_X1 i_1100 (.ZN (n_1036), .A (n_1045), .B (n_1044), .C1 (n_1042), .C2 (n_1041));
AOI21_X1 i_1099 (.ZN (n_1035), .A (n_4209), .B1 (n_4097), .B2 (n_4024));
INV_X1 i_1098 (.ZN (n_1034), .A (n_4021));
OAI21_X1 i_1097 (.ZN (n_1033), .A (n_4015), .B1 (n_1035), .B2 (n_1034));
NAND2_X1 i_1096 (.ZN (n_1032), .A1 (n_1045), .A2 (n_1044));
NAND3_X2 i_1095 (.ZN (n_1031), .A1 (n_1032), .A2 (n_1043), .A3 (n_1033));
NAND2_X1 i_1094 (.ZN (n_1030), .A1 (n_1070), .A2 (n_1094));
NAND2_X1 i_1093 (.ZN (n_1029), .A1 (n_1030), .A2 (n_1092));
NAND3_X2 i_1092 (.ZN (n_1028), .A1 (n_1031), .A2 (n_1029), .A3 (n_1036));
NAND2_X1 i_1091 (.ZN (n_1027), .A1 (n_1031), .A2 (n_1036));
INV_X1 i_1090 (.ZN (n_1026), .A (n_1029));
NAND2_X1 i_1089 (.ZN (n_1025), .A1 (n_1027), .A2 (n_1026));
AOI21_X2 i_1088 (.ZN (n_1024), .A (n_1062), .B1 (n_1025), .B2 (n_1028));
INV_X2 i_1087 (.ZN (n_1023), .A (n_1028));
NAND2_X1 i_1086 (.ZN (n_1022), .A1 (n_1054), .A2 (n_1057));
INV_X1 i_1085 (.ZN (n_1021), .A (n_1039));
NAND2_X1 i_1084 (.ZN (n_1020), .A1 (n_1022), .A2 (n_1021));
AOI21_X2 i_1083 (.ZN (n_1019), .A (n_1023), .B1 (n_1020), .B2 (n_1038));
NOR2_X2 i_1082 (.ZN (n_1018), .A1 (n_1019), .A2 (n_1024));
NAND3_X1 i_1081 (.ZN (n_1017), .A1 (n_1018), .A2 (n_1060), .A3 (n_1037));
INV_X1 i_1080 (.ZN (n_1016), .A (n_1017));
NAND2_X4 i_1079 (.ZN (n_1015), .A1 (n_1101), .A2 (n_1016));
INV_X1 i_1078 (.ZN (n_1014), .A (n_1061));
NAND3_X1 i_1077 (.ZN (n_1013), .A1 (n_1014), .A2 (n_3081), .A3 (n_1063));
INV_X2 i_1076 (.ZN (n_1012), .A (n_1013));
NAND3_X1 i_1075 (.ZN (n_1011), .A1 (n_1018), .A2 (n_1037), .A3 (n_1012));
INV_X1 i_1074 (.ZN (n_1010), .A (n_1058));
NAND3_X1 i_1073 (.ZN (n_1009), .A1 (n_1025), .A2 (n_1062), .A3 (n_1028));
NAND2_X1 i_1072 (.ZN (n_1008), .A1 (n_1009), .A2 (n_1028));
OAI21_X2 sgo__sro_c303 (.ZN (n_1856), .A (sgo__sro_n156), .B1 (n_6584), .B2 (n_8644));
INV_X1 i_1070 (.ZN (n_1006), .A (n_1038));
NAND2_X1 i_1069 (.ZN (n_1005), .A1 (n_1010), .A2 (n_1006));
NAND3_X1 i_1068 (.ZN (n_1004), .A1 (n_1011), .A2 (n_1007), .A3 (n_1005));
INV_X2 i_1067 (.ZN (n_1003), .A (n_1004));
NAND2_X4 i_1066 (.ZN (n_1002), .A1 (n_1003), .A2 (n_1015));
NAND2_X1 i_1065 (.ZN (n_1001), .A1 (n_3993), .A2 (n_3996));
NAND2_X1 i_1064 (.ZN (n_1000), .A1 (n_1001), .A2 (n_3998));
NAND3_X1 i_1063 (.ZN (n_999), .A1 (n_4221), .A2 (n_1000), .A3 (n_4252));
NAND2_X2 i_1061 (.ZN (n_997), .A1 (CLOCK_opt_ipo_n326), .A2 (n_5109));
NAND2_X2 i_1059 (.ZN (n_995), .A1 (n_1002), .A2 (CLOCK_opt_ipo_n324));
INV_X1 i_1058 (.ZN (n_994), .A (n_6010));
OAI21_X2 i_1057 (.ZN (n_993), .A (n_5726), .B1 (n_994), .B2 (n_6009));
NAND2_X1 i_1056 (.ZN (n_992), .A1 (n_5692), .A2 (n_5695));
NAND2_X1 i_1055 (.ZN (n_991), .A1 (n_5690), .A2 (n_6089));
NAND2_X1 i_1054 (.ZN (n_990), .A1 (n_992), .A2 (n_991));
NAND2_X2 i_1053 (.ZN (n_989), .A1 (n_993), .A2 (n_990));
INV_X2 i_1052 (.ZN (n_988), .A (n_5666));
INV_X1 i_1051 (.ZN (n_987), .A (n_5665));
AOI21_X1 i_1050 (.ZN (n_986), .A (n_5669), .B1 (n_5678), .B2 (n_5675));
OAI21_X2 i_1049 (.ZN (n_985), .A (n_5660), .B1 (n_987), .B2 (n_986));
NAND2_X1 i_1048 (.ZN (n_984), .A1 (n_7476), .A2 (n_7475));
NAND2_X1 i_1047 (.ZN (n_983), .A1 (n_984), .A2 (n_7470));
NAND3_X1 i_1046 (.ZN (n_982), .A1 (n_5668), .A2 (n_983), .A3 (n_5688));
OAI21_X2 i_1045 (.ZN (n_981), .A (n_982), .B1 (n_988), .B2 (n_985));
AOI21_X2 i_1044 (.ZN (n_980), .A (n_981), .B1 (n_989), .B2 (CLOCK_opt_ipo_n351));
NAND3_X1 i_1043 (.ZN (n_979), .A1 (n_6936), .A2 (n_6964), .A3 (n_6943));
NAND2_X1 i_1042 (.ZN (n_978), .A1 (n_6939), .A2 (n_6942));
NAND2_X1 i_1041 (.ZN (n_977), .A1 (n_978), .A2 (n_6938));
NAND3_X1 i_1040 (.ZN (n_976), .A1 (n_7733), .A2 (n_7467), .A3 (n_7737));
NAND2_X1 i_1039 (.ZN (n_975), .A1 (n_977), .A2 (n_976));
INV_X1 i_1038 (.ZN (n_974), .A (n_975));
NAND2_X1 i_1037 (.ZN (n_973), .A1 (n_6941), .A2 (n_6952));
AOI22_X1 i_1036 (.ZN (n_972), .A1 (n_6963), .A2 (n_6961), .B1 (n_973), .B2 (n_6954));
AOI22_X1 i_1035 (.ZN (n_971), .A1 (n_7000), .A2 (n_6997), .B1 (n_6965), .B2 (n_6975));
AOI21_X1 i_1034 (.ZN (n_970), .A (n_971), .B1 (n_6964), .B2 (n_972));
OAI21_X1 i_1033 (.ZN (n_969), .A (n_970), .B1 (n_974), .B2 (n_979));
INV_X1 i_1032 (.ZN (n_968), .A (n_969));
OAI21_X1 i_1031 (.ZN (n_967), .A (n_968), .B1 (n_980), .B2 (n_6935));
NAND3_X1 i_1030 (.ZN (n_966), .A1 (n_5112), .A2 (n_5139), .A3 (n_5121));
INV_X1 i_1029 (.ZN (n_965), .A (n_5116));
NAND2_X1 i_1028 (.ZN (n_964), .A1 (n_965), .A2 (n_5114));
NAND2_X1 i_1027 (.ZN (n_963), .A1 (n_5655), .A2 (n_7200));
NAND2_X1 i_1026 (.ZN (n_962), .A1 (n_5506), .A2 (n_5509));
NAND2_X1 i_1025 (.ZN (n_961), .A1 (n_962), .A2 (n_963));
AND2_X1 i_1024 (.ZN (n_960), .A1 (n_964), .A2 (n_961));
NAND2_X1 i_1023 (.ZN (n_959), .A1 (n_5135), .A2 (n_5138));
NAND2_X1 i_1022 (.ZN (n_958), .A1 (n_5122), .A2 (n_5130));
NAND3_X1 i_1021 (.ZN (n_957), .A1 (n_5139), .A2 (n_959), .A3 (n_958));
NAND2_X1 i_1020 (.ZN (n_956), .A1 (n_5168), .A2 (n_5172));
INV_X1 i_1019 (.ZN (n_955), .A (n_5140));
OAI21_X2 i_1018 (.ZN (n_954), .A (n_956), .B1 (n_5137), .B2 (n_955));
OAI211_X2 i_1017 (.ZN (n_953), .A (n_957), .B (n_954), .C1 (n_960), .C2 (n_966));
AOI21_X2 i_1016 (.ZN (n_952), .A (n_953), .B1 (n_967), .B2 (CLOCK_opt_ipo_n528));
NAND3_X4 i_1015 (.ZN (n_951), .A1 (n_952), .A2 (n_995), .A3 (n_3980));
NAND2_X1 i_1014 (.ZN (n_950), .A1 (n_5344), .A2 (n_5358));
INV_X1 i_1013 (.ZN (n_949), .A (n_5253));
OAI21_X1 i_1012 (.ZN (n_948), .A (n_5255), .B1 (n_5259), .B2 (n_949));
INV_X1 i_1011 (.ZN (n_947), .A (n_948));
NAND3_X1 i_1010 (.ZN (n_946), .A1 (n_950), .A2 (n_5345), .A3 (n_947));
NAND2_X1 i_1009 (.ZN (n_945), .A1 (n_950), .A2 (n_5345));
NAND2_X1 i_1008 (.ZN (n_944), .A1 (n_945), .A2 (n_948));
NAND2_X1 i_1007 (.ZN (n_943), .A1 (n_944), .A2 (n_946));
NAND2_X1 i_1006 (.ZN (n_942), .A1 (n_5323), .A2 (n_5333));
NAND2_X1 i_1005 (.ZN (n_941), .A1 (n_5324), .A2 (n_942));
INV_X1 i_1004 (.ZN (n_940), .A (n_941));
XNOR2_X1 i_1003 (.ZN (n_939), .A (n_943), .B (n_940));
NAND2_X1 i_1002 (.ZN (n_938), .A1 (n_5248), .A2 (n_5265));
NAND2_X1 i_1001 (.ZN (n_937), .A1 (n_938), .A2 (n_5249));
OR2_X1 i_1000 (.ZN (n_936), .A1 (n_939), .A2 (n_937));
NAND2_X1 i_999 (.ZN (n_935), .A1 (n_939), .A2 (n_937));
NAND2_X1 i_998 (.ZN (n_934), .A1 (n_936), .A2 (n_935));
INV_X1 i_997 (.ZN (n_933), .A (n_5350));
INV_X1 i_996 (.ZN (n_932), .A (n_5348));
OAI21_X1 i_995 (.ZN (n_931), .A (n_5349), .B1 (n_933), .B2 (n_932));
INV_X1 i_994 (.ZN (n_930), .A (n_5261));
OAI21_X1 i_993 (.ZN (n_929), .A (n_5262), .B1 (n_5263), .B2 (n_930));
OAI21_X1 i_992 (.ZN (n_928), .A (n_929), .B1 (n_8958), .B2 (n_7912));
INV_X1 i_991 (.ZN (n_927), .A (n_929));
NAND3_X1 i_990 (.ZN (n_926), .A1 (n_927), .A2 (B_imm[22]), .A3 (A_imm[27]));
NAND2_X1 i_989 (.ZN (n_925), .A1 (n_926), .A2 (n_928));
XNOR2_X1 i_988 (.ZN (n_924), .A (n_925), .B (n_931));
NAND2_X1 i_987 (.ZN (n_923), .A1 (A_imm[28]), .A2 (B_imm[21]));
OAI22_X1 i_986 (.ZN (n_922), .A1 (n_9006), .A2 (n_8893), .B1 (CLOCK_opt_ipo_n433), .B2 (n_8906));
NAND4_X1 i_985 (.ZN (n_921), .A1 (B_imm[29]), .A2 (B_imm[27]), .A3 (A_imm[22]), .A4 (A_imm[20]));
NAND2_X1 i_984 (.ZN (n_920), .A1 (n_922), .A2 (n_921));
XNOR2_X1 i_983 (.ZN (n_919), .A (n_920), .B (n_923));
NAND2_X1 i_982 (.ZN (n_918), .A1 (n_924), .A2 (n_919));
OR2_X1 i_981 (.ZN (n_917), .A1 (n_924), .A2 (n_919));
NAND2_X1 i_980 (.ZN (n_916), .A1 (n_917), .A2 (n_918));
INV_X1 i_979 (.ZN (n_915), .A (n_5327));
OAI21_X1 i_978 (.ZN (n_914), .A (n_5328), .B1 (n_5329), .B2 (n_915));
INV_X1 i_977 (.ZN (n_913), .A (n_914));
OAI22_X1 i_976 (.ZN (n_912), .A1 (n_9038), .A2 (n_8956), .B1 (n_9004), .B2 (n_8892));
NAND4_X1 i_975 (.ZN (n_911), .A1 (B_imm[31]), .A2 (B_imm[30]), .A3 (A_imm[19]), .A4 (A_imm[18]));
NAND2_X1 i_974 (.ZN (n_910), .A1 (n_912), .A2 (n_911));
XNOR2_X1 i_973 (.ZN (n_909), .A (n_910), .B (n_913));
XNOR2_X1 i_972 (.ZN (n_908), .A (n_916), .B (n_909));
XOR2_X1 i_971 (.Z (n_907), .A (n_908), .B (n_934));
NAND2_X1 i_970 (.ZN (n_906), .A1 (n_5368), .A2 (n_5271));
AND2_X1 i_969 (.ZN (n_905), .A1 (n_906), .A2 (n_5273));
NAND2_X1 i_968 (.ZN (n_904), .A1 (n_907), .A2 (n_905));
OR2_X1 i_967 (.ZN (n_903), .A1 (n_907), .A2 (n_905));
NAND2_X1 i_966 (.ZN (n_902), .A1 (n_5225), .A2 (n_5223));
NAND2_X1 i_965 (.ZN (n_901), .A1 (n_902), .A2 (n_5226));
INV_X1 i_964 (.ZN (n_900), .A (n_5243));
INV_X1 i_963 (.ZN (n_899), .A (n_5241));
OAI21_X1 i_962 (.ZN (n_898), .A (n_5242), .B1 (n_900), .B2 (n_899));
OAI21_X1 i_961 (.ZN (n_897), .A (n_898), .B1 (n_8860), .B2 (n_8994));
OR3_X1 i_960 (.ZN (n_896), .A1 (n_898), .A2 (n_8860), .A3 (n_8994));
NAND2_X1 i_959 (.ZN (n_895), .A1 (n_896), .A2 (n_897));
NAND2_X1 i_958 (.ZN (n_894), .A1 (B_imm[23]), .A2 (A_imm[26]));
OAI22_X1 i_957 (.ZN (n_893), .A1 (n_8423), .A2 (n_9037), .B1 (n_8948), .B2 (n_8794));
NAND4_X1 i_956 (.ZN (n_892), .A1 (B_imm[24]), .A2 (opt_ipoPP_0), .A3 (B_imm[18]), .A4 (A_imm[25]));
NAND2_X1 i_955 (.ZN (n_891), .A1 (n_893), .A2 (n_892));
XNOR2_X1 i_954 (.ZN (n_890), .A (n_891), .B (n_894));
XNOR2_X1 i_953 (.ZN (n_889), .A (n_895), .B (n_890));
INV_X1 i_952 (.ZN (n_888), .A (n_889));
NAND2_X1 i_951 (.ZN (n_887), .A1 (n_888), .A2 (n_901));
NAND3_X1 i_950 (.ZN (n_886), .A1 (n_889), .A2 (n_902), .A3 (n_5226));
NAND2_X1 i_949 (.ZN (n_885), .A1 (n_886), .A2 (n_887));
NAND2_X1 i_948 (.ZN (n_884), .A1 (A_imm[30]), .A2 (B_imm[19]));
INV_X1 i_947 (.ZN (n_883), .A (n_5229));
OAI21_X1 i_946 (.ZN (n_882), .A (n_5231), .B1 (n_883), .B2 (n_5235));
NAND2_X1 i_945 (.ZN (n_881), .A1 (B_imm[26]), .A2 (A_imm[23]));
OAI22_X1 i_944 (.ZN (n_880), .A1 (n_9021), .A2 (n_8859), .B1 (n_8974), .B2 (n_8767));
NAND4_X1 i_943 (.ZN (n_879), .A1 (B_imm[28]), .A2 (B_imm[25]), .A3 (A_imm[24]), .A4 (A_imm[21]));
NAND2_X1 i_942 (.ZN (n_878), .A1 (n_880), .A2 (n_879));
XNOR2_X1 i_941 (.ZN (n_877), .A (n_878), .B (n_881));
OR2_X1 i_940 (.ZN (n_876), .A1 (n_882), .A2 (n_877));
NAND2_X1 i_939 (.ZN (n_875), .A1 (n_882), .A2 (n_877));
NAND2_X1 i_938 (.ZN (n_874), .A1 (n_876), .A2 (n_875));
XNOR2_X1 i_937 (.ZN (n_873), .A (n_874), .B (n_884));
XNOR2_X1 i_936 (.ZN (n_872), .A (n_885), .B (n_873));
INV_X1 i_935 (.ZN (n_871), .A (n_5335));
OAI21_X1 i_934 (.ZN (n_870), .A (n_5338), .B1 (n_871), .B2 (n_5321));
INV_X1 i_933 (.ZN (n_869), .A (n_870));
NAND2_X1 i_932 (.ZN (n_868), .A1 (n_872), .A2 (n_869));
INV_X1 i_931 (.ZN (n_867), .A (n_872));
NAND2_X1 i_930 (.ZN (n_866), .A1 (n_867), .A2 (n_870));
NAND2_X1 i_929 (.ZN (n_865), .A1 (n_866), .A2 (n_868));
NAND2_X1 i_928 (.ZN (n_864), .A1 (n_5246), .A2 (n_5216));
AND2_X1 i_927 (.ZN (n_863), .A1 (n_864), .A2 (n_5217));
XNOR2_X1 i_926 (.ZN (n_862), .A (n_865), .B (n_863));
INV_X1 i_925 (.ZN (n_861), .A (n_862));
NAND3_X1 i_924 (.ZN (n_860), .A1 (n_903), .A2 (n_904), .A3 (n_861));
NAND2_X1 i_923 (.ZN (n_859), .A1 (n_903), .A2 (n_904));
NAND2_X1 i_922 (.ZN (n_858), .A1 (n_859), .A2 (n_862));
NAND2_X1 i_921 (.ZN (n_857), .A1 (n_858), .A2 (n_860));
NAND2_X1 i_920 (.ZN (n_856), .A1 (n_5171), .A2 (n_5173));
NAND3_X1 i_919 (.ZN (n_855), .A1 (n_857), .A2 (n_5175), .A3 (n_856));
NAND2_X1 i_918 (.ZN (n_854), .A1 (n_936), .A2 (n_908));
NAND2_X1 i_917 (.ZN (n_853), .A1 (n_854), .A2 (n_935));
INV_X1 i_916 (.ZN (n_852), .A (n_853));
NAND2_X1 i_915 (.ZN (n_851), .A1 (n_918), .A2 (n_909));
NAND2_X1 i_914 (.ZN (n_850), .A1 (n_917), .A2 (n_851));
INV_X1 i_913 (.ZN (n_849), .A (n_875));
OAI21_X1 i_912 (.ZN (n_848), .A (n_876), .B1 (n_884), .B2 (n_849));
NAND2_X1 i_911 (.ZN (n_847), .A1 (n_850), .A2 (n_848));
OR2_X1 i_910 (.ZN (n_846), .A1 (n_850), .A2 (n_848));
NAND2_X1 i_909 (.ZN (n_845), .A1 (n_846), .A2 (n_847));
NAND2_X1 i_908 (.ZN (n_844), .A1 (n_926), .A2 (n_931));
NAND2_X1 i_907 (.ZN (n_843), .A1 (n_844), .A2 (n_928));
INV_X1 i_906 (.ZN (n_842), .A (n_843));
NAND2_X1 i_905 (.ZN (n_841), .A1 (B_imm[28]), .A2 (A_imm[22]));
INV_X1 i_904 (.ZN (n_840), .A (n_841));
OAI22_X1 i_903 (.ZN (n_839), .A1 (n_8974), .A2 (n_8794), .B1 (n_8948), .B2 (n_8972));
NAND4_X1 i_902 (.ZN (n_838), .A1 (B_imm[25]), .A2 (B_imm[24]), .A3 (A_imm[26]), .A4 (A_imm[25]));
NAND2_X1 i_901 (.ZN (n_837), .A1 (n_839), .A2 (n_838));
XNOR2_X1 i_900 (.ZN (n_836), .A (n_837), .B (n_840));
NAND2_X1 i_899 (.ZN (n_835), .A1 (n_842), .A2 (n_836));
INV_X1 i_898 (.ZN (n_834), .A (n_835));
NOR2_X1 i_897 (.ZN (n_833), .A1 (n_842), .A2 (n_836));
NOR2_X1 i_896 (.ZN (n_832), .A1 (n_834), .A2 (n_833));
NAND2_X1 i_895 (.ZN (n_831), .A1 (B_imm[27]), .A2 (A_imm[23]));
OAI22_X1 i_894 (.ZN (n_830), .A1 (n_8525), .A2 (n_9037), .B1 (n_8993), .B2 (n_8767));
NAND4_X1 i_893 (.ZN (n_829), .A1 (B_imm[19]), .A2 (B_imm[26]), .A3 (A_imm[31]), .A4 (A_imm[24]));
NAND2_X1 i_892 (.ZN (n_828), .A1 (n_830), .A2 (n_829));
XNOR2_X1 i_891 (.ZN (n_827), .A (n_828), .B (n_831));
XNOR2_X1 i_890 (.ZN (n_826), .A (n_832), .B (n_827));
XNOR2_X1 i_889 (.ZN (n_825), .A (n_845), .B (n_826));
INV_X1 i_888 (.ZN (n_824), .A (n_873));
NAND2_X1 i_887 (.ZN (n_823), .A1 (n_886), .A2 (n_824));
NAND2_X1 i_886 (.ZN (n_822), .A1 (n_823), .A2 (n_887));
NAND2_X1 i_885 (.ZN (n_821), .A1 (n_825), .A2 (n_822));
INV_X1 i_884 (.ZN (n_820), .A (n_825));
NAND3_X1 i_883 (.ZN (n_819), .A1 (n_820), .A2 (n_887), .A3 (n_823));
NAND2_X1 i_882 (.ZN (n_818), .A1 (n_819), .A2 (n_821));
XNOR2_X1 i_881 (.ZN (n_817), .A (n_818), .B (n_852));
NAND2_X1 i_880 (.ZN (n_816), .A1 (n_866), .A2 (n_863));
NAND2_X1 i_879 (.ZN (n_815), .A1 (n_816), .A2 (n_868));
INV_X1 i_878 (.ZN (n_814), .A (n_815));
INV_X1 i_877 (.ZN (n_813), .A (n_923));
INV_X1 i_876 (.ZN (n_812), .A (n_921));
OAI21_X1 i_875 (.ZN (n_811), .A (n_922), .B1 (n_813), .B2 (n_812));
AOI22_X1 i_874 (.ZN (n_810), .A1 (A_imm[29]), .A2 (B_imm[21]), .B1 (B_imm[31]), .B2 (A_imm[19]));
INV_X1 i_873 (.ZN (n_809), .A (n_810));
NAND4_X1 i_872 (.ZN (n_808), .A1 (A_imm[29]), .A2 (B_imm[31]), .A3 (B_imm[21]), .A4 (A_imm[19]));
NAND2_X1 i_871 (.ZN (n_807), .A1 (n_809), .A2 (n_808));
XOR2_X1 i_870 (.Z (n_806), .A (n_811), .B (n_807));
INV_X1 i_869 (.ZN (n_805), .A (n_897));
OAI21_X1 i_868 (.ZN (n_804), .A (n_896), .B1 (n_805), .B2 (n_890));
INV_X1 i_867 (.ZN (n_803), .A (n_804));
INV_X1 i_866 (.ZN (n_802), .A (n_881));
INV_X1 i_865 (.ZN (n_801), .A (n_879));
OAI21_X1 i_864 (.ZN (n_800), .A (n_880), .B1 (n_802), .B2 (n_801));
OAI22_X1 i_863 (.ZN (n_799), .A1 (n_9004), .A2 (n_8893), .B1 (n_7912), .B2 (n_8821));
NAND4_X1 i_862 (.ZN (n_798), .A1 (B_imm[30]), .A2 (A_imm[27]), .A3 (B_imm[23]), .A4 (A_imm[20]));
NAND2_X1 i_861 (.ZN (n_797), .A1 (n_799), .A2 (n_798));
XNOR2_X1 i_860 (.ZN (n_796), .A (n_797), .B (n_800));
OR2_X1 i_859 (.ZN (n_795), .A1 (n_803), .A2 (n_796));
NAND2_X1 i_858 (.ZN (n_794), .A1 (n_803), .A2 (n_796));
NAND2_X1 i_857 (.ZN (n_793), .A1 (n_795), .A2 (n_794));
XNOR2_X1 i_856 (.ZN (n_792), .A (n_793), .B (n_806));
NAND2_X1 i_855 (.ZN (n_791), .A1 (n_892), .A2 (n_894));
NAND2_X1 i_854 (.ZN (n_790), .A1 (n_893), .A2 (n_791));
INV_X1 i_853 (.ZN (n_789), .A (n_790));
OAI22_X1 i_852 (.ZN (n_788), .A1 (n_9020), .A2 (n_8958), .B1 (n_9006), .B2 (n_8859));
NAND4_X1 i_851 (.ZN (n_787), .A1 (A_imm[28]), .A2 (B_imm[29]), .A3 (B_imm[22]), .A4 (A_imm[21]));
NAND2_X1 i_850 (.ZN (n_786), .A1 (n_788), .A2 (n_787));
XNOR2_X1 i_849 (.ZN (n_785), .A (n_786), .B (n_789));
INV_X1 i_848 (.ZN (n_784), .A (n_911));
OAI21_X1 i_847 (.ZN (n_783), .A (n_912), .B1 (n_913), .B2 (n_784));
OR3_X1 i_846 (.ZN (n_782), .A1 (n_783), .A2 (n_8860), .A3 (n_9005));
OAI21_X1 i_845 (.ZN (n_781), .A (n_783), .B1 (n_8860), .B2 (n_9005));
NAND2_X1 i_844 (.ZN (n_780), .A1 (n_782), .A2 (n_781));
XNOR2_X1 i_843 (.ZN (n_779), .A (n_780), .B (n_785));
INV_X1 i_842 (.ZN (n_778), .A (n_946));
OAI21_X1 i_841 (.ZN (n_777), .A (n_944), .B1 (n_778), .B2 (n_940));
INV_X1 i_840 (.ZN (n_776), .A (n_777));
NAND2_X1 i_839 (.ZN (n_775), .A1 (n_779), .A2 (n_776));
OR2_X1 i_838 (.ZN (n_774), .A1 (n_779), .A2 (n_776));
NAND2_X1 i_837 (.ZN (n_773), .A1 (n_774), .A2 (n_775));
XNOR2_X1 i_836 (.ZN (n_772), .A (n_792), .B (n_773));
NAND2_X1 i_835 (.ZN (n_771), .A1 (n_814), .A2 (n_772));
NOR2_X1 i_834 (.ZN (n_770), .A1 (n_814), .A2 (n_772));
INV_X1 i_833 (.ZN (n_769), .A (n_770));
NAND3_X1 i_832 (.ZN (n_768), .A1 (n_817), .A2 (n_769), .A3 (n_771));
INV_X1 i_831 (.ZN (n_767), .A (n_817));
INV_X1 i_830 (.ZN (n_766), .A (n_771));
OAI21_X1 i_829 (.ZN (n_765), .A (n_767), .B1 (n_766), .B2 (n_770));
NAND2_X1 i_828 (.ZN (n_764), .A1 (n_861), .A2 (n_904));
NAND2_X1 i_827 (.ZN (n_763), .A1 (n_764), .A2 (n_903));
INV_X1 i_826 (.ZN (n_762), .A (n_763));
NAND3_X1 i_825 (.ZN (n_761), .A1 (n_762), .A2 (n_768), .A3 (n_765));
INV_X1 i_824 (.ZN (n_760), .A (n_800));
INV_X1 i_823 (.ZN (n_759), .A (n_798));
OAI21_X1 i_822 (.ZN (n_758), .A (n_799), .B1 (n_760), .B2 (n_759));
NAND2_X1 i_821 (.ZN (n_757), .A1 (B_imm[28]), .A2 (A_imm[23]));
OAI22_X1 i_820 (.ZN (n_756), .A1 (n_8860), .A2 (n_9037), .B1 (n_8974), .B2 (n_8972));
NAND4_X1 i_819 (.ZN (n_755), .A1 (B_imm[20]), .A2 (B_imm[25]), .A3 (opt_ipoPP_0), .A4 (A_imm[26]));
NAND2_X1 i_818 (.ZN (n_754), .A1 (n_756), .A2 (n_755));
XNOR2_X1 i_817 (.ZN (n_753), .A (n_754), .B (n_757));
INV_X1 i_816 (.ZN (n_752), .A (n_753));
NAND3_X1 i_815 (.ZN (n_751), .A1 (n_752), .A2 (B_imm[21]), .A3 (A_imm[30]));
OAI21_X1 i_814 (.ZN (n_750), .A (n_753), .B1 (n_8957), .B2 (n_9005));
NAND2_X1 i_813 (.ZN (n_749), .A1 (n_751), .A2 (n_750));
XNOR2_X1 i_812 (.ZN (n_748), .A (n_749), .B (n_758));
NAND2_X1 i_811 (.ZN (n_747), .A1 (n_794), .A2 (n_806));
NAND2_X1 i_810 (.ZN (n_746), .A1 (n_795), .A2 (n_747));
INV_X1 i_809 (.ZN (n_745), .A (n_746));
NAND2_X1 i_808 (.ZN (n_744), .A1 (n_745), .A2 (n_748));
OR2_X1 i_807 (.ZN (n_743), .A1 (n_745), .A2 (n_748));
NAND2_X1 i_806 (.ZN (n_742), .A1 (n_743), .A2 (n_744));
AOI21_X1 i_805 (.ZN (n_741), .A (n_810), .B1 (n_811), .B2 (n_808));
INV_X1 i_804 (.ZN (n_740), .A (n_838));
OAI21_X1 i_803 (.ZN (n_739), .A (n_839), .B1 (n_740), .B2 (n_840));
AOI22_X1 i_802 (.ZN (n_738), .A1 (A_imm[27]), .A2 (B_imm[24]), .B1 (A_imm[28]), .B2 (B_imm[23]));
INV_X1 i_801 (.ZN (n_737), .A (n_738));
NAND4_X1 i_800 (.ZN (n_736), .A1 (A_imm[27]), .A2 (B_imm[24]), .A3 (B_imm[23]), .A4 (A_imm[28]));
NAND2_X1 i_799 (.ZN (n_735), .A1 (n_737), .A2 (n_736));
XOR2_X1 i_798 (.Z (n_734), .A (n_739), .B (n_735));
OR2_X1 i_797 (.ZN (n_733), .A1 (n_734), .A2 (n_741));
NAND2_X1 i_796 (.ZN (n_732), .A1 (n_734), .A2 (n_741));
NAND2_X1 i_795 (.ZN (n_731), .A1 (n_733), .A2 (n_732));
OAI22_X1 i_794 (.ZN (n_730), .A1 (n_9038), .A2 (n_8893), .B1 (n_9004), .B2 (n_8859));
NAND4_X1 i_793 (.ZN (n_729), .A1 (B_imm[31]), .A2 (B_imm[30]), .A3 (A_imm[21]), .A4 (A_imm[20]));
NAND2_X1 i_792 (.ZN (n_728), .A1 (n_730), .A2 (n_729));
NAND2_X1 i_791 (.ZN (n_727), .A1 (n_829), .A2 (n_831));
NAND2_X1 i_790 (.ZN (n_726), .A1 (n_727), .A2 (n_830));
INV_X1 i_789 (.ZN (n_725), .A (n_726));
XNOR2_X1 i_788 (.ZN (n_724), .A (n_728), .B (n_725));
XOR2_X1 i_787 (.Z (n_723), .A (n_724), .B (n_731));
XNOR2_X1 i_786 (.ZN (n_722), .A (n_742), .B (n_723));
NAND2_X1 i_785 (.ZN (n_721), .A1 (n_819), .A2 (n_853));
NAND3_X1 i_784 (.ZN (n_720), .A1 (n_722), .A2 (n_821), .A3 (n_721));
INV_X1 i_783 (.ZN (n_719), .A (n_722));
NAND2_X1 i_782 (.ZN (n_718), .A1 (n_721), .A2 (n_821));
NAND2_X1 i_781 (.ZN (n_717), .A1 (n_718), .A2 (n_719));
NAND2_X1 i_780 (.ZN (n_716), .A1 (n_781), .A2 (n_785));
NAND2_X1 i_779 (.ZN (n_715), .A1 (n_782), .A2 (n_716));
OAI21_X1 i_778 (.ZN (n_714), .A (n_835), .B1 (n_833), .B2 (n_827));
NAND2_X1 i_777 (.ZN (n_713), .A1 (n_715), .A2 (n_714));
OR2_X1 i_776 (.ZN (n_712), .A1 (n_714), .A2 (n_715));
NAND2_X1 i_775 (.ZN (n_711), .A1 (n_712), .A2 (n_713));
INV_X1 i_774 (.ZN (n_710), .A (n_787));
OAI21_X1 i_773 (.ZN (n_709), .A (n_788), .B1 (n_789), .B2 (n_710));
INV_X1 i_772 (.ZN (n_708), .A (n_709));
NAND3_X1 i_771 (.ZN (n_707), .A1 (n_708), .A2 (B_imm[22]), .A3 (A_imm[29]));
INV_X1 i_770 (.ZN (n_706), .A (n_707));
AOI21_X1 i_769 (.ZN (n_705), .A (n_708), .B1 (B_imm[22]), .B2 (A_imm[29]));
OR2_X1 i_768 (.ZN (n_704), .A1 (n_706), .A2 (n_705));
INV_X1 i_767 (.ZN (n_703), .A (n_704));
NAND2_X1 i_766 (.ZN (n_702), .A1 (B_imm[29]), .A2 (A_imm[22]));
OAI22_X1 i_765 (.ZN (n_701), .A1 (CLOCK_opt_ipo_n433), .A2 (n_8767), .B1 (n_8993), .B2 (n_8794));
NAND4_X1 i_764 (.ZN (n_700), .A1 (B_imm[27]), .A2 (B_imm[26]), .A3 (A_imm[25]), .A4 (A_imm[24]));
NAND2_X1 i_763 (.ZN (n_699), .A1 (n_701), .A2 (n_700));
XNOR2_X1 i_762 (.ZN (n_698), .A (n_699), .B (n_702));
XNOR2_X1 i_761 (.ZN (n_697), .A (n_703), .B (n_698));
INV_X1 i_760 (.ZN (n_696), .A (n_697));
XNOR2_X1 i_759 (.ZN (n_695), .A (n_711), .B (n_696));
INV_X1 i_758 (.ZN (n_694), .A (n_847));
AOI21_X1 i_757 (.ZN (n_693), .A (n_694), .B1 (n_846), .B2 (n_826));
NAND2_X1 i_756 (.ZN (n_692), .A1 (n_693), .A2 (n_695));
OR2_X1 i_755 (.ZN (n_691), .A1 (n_695), .A2 (n_693));
NAND2_X1 i_754 (.ZN (n_690), .A1 (n_691), .A2 (n_692));
INV_X1 i_753 (.ZN (n_689), .A (n_690));
INV_X1 i_752 (.ZN (n_688), .A (n_775));
AOI21_X1 i_751 (.ZN (n_687), .A (n_688), .B1 (n_792), .B2 (n_774));
XNOR2_X1 i_750 (.ZN (n_686), .A (n_689), .B (n_687));
NAND3_X1 i_749 (.ZN (n_685), .A1 (n_686), .A2 (n_717), .A3 (n_720));
NAND2_X1 i_748 (.ZN (n_684), .A1 (n_717), .A2 (n_720));
INV_X1 i_747 (.ZN (n_683), .A (n_686));
NAND2_X1 i_746 (.ZN (n_682), .A1 (n_684), .A2 (n_683));
NAND2_X1 i_745 (.ZN (n_681), .A1 (n_682), .A2 (n_685));
OAI21_X1 i_744 (.ZN (n_680), .A (n_771), .B1 (n_817), .B2 (n_770));
INV_X1 i_743 (.ZN (n_679), .A (n_680));
NAND2_X1 i_742 (.ZN (n_678), .A1 (n_679), .A2 (n_681));
NAND2_X1 i_741 (.ZN (n_677), .A1 (A_imm[30]), .A2 (B_imm[22]));
AOI21_X1 i_740 (.ZN (n_676), .A (n_738), .B1 (n_739), .B2 (n_736));
INV_X1 i_739 (.ZN (n_675), .A (n_676));
NAND2_X1 i_738 (.ZN (n_674), .A1 (B_imm[26]), .A2 (A_imm[26]));
OAI22_X1 i_737 (.ZN (n_673), .A1 (n_9021), .A2 (n_8767), .B1 (n_8957), .B2 (n_9037));
NAND4_X1 i_736 (.ZN (n_672), .A1 (B_imm[28]), .A2 (B_imm[21]), .A3 (opt_ipoPP_0), .A4 (A_imm[24]));
NAND2_X1 i_735 (.ZN (n_671), .A1 (n_673), .A2 (n_672));
XNOR2_X1 i_734 (.ZN (n_670), .A (n_671), .B (n_674));
OR2_X1 i_733 (.ZN (n_669), .A1 (n_670), .A2 (n_675));
NAND2_X1 i_732 (.ZN (n_668), .A1 (n_670), .A2 (n_675));
NAND2_X1 i_731 (.ZN (n_667), .A1 (n_669), .A2 (n_668));
XOR2_X1 i_730 (.Z (n_666), .A (n_677), .B (n_667));
NAND2_X1 i_729 (.ZN (n_665), .A1 (n_733), .A2 (n_724));
NAND2_X1 i_728 (.ZN (n_664), .A1 (n_665), .A2 (n_732));
NAND2_X1 i_727 (.ZN (n_663), .A1 (n_666), .A2 (n_664));
OR2_X1 i_726 (.ZN (n_662), .A1 (n_666), .A2 (n_664));
NAND2_X1 i_725 (.ZN (n_661), .A1 (n_662), .A2 (n_663));
INV_X1 i_724 (.ZN (n_660), .A (n_729));
OAI21_X1 i_723 (.ZN (n_659), .A (n_730), .B1 (n_725), .B2 (n_660));
NAND2_X1 i_722 (.ZN (n_658), .A1 (A_imm[28]), .A2 (B_imm[24]));
OAI22_X1 i_721 (.ZN (n_657), .A1 (n_9006), .A2 (n_8907), .B1 (CLOCK_opt_ipo_n433), .B2 (n_8794));
NAND4_X1 i_720 (.ZN (n_656), .A1 (B_imm[29]), .A2 (B_imm[27]), .A3 (A_imm[25]), .A4 (A_imm[23]));
NAND2_X1 i_719 (.ZN (n_655), .A1 (n_657), .A2 (n_656));
XNOR2_X1 i_718 (.ZN (n_654), .A (n_655), .B (n_658));
OR2_X1 i_717 (.ZN (n_653), .A1 (n_654), .A2 (n_659));
NAND2_X1 i_716 (.ZN (n_652), .A1 (n_654), .A2 (n_659));
NAND2_X1 i_715 (.ZN (n_651), .A1 (n_653), .A2 (n_652));
OAI22_X1 i_714 (.ZN (n_650), .A1 (n_9004), .A2 (n_8906), .B1 (n_7912), .B2 (n_8974));
INV_X1 i_713 (.ZN (n_649), .A (n_650));
NAND4_X1 i_712 (.ZN (n_648), .A1 (B_imm[30]), .A2 (A_imm[27]), .A3 (B_imm[25]), .A4 (A_imm[22]));
NAND2_X1 i_711 (.ZN (n_647), .A1 (n_650), .A2 (n_648));
INV_X1 i_710 (.ZN (n_646), .A (n_647));
NAND2_X1 i_709 (.ZN (n_645), .A1 (n_755), .A2 (n_757));
NAND2_X1 i_708 (.ZN (n_644), .A1 (n_645), .A2 (n_756));
NAND2_X1 i_707 (.ZN (n_643), .A1 (n_648), .A2 (n_644));
OAI22_X1 i_706 (.ZN (n_642), .A1 (n_646), .A2 (n_644), .B1 (n_649), .B2 (n_643));
XNOR2_X1 i_705 (.ZN (n_641), .A (n_651), .B (n_642));
XOR2_X1 i_704 (.Z (n_640), .A (n_641), .B (n_661));
INV_X1 i_703 (.ZN (n_639), .A (n_692));
OAI21_X1 i_702 (.ZN (n_638), .A (n_691), .B1 (n_687), .B2 (n_639));
INV_X1 i_701 (.ZN (n_637), .A (n_638));
OR2_X1 i_700 (.ZN (n_636), .A1 (n_637), .A2 (n_640));
NAND2_X1 i_699 (.ZN (n_635), .A1 (n_640), .A2 (n_637));
NAND2_X1 i_698 (.ZN (n_634), .A1 (n_636), .A2 (n_635));
OAI21_X1 i_697 (.ZN (n_633), .A (n_707), .B1 (n_705), .B2 (n_698));
NAND2_X1 i_696 (.ZN (n_632), .A1 (n_751), .A2 (n_758));
NAND3_X1 i_695 (.ZN (n_631), .A1 (n_633), .A2 (n_632), .A3 (n_750));
INV_X1 i_694 (.ZN (n_630), .A (n_633));
NAND2_X1 i_693 (.ZN (n_629), .A1 (n_632), .A2 (n_750));
NAND2_X1 i_692 (.ZN (n_628), .A1 (n_629), .A2 (n_630));
NAND2_X1 i_691 (.ZN (n_627), .A1 (n_628), .A2 (n_631));
NAND2_X1 i_690 (.ZN (n_626), .A1 (A_imm[29]), .A2 (B_imm[23]));
NAND2_X1 i_689 (.ZN (n_625), .A1 (n_700), .A2 (n_702));
NAND2_X1 i_688 (.ZN (n_624), .A1 (n_625), .A2 (n_701));
INV_X1 i_687 (.ZN (n_623), .A (n_624));
NAND3_X1 i_686 (.ZN (n_622), .A1 (n_623), .A2 (B_imm[31]), .A3 (A_imm[21]));
AOI21_X1 i_685 (.ZN (n_621), .A (n_623), .B1 (B_imm[31]), .B2 (A_imm[21]));
INV_X1 i_684 (.ZN (n_620), .A (n_621));
NAND2_X1 i_683 (.ZN (n_619), .A1 (n_620), .A2 (n_622));
XOR2_X1 i_682 (.Z (n_618), .A (n_626), .B (n_619));
XOR2_X1 i_681 (.Z (n_617), .A (n_627), .B (n_618));
INV_X1 i_680 (.ZN (n_616), .A (n_712));
OAI21_X1 i_679 (.ZN (n_615), .A (n_713), .B1 (n_696), .B2 (n_616));
INV_X1 i_678 (.ZN (n_614), .A (n_615));
OR2_X1 i_677 (.ZN (n_613), .A1 (n_617), .A2 (n_614));
NAND2_X1 i_676 (.ZN (n_612), .A1 (n_617), .A2 (n_614));
NAND2_X1 i_675 (.ZN (n_611), .A1 (n_613), .A2 (n_612));
INV_X1 i_674 (.ZN (n_610), .A (n_744));
OAI21_X1 i_673 (.ZN (n_609), .A (n_743), .B1 (n_723), .B2 (n_610));
INV_X1 i_672 (.ZN (n_608), .A (n_609));
XNOR2_X1 i_671 (.ZN (n_607), .A (n_611), .B (n_608));
INV_X1 i_670 (.ZN (n_606), .A (n_607));
NAND2_X1 i_669 (.ZN (n_605), .A1 (n_634), .A2 (n_606));
NAND3_X1 i_668 (.ZN (n_604), .A1 (n_636), .A2 (n_635), .A3 (n_607));
NAND2_X1 i_667 (.ZN (n_603), .A1 (n_605), .A2 (n_604));
NAND2_X1 i_666 (.ZN (n_602), .A1 (n_686), .A2 (n_720));
NAND2_X1 i_665 (.ZN (n_601), .A1 (n_602), .A2 (n_717));
OR2_X1 i_664 (.ZN (n_600), .A1 (n_603), .A2 (n_601));
NAND4_X1 i_663 (.ZN (n_599), .A1 (n_855), .A2 (n_761), .A3 (n_678), .A4 (n_600));
INV_X1 i_662 (.ZN (n_598), .A (n_599));
NAND3_X1 i_661 (.ZN (n_597), .A1 (n_600), .A2 (n_761), .A3 (n_678));
INV_X1 i_660 (.ZN (n_596), .A (n_678));
NAND2_X1 i_659 (.ZN (n_595), .A1 (n_765), .A2 (n_768));
NAND2_X1 i_658 (.ZN (n_594), .A1 (n_595), .A2 (n_763));
NAND3_X1 i_657 (.ZN (n_593), .A1 (n_680), .A2 (n_685), .A3 (n_682));
OAI21_X1 i_656 (.ZN (n_592), .A (n_593), .B1 (n_594), .B2 (n_596));
NAND2_X1 i_655 (.ZN (n_591), .A1 (n_592), .A2 (n_600));
NAND2_X1 i_654 (.ZN (n_590), .A1 (n_856), .A2 (n_5175));
NAND3_X1 i_653 (.ZN (n_589), .A1 (n_858), .A2 (n_860), .A3 (n_590));
NAND2_X1 i_652 (.ZN (n_588), .A1 (n_603), .A2 (n_601));
OAI211_X1 i_651 (.ZN (n_587), .A (n_591), .B (n_588), .C1 (n_597), .C2 (n_589));
AOI21_X4 i_650 (.ZN (n_586), .A (n_587), .B1 (n_951), .B2 (n_598));
NAND2_X1 i_649 (.ZN (n_585), .A1 (n_656), .A2 (n_658));
NAND2_X1 i_648 (.ZN (n_584), .A1 (n_585), .A2 (n_657));
INV_X1 i_647 (.ZN (n_583), .A (n_584));
NAND3_X1 i_646 (.ZN (n_582), .A1 (n_583), .A2 (B_imm[24]), .A3 (A_imm[29]));
OAI21_X1 i_645 (.ZN (n_581), .A (n_584), .B1 (n_8948), .B2 (n_8994));
NAND2_X1 i_644 (.ZN (n_580), .A1 (n_582), .A2 (n_581));
NAND2_X1 i_643 (.ZN (n_579), .A1 (B_imm[27]), .A2 (A_imm[26]));
OAI22_X1 i_642 (.ZN (n_578), .A1 (n_9021), .A2 (n_8794), .B1 (n_8958), .B2 (n_9037));
NAND4_X1 i_641 (.ZN (n_577), .A1 (B_imm[28]), .A2 (B_imm[22]), .A3 (opt_ipoPP_0), .A4 (A_imm[25]));
NAND2_X1 i_640 (.ZN (n_576), .A1 (n_578), .A2 (n_577));
XOR2_X1 i_639 (.Z (n_575), .A (n_579), .B (n_576));
XNOR2_X1 i_638 (.ZN (n_574), .A (n_575), .B (n_580));
NAND2_X1 i_637 (.ZN (n_573), .A1 (n_652), .A2 (n_642));
NAND2_X1 i_636 (.ZN (n_572), .A1 (n_653), .A2 (n_573));
NAND2_X1 i_635 (.ZN (n_571), .A1 (n_574), .A2 (n_572));
OR2_X1 i_634 (.ZN (n_570), .A1 (n_574), .A2 (n_572));
NAND2_X1 i_633 (.ZN (n_569), .A1 (n_570), .A2 (n_571));
NAND4_X1 i_632 (.ZN (n_568), .A1 (n_643), .A2 (n_650), .A3 (A_imm[30]), .A4 (B_imm[23]));
NAND2_X1 i_631 (.ZN (n_567), .A1 (n_643), .A2 (n_650));
OAI21_X1 i_630 (.ZN (n_566), .A (n_567), .B1 (n_8821), .B2 (n_9005));
NAND2_X1 i_629 (.ZN (n_565), .A1 (n_566), .A2 (n_568));
AOI21_X1 i_628 (.ZN (n_564), .A (n_621), .B1 (n_626), .B2 (n_622));
XNOR2_X1 i_627 (.ZN (n_563), .A (n_565), .B (n_564));
XNOR2_X1 i_626 (.ZN (n_562), .A (n_569), .B (n_563));
INV_X1 i_625 (.ZN (n_561), .A (n_612));
OAI21_X1 i_624 (.ZN (n_560), .A (n_613), .B1 (n_561), .B2 (n_608));
OR2_X1 i_623 (.ZN (n_559), .A1 (n_560), .A2 (n_562));
NAND2_X1 i_622 (.ZN (n_558), .A1 (n_560), .A2 (n_562));
NAND2_X1 i_621 (.ZN (n_557), .A1 (n_559), .A2 (n_558));
NAND2_X1 i_620 (.ZN (n_556), .A1 (A_imm[27]), .A2 (B_imm[26]));
OAI22_X1 i_619 (.ZN (n_555), .A1 (n_9020), .A2 (n_8974), .B1 (n_9006), .B2 (n_8767));
NAND4_X1 i_618 (.ZN (n_554), .A1 (A_imm[28]), .A2 (B_imm[29]), .A3 (B_imm[25]), .A4 (A_imm[24]));
NAND2_X1 i_617 (.ZN (n_553), .A1 (n_555), .A2 (n_554));
XNOR2_X1 i_616 (.ZN (n_552), .A (n_553), .B (n_556));
NAND2_X1 i_615 (.ZN (n_551), .A1 (B_imm[31]), .A2 (A_imm[22]));
INV_X1 i_614 (.ZN (n_550), .A (n_551));
NAND2_X1 i_613 (.ZN (n_549), .A1 (n_672), .A2 (n_674));
NAND2_X1 i_612 (.ZN (n_548), .A1 (n_549), .A2 (n_673));
OAI21_X1 i_611 (.ZN (n_547), .A (n_548), .B1 (n_9004), .B2 (n_8907));
INV_X1 i_610 (.ZN (n_546), .A (n_548));
NAND3_X1 i_609 (.ZN (n_545), .A1 (n_546), .A2 (B_imm[30]), .A3 (A_imm[23]));
NAND2_X1 i_608 (.ZN (n_544), .A1 (n_545), .A2 (n_547));
XNOR2_X1 i_607 (.ZN (n_543), .A (n_544), .B (n_550));
INV_X1 i_606 (.ZN (n_542), .A (n_543));
OR2_X1 i_605 (.ZN (n_541), .A1 (n_542), .A2 (n_552));
NAND2_X1 i_604 (.ZN (n_540), .A1 (n_542), .A2 (n_552));
NAND2_X1 i_603 (.ZN (n_539), .A1 (n_541), .A2 (n_540));
INV_X1 i_602 (.ZN (n_538), .A (n_668));
OAI21_X1 i_601 (.ZN (n_537), .A (n_669), .B1 (n_677), .B2 (n_538));
XNOR2_X1 i_600 (.ZN (n_536), .A (n_539), .B (n_537));
NAND2_X1 i_599 (.ZN (n_535), .A1 (n_618), .A2 (n_628));
NAND2_X1 i_598 (.ZN (n_534), .A1 (n_535), .A2 (n_631));
NAND2_X1 i_597 (.ZN (n_533), .A1 (n_536), .A2 (n_534));
OR2_X1 i_596 (.ZN (n_532), .A1 (n_536), .A2 (n_534));
NAND2_X1 i_595 (.ZN (n_531), .A1 (n_532), .A2 (n_533));
NAND2_X1 i_594 (.ZN (n_530), .A1 (n_662), .A2 (n_641));
NAND2_X1 i_593 (.ZN (n_529), .A1 (n_530), .A2 (n_663));
XOR2_X1 i_592 (.Z (n_528), .A (n_529), .B (n_531));
INV_X1 i_591 (.ZN (n_527), .A (n_528));
XNOR2_X1 i_590 (.ZN (n_526), .A (n_527), .B (n_557));
INV_X1 i_589 (.ZN (n_525), .A (n_526));
NAND2_X1 i_588 (.ZN (n_524), .A1 (n_606), .A2 (n_635));
NAND2_X1 i_587 (.ZN (n_523), .A1 (n_636), .A2 (n_524));
INV_X1 i_586 (.ZN (n_522), .A (n_523));
NAND2_X1 i_585 (.ZN (n_521), .A1 (n_525), .A2 (n_522));
NAND2_X1 i_584 (.ZN (n_520), .A1 (A_imm[30]), .A2 (B_imm[26]));
INV_X1 i_583 (.ZN (n_519), .A (n_520));
OAI22_X1 i_582 (.ZN (n_518), .A1 (n_9004), .A2 (n_8794), .B1 (n_7912), .B2 (n_9021));
NAND2_X1 i_581 (.ZN (n_517), .A1 (B_imm[31]), .A2 (A_imm[24]));
INV_X1 i_580 (.ZN (n_516), .A (n_517));
NAND4_X1 i_579 (.ZN (n_515), .A1 (B_imm[30]), .A2 (A_imm[27]), .A3 (B_imm[28]), .A4 (A_imm[25]));
INV_X1 i_578 (.ZN (n_514), .A (n_515));
OAI21_X1 i_577 (.ZN (n_513), .A (n_518), .B1 (n_516), .B2 (n_514));
OAI22_X1 i_576 (.ZN (n_512), .A1 (n_9006), .A2 (n_8972), .B1 (n_8948), .B2 (n_9037));
NAND2_X1 i_575 (.ZN (n_511), .A1 (A_imm[28]), .A2 (B_imm[27]));
NAND4_X1 i_574 (.ZN (n_510), .A1 (B_imm[29]), .A2 (B_imm[24]), .A3 (opt_ipoPP_0), .A4 (A_imm[26]));
NAND2_X1 i_573 (.ZN (n_509), .A1 (n_510), .A2 (n_511));
NAND2_X1 i_572 (.ZN (n_508), .A1 (n_509), .A2 (n_512));
NAND2_X1 i_571 (.ZN (n_507), .A1 (n_513), .A2 (n_508));
INV_X1 i_570 (.ZN (n_506), .A (n_513));
INV_X1 i_569 (.ZN (n_505), .A (n_508));
NAND2_X1 i_568 (.ZN (n_504), .A1 (n_506), .A2 (n_505));
NAND2_X1 i_567 (.ZN (n_503), .A1 (n_504), .A2 (n_507));
XNOR2_X1 i_566 (.ZN (n_502), .A (n_503), .B (n_519));
NAND2_X1 i_565 (.ZN (n_501), .A1 (n_577), .A2 (n_579));
NAND2_X1 i_564 (.ZN (n_500), .A1 (n_501), .A2 (n_578));
OAI21_X1 i_563 (.ZN (n_499), .A (n_500), .B1 (n_9038), .B2 (n_8907));
NAND2_X1 i_562 (.ZN (n_498), .A1 (A_imm[29]), .A2 (B_imm[25]));
NAND4_X1 i_561 (.ZN (n_497), .A1 (n_501), .A2 (n_578), .A3 (B_imm[31]), .A4 (A_imm[23]));
NAND2_X1 i_560 (.ZN (n_496), .A1 (n_497), .A2 (n_498));
NAND2_X1 i_559 (.ZN (n_495), .A1 (n_496), .A2 (n_499));
INV_X1 i_558 (.ZN (n_494), .A (n_495));
NAND3_X1 i_557 (.ZN (n_493), .A1 (n_494), .A2 (B_imm[25]), .A3 (A_imm[30]));
AOI21_X1 i_556 (.ZN (n_492), .A (n_494), .B1 (B_imm[25]), .B2 (A_imm[30]));
NAND2_X1 i_555 (.ZN (n_491), .A1 (n_512), .A2 (n_510));
XOR2_X1 i_554 (.Z (n_490), .A (n_511), .B (n_491));
INV_X1 i_553 (.ZN (n_489), .A (n_490));
OAI21_X1 i_552 (.ZN (n_488), .A (n_493), .B1 (n_489), .B2 (n_492));
OR2_X1 i_551 (.ZN (n_487), .A1 (n_502), .A2 (n_488));
NAND2_X1 i_550 (.ZN (n_486), .A1 (n_502), .A2 (n_488));
NAND2_X1 i_549 (.ZN (n_485), .A1 (n_487), .A2 (n_486));
NAND2_X1 i_548 (.ZN (n_484), .A1 (n_518), .A2 (n_515));
XNOR2_X1 i_547 (.ZN (n_483), .A (n_484), .B (n_517));
NAND2_X1 i_546 (.ZN (n_482), .A1 (n_554), .A2 (n_556));
NAND2_X1 i_545 (.ZN (n_481), .A1 (n_482), .A2 (n_555));
NAND2_X1 i_544 (.ZN (n_480), .A1 (B_imm[29]), .A2 (A_imm[25]));
OAI22_X1 i_543 (.ZN (n_479), .A1 (n_9021), .A2 (n_8972), .B1 (n_8821), .B2 (n_9037));
NAND4_X1 i_542 (.ZN (n_478), .A1 (B_imm[28]), .A2 (B_imm[23]), .A3 (opt_ipoPP_0), .A4 (A_imm[26]));
NAND2_X1 i_541 (.ZN (n_477), .A1 (n_479), .A2 (n_478));
XNOR2_X1 i_540 (.ZN (n_476), .A (n_477), .B (n_480));
OR2_X1 i_539 (.ZN (n_475), .A1 (n_476), .A2 (n_481));
NAND2_X1 i_538 (.ZN (n_474), .A1 (A_imm[30]), .A2 (B_imm[24]));
NAND2_X1 i_537 (.ZN (n_473), .A1 (n_476), .A2 (n_481));
INV_X1 i_536 (.ZN (n_472), .A (n_473));
OAI21_X1 i_535 (.ZN (n_471), .A (n_475), .B1 (n_474), .B2 (n_472));
INV_X1 i_534 (.ZN (n_470), .A (n_471));
OR2_X1 i_533 (.ZN (n_469), .A1 (n_470), .A2 (n_483));
NAND2_X1 i_532 (.ZN (n_468), .A1 (n_470), .A2 (n_483));
OAI22_X1 i_531 (.ZN (n_467), .A1 (n_7912), .A2 (CLOCK_opt_ipo_n433), .B1 (n_9020), .B2 (n_8993));
NAND2_X1 i_530 (.ZN (n_466), .A1 (B_imm[30]), .A2 (A_imm[24]));
INV_X1 i_529 (.ZN (n_465), .A (n_466));
NAND4_X1 i_528 (.ZN (n_464), .A1 (A_imm[27]), .A2 (B_imm[27]), .A3 (B_imm[26]), .A4 (A_imm[28]));
INV_X1 i_527 (.ZN (n_463), .A (n_464));
OAI21_X1 i_526 (.ZN (n_462), .A (n_467), .B1 (n_463), .B2 (n_465));
NAND2_X1 i_525 (.ZN (n_461), .A1 (n_478), .A2 (n_480));
NAND2_X1 i_524 (.ZN (n_460), .A1 (n_461), .A2 (n_479));
OAI21_X1 i_523 (.ZN (n_459), .A (n_460), .B1 (n_8994), .B2 (n_8993));
NAND4_X1 i_522 (.ZN (n_458), .A1 (A_imm[29]), .A2 (n_461), .A3 (n_479), .A4 (B_imm[26]));
NAND2_X1 i_521 (.ZN (n_457), .A1 (n_459), .A2 (n_458));
XOR2_X1 i_520 (.Z (n_456), .A (n_462), .B (n_457));
NAND2_X1 i_519 (.ZN (n_455), .A1 (n_468), .A2 (n_456));
NAND2_X1 i_518 (.ZN (n_454), .A1 (n_469), .A2 (n_455));
XOR2_X1 i_517 (.Z (n_453), .A (n_454), .B (n_485));
INV_X1 i_516 (.ZN (n_452), .A (n_453));
NAND2_X1 i_515 (.ZN (n_451), .A1 (n_462), .A2 (n_458));
NAND2_X1 i_514 (.ZN (n_450), .A1 (n_451), .A2 (n_459));
INV_X1 i_513 (.ZN (n_449), .A (n_450));
NAND2_X1 i_512 (.ZN (n_448), .A1 (A_imm[27]), .A2 (B_imm[29]));
INV_X1 i_511 (.ZN (n_447), .A (n_448));
OAI22_X1 i_510 (.ZN (n_446), .A1 (n_9020), .A2 (n_9021), .B1 (n_8974), .B2 (n_9037));
NAND4_X1 i_509 (.ZN (n_445), .A1 (A_imm[28]), .A2 (B_imm[28]), .A3 (B_imm[25]), .A4 (opt_ipoPP_0));
NAND2_X1 i_508 (.ZN (n_444), .A1 (n_446), .A2 (n_445));
XNOR2_X1 i_507 (.ZN (n_443), .A (n_444), .B (n_447));
NOR2_X1 i_506 (.ZN (n_442), .A1 (n_449), .A2 (n_443));
NAND2_X1 i_505 (.ZN (n_441), .A1 (n_449), .A2 (n_443));
INV_X1 i_504 (.ZN (n_440), .A (n_441));
OR2_X1 i_503 (.ZN (n_439), .A1 (n_440), .A2 (n_442));
NAND2_X1 i_502 (.ZN (n_438), .A1 (A_imm[29]), .A2 (B_imm[27]));
INV_X1 i_501 (.ZN (n_437), .A (n_438));
OAI22_X1 i_500 (.ZN (n_436), .A1 (n_9038), .A2 (n_8794), .B1 (n_9004), .B2 (n_8972));
NAND4_X1 i_499 (.ZN (n_435), .A1 (B_imm[31]), .A2 (B_imm[30]), .A3 (A_imm[26]), .A4 (A_imm[25]));
NAND2_X1 i_498 (.ZN (n_434), .A1 (n_436), .A2 (n_435));
XNOR2_X1 i_497 (.ZN (n_433), .A (n_434), .B (n_437));
XNOR2_X1 i_496 (.ZN (n_432), .A (n_439), .B (n_433));
NOR2_X1 i_495 (.ZN (n_431), .A1 (n_452), .A2 (n_432));
NAND2_X1 i_494 (.ZN (n_430), .A1 (n_452), .A2 (n_432));
INV_X1 i_493 (.ZN (n_429), .A (n_430));
NOR2_X1 i_492 (.ZN (n_428), .A1 (n_429), .A2 (n_431));
INV_X1 i_491 (.ZN (n_427), .A (n_493));
NOR2_X1 i_490 (.ZN (n_426), .A1 (n_492), .A2 (n_427));
XNOR2_X1 i_489 (.ZN (n_425), .A (n_426), .B (n_489));
INV_X1 i_488 (.ZN (n_424), .A (n_545));
OAI21_X1 i_487 (.ZN (n_423), .A (n_547), .B1 (n_424), .B2 (n_550));
NAND2_X1 i_486 (.ZN (n_422), .A1 (n_467), .A2 (n_464));
XNOR2_X1 i_485 (.ZN (n_421), .A (n_422), .B (n_465));
INV_X1 i_484 (.ZN (n_420), .A (n_421));
OR2_X1 i_483 (.ZN (n_419), .A1 (n_420), .A2 (n_423));
NAND2_X1 i_482 (.ZN (n_418), .A1 (n_420), .A2 (n_423));
NAND2_X1 i_481 (.ZN (n_417), .A1 (n_499), .A2 (n_497));
XOR2_X1 i_480 (.Z (n_416), .A (n_498), .B (n_417));
NAND2_X1 i_479 (.ZN (n_415), .A1 (n_416), .A2 (n_418));
NAND2_X1 i_478 (.ZN (n_414), .A1 (n_415), .A2 (n_419));
NAND2_X1 i_477 (.ZN (n_413), .A1 (n_425), .A2 (n_414));
OR2_X1 i_476 (.ZN (n_412), .A1 (n_425), .A2 (n_414));
NAND2_X1 i_475 (.ZN (n_411), .A1 (n_469), .A2 (n_468));
XNOR2_X1 i_474 (.ZN (n_410), .A (n_411), .B (n_456));
NAND2_X1 i_473 (.ZN (n_409), .A1 (n_410), .A2 (n_412));
AND2_X1 i_472 (.ZN (n_408), .A1 (n_409), .A2 (n_413));
XOR2_X1 i_471 (.Z (n_407), .A (n_408), .B (n_428));
INV_X1 i_470 (.ZN (n_406), .A (n_568));
OAI21_X1 i_469 (.ZN (n_405), .A (n_566), .B1 (n_564), .B2 (n_406));
INV_X1 i_468 (.ZN (n_404), .A (n_582));
OAI21_X1 i_467 (.ZN (n_403), .A (n_581), .B1 (n_575), .B2 (n_404));
NAND2_X1 i_466 (.ZN (n_402), .A1 (n_405), .A2 (n_403));
OR2_X1 i_465 (.ZN (n_401), .A1 (n_405), .A2 (n_403));
NAND2_X1 i_464 (.ZN (n_400), .A1 (n_475), .A2 (n_473));
XNOR2_X1 i_463 (.ZN (n_399), .A (n_400), .B (n_474));
NAND2_X1 i_462 (.ZN (n_398), .A1 (n_399), .A2 (n_401));
NAND2_X1 i_461 (.ZN (n_397), .A1 (n_398), .A2 (n_402));
NAND2_X1 i_460 (.ZN (n_396), .A1 (n_419), .A2 (n_418));
XNOR2_X1 i_459 (.ZN (n_395), .A (n_396), .B (n_416));
NAND2_X1 i_458 (.ZN (n_394), .A1 (n_540), .A2 (n_537));
NAND2_X1 i_457 (.ZN (n_393), .A1 (n_541), .A2 (n_394));
NAND2_X1 i_456 (.ZN (n_392), .A1 (n_395), .A2 (n_393));
OR2_X1 i_455 (.ZN (n_391), .A1 (n_395), .A2 (n_393));
NAND2_X1 i_454 (.ZN (n_390), .A1 (n_570), .A2 (n_563));
NAND2_X1 i_453 (.ZN (n_389), .A1 (n_390), .A2 (n_571));
NAND2_X1 i_452 (.ZN (n_388), .A1 (n_391), .A2 (n_389));
NAND2_X1 i_451 (.ZN (n_387), .A1 (n_388), .A2 (n_392));
INV_X1 i_450 (.ZN (n_386), .A (n_387));
NAND2_X1 i_449 (.ZN (n_385), .A1 (n_386), .A2 (n_397));
NOR2_X1 i_448 (.ZN (n_384), .A1 (n_386), .A2 (n_397));
NAND2_X1 i_447 (.ZN (n_383), .A1 (n_412), .A2 (n_413));
XOR2_X1 i_446 (.Z (n_382), .A (n_383), .B (n_410));
INV_X1 i_445 (.ZN (n_381), .A (n_382));
OAI21_X1 i_444 (.ZN (n_380), .A (n_385), .B1 (n_381), .B2 (n_384));
NAND2_X1 i_443 (.ZN (n_379), .A1 (n_407), .A2 (n_380));
NAND2_X1 i_442 (.ZN (n_378), .A1 (n_527), .A2 (n_559));
NAND2_X1 i_441 (.ZN (n_377), .A1 (n_401), .A2 (n_402));
XNOR2_X1 i_440 (.ZN (n_376), .A (n_399), .B (n_377));
NAND2_X1 i_439 (.ZN (n_375), .A1 (n_532), .A2 (n_529));
NAND2_X1 i_438 (.ZN (n_374), .A1 (n_375), .A2 (n_533));
INV_X1 i_437 (.ZN (n_373), .A (n_374));
NOR2_X1 i_436 (.ZN (n_372), .A1 (n_373), .A2 (n_376));
INV_X1 i_435 (.ZN (n_371), .A (n_372));
NAND2_X1 i_434 (.ZN (n_370), .A1 (n_373), .A2 (n_376));
NAND2_X1 i_433 (.ZN (n_369), .A1 (n_371), .A2 (n_370));
NAND2_X1 i_432 (.ZN (n_368), .A1 (n_391), .A2 (n_392));
XOR2_X1 i_431 (.Z (n_367), .A (n_389), .B (n_368));
INV_X1 i_430 (.ZN (n_366), .A (n_367));
XNOR2_X1 i_429 (.ZN (n_365), .A (n_369), .B (n_366));
INV_X1 i_428 (.ZN (n_364), .A (n_365));
NAND3_X1 i_427 (.ZN (n_363), .A1 (n_364), .A2 (n_558), .A3 (n_378));
INV_X1 i_426 (.ZN (n_362), .A (n_384));
NAND2_X1 i_425 (.ZN (n_361), .A1 (n_362), .A2 (n_385));
XNOR2_X1 i_424 (.ZN (n_360), .A (n_381), .B (n_361));
INV_X1 i_423 (.ZN (n_359), .A (n_360));
NAND2_X1 i_422 (.ZN (n_358), .A1 (n_366), .A2 (n_370));
NAND2_X1 i_421 (.ZN (n_357), .A1 (n_358), .A2 (n_371));
INV_X1 i_420 (.ZN (n_356), .A (n_357));
NAND2_X1 i_419 (.ZN (n_355), .A1 (n_359), .A2 (n_356));
NAND3_X1 i_418 (.ZN (n_354), .A1 (n_363), .A2 (n_379), .A3 (n_355));
INV_X1 i_417 (.ZN (n_353), .A (n_354));
NAND2_X1 i_416 (.ZN (n_352), .A1 (n_8995), .A2 (n_8996));
XOR2_X1 i_415 (.Z (n_351), .A (n_8981), .B (n_352));
INV_X1 i_414 (.ZN (n_350), .A (n_351));
NAND2_X1 i_413 (.ZN (n_349), .A1 (n_9019), .A2 (n_9016));
XNOR2_X1 i_412 (.ZN (n_348), .A (n_349), .B (n_9017));
INV_X1 i_411 (.ZN (n_347), .A (n_348));
NAND2_X1 i_410 (.ZN (n_346), .A1 (n_350), .A2 (n_347));
NOR2_X1 i_409 (.ZN (n_345), .A1 (n_350), .A2 (n_347));
AOI22_X1 i_408 (.ZN (n_344), .A1 (A_imm[29]), .A2 (B_imm[28]), .B1 (B_imm[31]), .B2 (A_imm[26]));
INV_X1 i_407 (.ZN (n_343), .A (n_445));
OAI21_X1 i_406 (.ZN (n_342), .A (n_446), .B1 (n_447), .B2 (n_343));
NAND4_X1 i_405 (.ZN (n_341), .A1 (A_imm[29]), .A2 (B_imm[31]), .A3 (B_imm[28]), .A4 (A_imm[26]));
AOI21_X1 i_404 (.ZN (n_340), .A (n_344), .B1 (n_342), .B2 (n_341));
INV_X1 i_403 (.ZN (n_339), .A (n_340));
NAND2_X1 i_402 (.ZN (n_338), .A1 (n_9002), .A2 (n_8999));
XNOR2_X1 i_401 (.ZN (n_337), .A (n_338), .B (n_9000));
INV_X1 i_400 (.ZN (n_336), .A (n_337));
NAND2_X1 i_399 (.ZN (n_335), .A1 (n_336), .A2 (n_339));
INV_X1 i_398 (.ZN (n_334), .A (n_335));
NAND2_X1 i_397 (.ZN (n_333), .A1 (n_337), .A2 (n_340));
INV_X1 i_396 (.ZN (n_332), .A (n_435));
OAI21_X1 i_395 (.ZN (n_331), .A (n_436), .B1 (n_437), .B2 (n_332));
OAI21_X1 i_394 (.ZN (n_330), .A (n_331), .B1 (CLOCK_opt_ipo_n433), .B2 (n_9005));
OR3_X1 i_393 (.ZN (n_329), .A1 (n_331), .A2 (CLOCK_opt_ipo_n433), .A3 (n_9005));
NAND2_X1 i_392 (.ZN (n_328), .A1 (n_8992), .A2 (n_8989));
XNOR2_X1 i_391 (.ZN (n_327), .A (n_328), .B (n_8990));
INV_X1 i_390 (.ZN (n_326), .A (n_327));
NAND2_X1 i_389 (.ZN (n_325), .A1 (n_329), .A2 (n_326));
NAND2_X1 i_388 (.ZN (n_324), .A1 (n_325), .A2 (n_330));
AOI21_X1 i_387 (.ZN (n_323), .A (n_334), .B1 (n_324), .B2 (n_333));
OAI21_X1 i_386 (.ZN (n_322), .A (n_346), .B1 (n_345), .B2 (n_323));
NAND2_X1 i_385 (.ZN (n_321), .A1 (n_9009), .A2 (n_9008));
XNOR2_X1 i_384 (.ZN (n_320), .A (n_321), .B (n_8979));
NAND2_X1 i_383 (.ZN (n_319), .A1 (n_322), .A2 (n_320));
INV_X1 i_382 (.ZN (n_318), .A (n_346));
NOR2_X1 i_381 (.ZN (n_317), .A1 (n_318), .A2 (n_345));
XOR2_X1 i_380 (.Z (n_316), .A (n_323), .B (n_317));
INV_X1 i_379 (.ZN (n_315), .A (n_316));
NAND2_X1 i_378 (.ZN (n_314), .A1 (n_8983), .A2 (n_8986));
XNOR2_X1 i_377 (.ZN (n_313), .A (n_314), .B (n_8984));
INV_X1 i_376 (.ZN (n_312), .A (n_344));
NAND2_X1 i_375 (.ZN (n_311), .A1 (n_312), .A2 (n_341));
XOR2_X1 i_374 (.Z (n_310), .A (n_342), .B (n_311));
INV_X1 i_373 (.ZN (n_309), .A (n_310));
INV_X1 i_372 (.ZN (n_308), .A (n_504));
OAI21_X1 i_371 (.ZN (n_307), .A (n_507), .B1 (n_308), .B2 (n_519));
OR2_X1 i_370 (.ZN (n_306), .A1 (n_309), .A2 (n_307));
NAND2_X1 i_369 (.ZN (n_305), .A1 (n_309), .A2 (n_307));
INV_X1 i_368 (.ZN (n_304), .A (n_305));
INV_X1 i_367 (.ZN (n_303), .A (n_433));
OAI21_X1 i_366 (.ZN (n_302), .A (n_441), .B1 (n_303), .B2 (n_442));
INV_X1 i_365 (.ZN (n_301), .A (n_302));
OAI21_X1 i_364 (.ZN (n_300), .A (n_306), .B1 (n_301), .B2 (n_304));
NAND2_X1 i_363 (.ZN (n_299), .A1 (n_300), .A2 (n_313));
OR2_X1 i_362 (.ZN (n_298), .A1 (n_300), .A2 (n_313));
INV_X1 i_361 (.ZN (n_297), .A (n_324));
NAND2_X1 i_360 (.ZN (n_296), .A1 (n_335), .A2 (n_333));
XNOR2_X1 i_359 (.ZN (n_295), .A (n_297), .B (n_296));
NAND2_X1 i_358 (.ZN (n_294), .A1 (n_298), .A2 (n_295));
NAND2_X1 i_357 (.ZN (n_293), .A1 (n_294), .A2 (n_299));
INV_X1 i_356 (.ZN (n_292), .A (n_293));
NAND2_X1 i_355 (.ZN (n_291), .A1 (n_315), .A2 (n_292));
NAND2_X1 i_354 (.ZN (n_290), .A1 (n_291), .A2 (n_319));
INV_X1 i_353 (.ZN (n_289), .A (n_290));
INV_X1 i_352 (.ZN (n_288), .A (n_295));
NAND2_X1 i_351 (.ZN (n_287), .A1 (n_298), .A2 (n_299));
XNOR2_X1 i_350 (.ZN (n_286), .A (n_287), .B (n_288));
NAND2_X1 i_349 (.ZN (n_285), .A1 (n_329), .A2 (n_330));
XNOR2_X1 i_348 (.ZN (n_284), .A (n_285), .B (n_326));
NAND2_X1 i_347 (.ZN (n_283), .A1 (n_454), .A2 (n_487));
NAND2_X1 i_346 (.ZN (n_282), .A1 (n_283), .A2 (n_486));
INV_X1 i_345 (.ZN (n_281), .A (n_282));
NOR2_X1 i_344 (.ZN (n_280), .A1 (n_281), .A2 (n_284));
INV_X1 i_343 (.ZN (n_279), .A (n_280));
NAND2_X1 i_342 (.ZN (n_278), .A1 (n_281), .A2 (n_284));
NAND2_X1 i_341 (.ZN (n_277), .A1 (n_306), .A2 (n_305));
XNOR2_X1 i_340 (.ZN (n_276), .A (n_277), .B (n_301));
INV_X1 i_339 (.ZN (n_275), .A (n_276));
NAND2_X1 i_338 (.ZN (n_274), .A1 (n_275), .A2 (n_278));
NAND3_X1 i_337 (.ZN (n_273), .A1 (n_286), .A2 (n_279), .A3 (n_274));
NAND2_X1 i_336 (.ZN (n_272), .A1 (n_279), .A2 (n_278));
XNOR2_X1 i_335 (.ZN (n_271), .A (n_272), .B (n_275));
OAI21_X1 i_334 (.ZN (n_270), .A (n_430), .B1 (n_431), .B2 (n_408));
OR2_X1 i_333 (.ZN (n_269), .A1 (n_270), .A2 (n_271));
NAND3_X1 i_332 (.ZN (n_268), .A1 (n_269), .A2 (n_289), .A3 (n_273));
INV_X1 i_331 (.ZN (n_267), .A (n_268));
NAND3_X1 i_330 (.ZN (n_266), .A1 (n_353), .A2 (n_521), .A3 (n_267));
NAND3_X1 i_329 (.ZN (n_265), .A1 (n_353), .A2 (n_526), .A3 (n_523));
INV_X1 i_328 (.ZN (n_264), .A (n_355));
NAND2_X1 i_327 (.ZN (n_263), .A1 (n_360), .A2 (n_357));
NAND2_X1 i_326 (.ZN (n_262), .A1 (n_378), .A2 (n_558));
NAND2_X1 i_325 (.ZN (n_261), .A1 (n_262), .A2 (n_365));
OAI21_X1 i_324 (.ZN (n_260), .A (n_263), .B1 (n_261), .B2 (n_264));
NAND2_X1 i_323 (.ZN (n_259), .A1 (n_260), .A2 (n_379));
OR2_X1 i_322 (.ZN (n_258), .A1 (n_407), .A2 (n_380));
NAND3_X1 i_321 (.ZN (n_257), .A1 (n_265), .A2 (n_259), .A3 (n_258));
NAND2_X1 i_320 (.ZN (n_256), .A1 (n_271), .A2 (n_270));
NAND2_X1 i_319 (.ZN (n_255), .A1 (n_289), .A2 (n_273));
INV_X1 i_318 (.ZN (n_254), .A (n_291));
INV_X1 i_317 (.ZN (n_253), .A (n_286));
INV_X1 i_316 (.ZN (n_252), .A (n_274));
OAI21_X1 i_315 (.ZN (n_251), .A (n_253), .B1 (n_280), .B2 (n_252));
OR2_X1 i_314 (.ZN (n_250), .A1 (n_322), .A2 (n_320));
NAND2_X1 i_313 (.ZN (n_249), .A1 (n_316), .A2 (n_293));
OAI211_X1 i_312 (.ZN (n_248), .A (n_250), .B (n_249), .C1 (n_254), .C2 (n_251));
NAND2_X1 i_311 (.ZN (n_247), .A1 (n_248), .A2 (n_319));
OAI21_X1 i_310 (.ZN (n_246), .A (n_247), .B1 (n_256), .B2 (n_255));
AOI21_X1 i_309 (.ZN (n_245), .A (n_246), .B1 (n_257), .B2 (n_267));
OAI21_X2 i_308 (.ZN (n_244), .A (n_245), .B1 (n_586), .B2 (n_266));
AOI21_X1 i_307 (.ZN (n_243), .A (n_8976), .B1 (n_244), .B2 (n_8975));
OAI21_X1 i_306 (.ZN (Res_imm[63]), .A (n_9027), .B1 (n_243), .B2 (n_9025));
INV_X1 i_305 (.ZN (n_242), .A (n_8976));
NAND2_X2 i_304 (.ZN (n_241), .A1 (n_244), .A2 (n_8975));
NAND2_X1 i_303 (.ZN (n_240), .A1 (n_9027), .A2 (n_9026));
AOI21_X2 i_302 (.ZN (n_239), .A (n_240), .B1 (n_241), .B2 (n_242));
NAND3_X1 i_301 (.ZN (n_238), .A1 (n_241), .A2 (n_242), .A3 (n_240));
NOR2_X2 i_299 (.ZN (Res_imm[62]), .A1 (CLOCK_opt_ipo_n345), .A2 (n_239));
NAND2_X1 i_298 (.ZN (n_236), .A1 (n_242), .A2 (n_8975));
INV_X1 i_297 (.ZN (n_235), .A (n_236));
XNOR2_X1 i_296 (.ZN (n_234), .A (n_244), .B (n_235));
INV_X1 i_295 (.ZN (Res_imm[61]), .A (n_234));
NAND2_X1 i_294 (.ZN (n_233), .A1 (n_250), .A2 (n_319));
INV_X1 i_293 (.ZN (n_232), .A (n_233));
NAND2_X1 i_292 (.ZN (n_231), .A1 (n_353), .A2 (n_521));
INV_X1 i_291 (.ZN (n_230), .A (n_257));
OAI21_X4 i_290 (.ZN (n_229), .A (n_230), .B1 (n_586), .B2 (n_231));
NAND2_X1 i_289 (.ZN (n_228), .A1 (n_269), .A2 (n_256));
INV_X1 i_288 (.ZN (n_227), .A (n_228));
NAND4_X1 i_287 (.ZN (n_226), .A1 (n_227), .A2 (n_273), .A3 (n_251), .A4 (n_249));
NAND2_X1 i_286 (.ZN (n_225), .A1 (n_269), .A2 (n_273));
NAND2_X1 i_285 (.ZN (n_224), .A1 (n_225), .A2 (n_251));
INV_X1 i_284 (.ZN (n_223), .A (n_224));
OAI21_X1 i_283 (.ZN (n_222), .A (n_249), .B1 (n_223), .B2 (n_254));
OAI21_X1 i_282 (.ZN (n_221), .A (n_222), .B1 (n_229), .B2 (n_226));
NAND2_X1 i_281 (.ZN (n_220), .A1 (n_221), .A2 (n_232));
OAI211_X1 i_280 (.ZN (n_219), .A (n_233), .B (n_222), .C1 (n_229), .C2 (n_226));
NAND2_X1 i_279 (.ZN (Res_imm[60]), .A1 (n_220), .A2 (n_219));
NAND2_X1 i_278 (.ZN (n_218), .A1 (n_227), .A2 (n_251));
OAI21_X1 i_277 (.ZN (n_217), .A (n_224), .B1 (n_229), .B2 (n_218));
NAND2_X1 i_276 (.ZN (n_216), .A1 (n_291), .A2 (n_249));
INV_X1 i_275 (.ZN (n_215), .A (n_216));
NAND2_X1 i_274 (.ZN (n_214), .A1 (n_217), .A2 (n_215));
OAI211_X1 i_273 (.ZN (n_213), .A (n_224), .B (n_216), .C1 (n_229), .C2 (n_218));
NAND2_X1 i_272 (.ZN (Res_imm[59]), .A1 (n_214), .A2 (n_213));
NAND2_X1 i_271 (.ZN (n_212), .A1 (n_229), .A2 (n_269));
NAND4_X1 i_270 (.ZN (n_211), .A1 (n_212), .A2 (n_273), .A3 (n_256), .A4 (n_251));
NAND2_X1 i_269 (.ZN (n_210), .A1 (n_251), .A2 (n_273));
NAND2_X1 i_268 (.ZN (n_209), .A1 (n_212), .A2 (n_256));
NAND2_X1 i_267 (.ZN (n_208), .A1 (n_209), .A2 (n_210));
NAND2_X2 i_266 (.ZN (Res_imm[58]), .A1 (n_208), .A2 (n_211));
XNOR2_X2 i_265 (.ZN (CLOCK_opt_ipo_n452), .A (n_229), .B (n_227));
NAND2_X1 i_263 (.ZN (n_206), .A1 (n_258), .A2 (n_379));
INV_X1 i_262 (.ZN (n_205), .A (n_206));
INV_X1 i_261 (.ZN (n_204), .A (n_521));
NAND2_X1 i_260 (.ZN (n_203), .A1 (n_526), .A2 (n_523));
OAI21_X2 i_259 (.ZN (n_202), .A (n_203), .B1 (n_586), .B2 (n_204));
NAND2_X1 i_258 (.ZN (n_201), .A1 (n_363), .A2 (n_261));
INV_X1 i_257 (.ZN (n_200), .A (n_201));
NAND2_X1 i_256 (.ZN (n_199), .A1 (n_200), .A2 (n_263));
INV_X1 i_255 (.ZN (n_198), .A (n_363));
OAI21_X1 i_254 (.ZN (n_197), .A (n_263), .B1 (n_198), .B2 (n_264));
OAI21_X1 i_253 (.ZN (n_196), .A (n_197), .B1 (n_202), .B2 (n_199));
NAND2_X1 i_252 (.ZN (n_195), .A1 (n_196), .A2 (n_205));
OAI211_X1 i_251 (.ZN (n_194), .A (n_206), .B (n_197), .C1 (n_202), .C2 (n_199));
NAND2_X2 i_250 (.ZN (Res_imm[56]), .A1 (n_195), .A2 (n_194));
NAND2_X1 i_249 (.ZN (n_193), .A1 (n_202), .A2 (n_363));
NAND4_X1 i_248 (.ZN (n_192), .A1 (n_193), .A2 (n_355), .A3 (n_263), .A4 (n_261));
NAND2_X1 i_247 (.ZN (n_191), .A1 (n_355), .A2 (n_263));
NAND2_X1 i_246 (.ZN (n_190), .A1 (n_193), .A2 (n_261));
NAND2_X2 i_245 (.ZN (n_189), .A1 (n_190), .A2 (n_191));
NAND2_X4 i_244 (.ZN (Res_imm[55]), .A1 (n_189), .A2 (n_192));
XNOR2_X1 i_243 (.ZN (n_188), .A (n_202), .B (n_200));
INV_X2 i_242 (.ZN (Res_imm[54]), .A (n_188));
NAND2_X1 i_241 (.ZN (n_187), .A1 (n_521), .A2 (n_203));
XOR2_X1 i_240 (.Z (Res_imm[53]), .A (n_187), .B (n_586));
INV_X1 i_239 (.ZN (n_186), .A (n_761));
INV_X1 i_238 (.ZN (n_185), .A (n_589));
AOI21_X2 i_237 (.ZN (n_184), .A (n_185), .B1 (n_951), .B2 (n_855));
OAI21_X2 i_236 (.ZN (n_183), .A (n_594), .B1 (n_184), .B2 (n_186));
NAND2_X1 i_235 (.ZN (n_182), .A1 (n_183), .A2 (n_678));
NAND4_X1 i_234 (.ZN (n_181), .A1 (n_182), .A2 (n_600), .A3 (n_593), .A4 (n_588));
NAND2_X1 i_233 (.ZN (n_180), .A1 (n_600), .A2 (n_588));
NAND2_X1 i_232 (.ZN (n_179), .A1 (n_182), .A2 (n_593));
NAND2_X1 i_231 (.ZN (n_178), .A1 (n_179), .A2 (n_180));
NAND2_X4 i_230 (.ZN (Res_imm[52]), .A1 (n_178), .A2 (n_181));
NAND2_X1 i_229 (.ZN (n_177), .A1 (n_593), .A2 (n_678));
INV_X1 i_228 (.ZN (n_176), .A (n_177));
XNOR2_X2 i_227 (.ZN (Res_imm[51]), .A (n_183), .B (n_176));
NAND2_X1 i_225 (.ZN (n_174), .A1 (n_761), .A2 (n_594));
XOR2_X2 i_224 (.Z (Res_imm[50]), .A (n_174), .B (n_184));
NAND2_X1 i_223 (.ZN (n_173), .A1 (n_855), .A2 (n_589));
XOR2_X1 i_222 (.Z (n_172), .A (n_173), .B (n_951));
INV_X1 i_221 (.ZN (Res_imm[49]), .A (n_172));
NAND2_X1 i_220 (.ZN (n_171), .A1 (n_5112), .A2 (n_5121));
NAND2_X1 i_219 (.ZN (n_170), .A1 (n_959), .A2 (n_958));
NAND2_X1 i_218 (.ZN (n_169), .A1 (n_954), .A2 (n_5139));
INV_X1 i_217 (.ZN (n_168), .A (n_169));
NAND2_X1 i_216 (.ZN (n_167), .A1 (n_964), .A2 (n_5112));
INV_X1 i_215 (.ZN (n_166), .A (n_167));
NAND3_X1 i_214 (.ZN (n_165), .A1 (n_6934), .A2 (n_5724), .A3 (CLOCK_opt_ipo_n351));
INV_X1 i_213 (.ZN (n_164), .A (n_967));
AOI21_X4 i_212 (.ZN (n_163), .A (n_3981), .B1 (n_1002), .B2 (CLOCK_opt_ipo_n326));
OAI21_X2 i_211 (.ZN (n_162), .A (n_164), .B1 (n_163), .B2 (n_165));
NAND2_X1 i_210 (.ZN (n_161), .A1 (n_162), .A2 (n_5505));
NAND3_X1 i_209 (.ZN (n_160), .A1 (n_161), .A2 (n_961), .A3 (n_166));
INV_X1 i_208 (.ZN (n_159), .A (n_160));
OAI211_X1 i_207 (.ZN (n_158), .A (n_170), .B (n_168), .C1 (n_159), .C2 (n_171));
OAI21_X1 i_206 (.ZN (n_157), .A (n_170), .B1 (n_159), .B2 (n_171));
NAND2_X1 i_205 (.ZN (n_156), .A1 (n_157), .A2 (n_169));
NAND2_X2 i_204 (.ZN (Res_imm[48]), .A1 (n_156), .A2 (n_158));
INV_X1 i_203 (.ZN (n_155), .A (n_961));
AOI21_X1 i_202 (.ZN (n_154), .A (n_155), .B1 (n_162), .B2 (n_5505));
NAND2_X1 i_201 (.ZN (n_153), .A1 (n_154), .A2 (n_964));
NAND2_X1 i_200 (.ZN (n_152), .A1 (n_153), .A2 (n_5112));
NAND3_X1 i_199 (.ZN (n_151), .A1 (n_152), .A2 (n_5121), .A3 (n_170));
NAND2_X1 i_198 (.ZN (n_150), .A1 (n_170), .A2 (n_5121));
NAND3_X1 i_197 (.ZN (n_149), .A1 (n_153), .A2 (n_5112), .A3 (n_150));
NAND2_X2 i_196 (.ZN (Res_imm[47]), .A1 (n_151), .A2 (n_149));
XNOR2_X1 i_195 (.ZN (Res_imm[46]), .A (n_154), .B (n_166));
NAND2_X1 i_194 (.ZN (n_148), .A1 (n_961), .A2 (n_5505));
XOR2_X1 i_193 (.Z (n_147), .A (n_148), .B (n_162));
INV_X1 i_192 (.ZN (Res_imm[45]), .A (n_147));
NAND2_X1 i_191 (.ZN (n_146), .A1 (n_6936), .A2 (n_6943));
INV_X1 i_190 (.ZN (n_145), .A (n_972));
INV_X1 i_189 (.ZN (n_144), .A (n_6964));
NOR2_X1 i_188 (.ZN (n_143), .A1 (n_144), .A2 (n_971));
NAND2_X1 i_187 (.ZN (n_142), .A1 (n_977), .A2 (n_6936));
INV_X1 i_186 (.ZN (n_141), .A (n_142));
NAND2_X1 i_185 (.ZN (n_140), .A1 (CLOCK_opt_ipo_n351), .A2 (n_5724));
OAI21_X2 i_184 (.ZN (n_139), .A (n_980), .B1 (n_163), .B2 (n_140));
NAND2_X1 i_183 (.ZN (n_138), .A1 (n_139), .A2 (n_7465));
NAND3_X1 i_182 (.ZN (n_137), .A1 (n_138), .A2 (n_976), .A3 (n_141));
INV_X1 i_181 (.ZN (n_136), .A (n_137));
OAI211_X2 i_180 (.ZN (n_135), .A (n_145), .B (n_143), .C1 (n_136), .C2 (n_146));
INV_X1 i_179 (.ZN (n_134), .A (n_976));
AOI21_X4 i_178 (.ZN (n_133), .A (n_134), .B1 (n_139), .B2 (n_7465));
AOI21_X1 i_177 (.ZN (n_132), .A (n_146), .B1 (n_133), .B2 (n_141));
INV_X1 sgo__sro_c300 (.ZN (sgo__sro_n158), .A (n_7691));
NAND2_X2 i_175 (.ZN (Res_imm[44]), .A1 (n_131), .A2 (n_135));
INV_X1 i_174 (.ZN (n_130), .A (n_6936));
OAI21_X4 i_173 (.ZN (n_129), .A (n_977), .B1 (n_133), .B2 (n_130));
INV_X1 i_172 (.ZN (n_128), .A (n_129));
NAND3_X2 i_171 (.ZN (n_127), .A1 (n_128), .A2 (n_6943), .A3 (n_145));
INV_X1 i_170 (.ZN (n_126), .A (n_6943));
OAI21_X1 i_169 (.ZN (n_125), .A (n_129), .B1 (n_126), .B2 (n_972));
NAND2_X4 i_168 (.ZN (Res_imm[43]), .A1 (n_127), .A2 (n_125));
XNOR2_X2 i_167 (.ZN (Res_imm[42]), .A (n_133), .B (n_141));
NAND2_X1 i_166 (.ZN (n_124), .A1 (n_7465), .A2 (n_976));
XOR2_X1 i_165 (.Z (CLOCK_opt_ipo_n363), .A (n_124), .B (n_139));
INV_X1 i_163 (.ZN (n_122), .A (n_5658));
INV_X1 i_162 (.ZN (n_121), .A (n_990));
INV_X1 i_161 (.ZN (n_120), .A (n_5724));
OAI21_X2 i_160 (.ZN (n_119), .A (n_993), .B1 (n_163), .B2 (n_120));
AOI21_X2 i_159 (.ZN (n_118), .A (n_121), .B1 (n_119), .B2 (n_5689));
OAI21_X2 i_158 (.ZN (n_117), .A (n_985), .B1 (n_118), .B2 (n_122));
INV_X1 i_157 (.ZN (n_116), .A (n_117));
NAND3_X1 i_156 (.ZN (n_115), .A1 (n_116), .A2 (n_5666), .A3 (n_982));
INV_X1 i_155 (.ZN (n_114), .A (n_982));
OAI21_X1 i_154 (.ZN (n_113), .A (n_117), .B1 (n_988), .B2 (n_114));
NAND2_X2 i_153 (.ZN (Res_imm[40]), .A1 (n_115), .A2 (n_113));
NAND2_X1 i_152 (.ZN (n_112), .A1 (n_985), .A2 (n_5658));
XOR2_X1 i_151 (.Z (Res_imm[39]), .A (n_112), .B (n_118));
NAND2_X1 i_150 (.ZN (n_111), .A1 (n_990), .A2 (n_5689));
XOR2_X1 i_149 (.Z (n_110), .A (n_111), .B (n_119));
INV_X1 i_148 (.ZN (Res_imm[38]), .A (n_110));
NAND2_X1 i_147 (.ZN (n_109), .A1 (n_5724), .A2 (n_993));
XOR2_X1 i_146 (.Z (Res_imm[37]), .A (n_109), .B (n_163));
NAND2_X1 i_145 (.ZN (n_108), .A1 (n_3984), .A2 (n_4222));
INV_X1 i_144 (.ZN (n_107), .A (n_3986));
INV_X1 i_143 (.ZN (n_106), .A (n_4252));
INV_X1 i_142 (.ZN (n_105), .A (n_3992));
AOI21_X1 i_141 (.ZN (n_104), .A (n_105), .B1 (n_1002), .B2 (n_1000));
OAI21_X2 i_140 (.ZN (n_103), .A (n_4217), .B1 (n_104), .B2 (n_106));
AOI21_X1 i_139 (.ZN (n_102), .A (n_107), .B1 (n_103), .B2 (n_4229));
XOR2_X1 i_138 (.Z (Res_imm[36]), .A (n_108), .B (n_102));
NAND2_X1 i_137 (.ZN (n_101), .A1 (n_3986), .A2 (n_4229));
XNOR2_X1 i_136 (.ZN (Res_imm[35]), .A (n_103), .B (n_101));
NAND2_X1 i_135 (.ZN (n_100), .A1 (n_4252), .A2 (n_4217));
XNOR2_X1 i_134 (.ZN (n_99), .A (n_104), .B (n_100));
INV_X2 i_133 (.ZN (Res_imm[34]), .A (n_99));
NAND2_X1 i_132 (.ZN (n_98), .A1 (n_1000), .A2 (n_3992));
XNOR2_X2 i_131 (.ZN (Res_imm[33]), .A (n_1002), .B (n_98));
NAND2_X1 i_130 (.ZN (n_97), .A1 (n_1005), .A2 (n_1037));
INV_X1 i_129 (.ZN (n_96), .A (n_1019));
NAND3_X1 i_128 (.ZN (n_95), .A1 (n_1020), .A2 (n_1038), .A3 (n_1023));
INV_X1 i_127 (.ZN (n_94), .A (n_95));
INV_X1 i_126 (.ZN (n_93), .A (n_1024));
NAND3_X1 i_125 (.ZN (n_92), .A1 (n_1138), .A2 (n_1131), .A3 (n_1124));
NAND3_X1 i_124 (.ZN (n_91), .A1 (n_92), .A2 (n_2323), .A3 (n_2104));
NAND3_X1 i_123 (.ZN (n_90), .A1 (n_91), .A2 (n_1119), .A3 (n_1114));
NAND3_X1 i_122 (.ZN (n_89), .A1 (n_90), .A2 (n_3077), .A3 (CLOCK_opt_ipo_n333));
NAND2_X2 i_121 (.ZN (n_88), .A1 (n_89), .A2 (n_1102));
AND2_X2 i_120 (.ZN (n_87), .A1 (n_88), .A2 (n_1060));
OAI21_X1 i_119 (.ZN (n_86), .A (n_93), .B1 (n_87), .B2 (n_1012));
NAND2_X1 i_118 (.ZN (n_85), .A1 (n_86), .A2 (n_1009));
OAI21_X2 i_117 (.ZN (n_84), .A (n_96), .B1 (n_85), .B2 (n_94));
XOR2_X2 i_116 (.Z (Res_imm[32]), .A (n_97), .B (n_84));
NAND2_X1 i_115 (.ZN (n_83), .A1 (n_96), .A2 (n_95));
XNOR2_X2 i_114 (.ZN (Res_imm[31]), .A (n_85), .B (n_83));
NOR2_X1 i_113 (.ZN (n_82), .A1 (n_87), .A2 (n_1012));
NAND2_X1 i_112 (.ZN (n_81), .A1 (n_93), .A2 (n_1009));
XNOR2_X1 i_111 (.ZN (n_80), .A (n_82), .B (n_81));
INV_X1 i_110 (.ZN (Res_imm[30]), .A (n_80));
NAND2_X1 i_109 (.ZN (n_79), .A1 (n_1013), .A2 (n_1060));
XNOR2_X1 i_108 (.ZN (Res_imm[29]), .A (n_88), .B (n_79));
NAND2_X1 i_107 (.ZN (n_78), .A1 (n_3077), .A2 (n_1105));
INV_X1 i_106 (.ZN (n_77), .A (n_1104));
INV_X1 i_105 (.ZN (n_76), .A (n_2769));
NAND4_X1 i_104 (.ZN (n_75), .A1 (n_2931), .A2 (n_2923), .A3 (n_2775), .A4 (n_2771));
NAND3_X1 i_103 (.ZN (n_74), .A1 (n_2774), .A2 (n_2636), .A3 (n_2633));
INV_X1 i_102 (.ZN (n_73), .A (n_74));
AOI21_X1 i_101 (.ZN (n_72), .A (n_73), .B1 (n_90), .B2 (n_2631));
OAI21_X1 i_100 (.ZN (n_71), .A (n_75), .B1 (n_72), .B2 (n_76));
AOI21_X1 i_99 (.ZN (n_70), .A (n_77), .B1 (n_71), .B2 (n_2928));
XNOR2_X1 i_98 (.ZN (n_69), .A (n_70), .B (n_78));
INV_X1 i_97 (.ZN (Res_imm[28]), .A (n_69));
NAND2_X1 i_96 (.ZN (n_68), .A1 (n_2928), .A2 (n_1104));
XNOR2_X2 i_95 (.ZN (Res_imm[27]), .A (n_71), .B (n_68));
NAND2_X1 i_94 (.ZN (n_67), .A1 (n_75), .A2 (n_2769));
XNOR2_X1 i_93 (.ZN (n_66), .A (n_72), .B (n_67));
INV_X1 i_92 (.ZN (Res_imm[26]), .A (n_66));
NAND2_X1 i_91 (.ZN (n_65), .A1 (n_2631), .A2 (n_74));
XNOR2_X1 i_90 (.ZN (Res_imm[25]), .A (n_90), .B (n_65));
XOR2_X1 i_89 (.Z (n_64), .A (n_2333), .B (n_1121));
INV_X1 i_88 (.ZN (n_63), .A (n_2339));
INV_X1 i_87 (.ZN (n_62), .A (n_2329));
NAND2_X1 i_86 (.ZN (n_61), .A1 (n_62), .A2 (n_63));
INV_X1 i_85 (.ZN (n_60), .A (n_61));
NAND2_X1 i_84 (.ZN (n_59), .A1 (n_1117), .A2 (n_2217));
INV_X1 i_83 (.ZN (n_58), .A (n_92));
OAI21_X1 i_82 (.ZN (n_57), .A (n_1116), .B1 (n_58), .B2 (CLOCK_opt_ipo_n425));
INV_X1 i_81 (.ZN (n_56), .A (n_57));
OAI21_X1 i_80 (.ZN (n_55), .A (n_59), .B1 (n_56), .B2 (n_2215));
AOI21_X1 i_79 (.ZN (n_54), .A (n_60), .B1 (n_55), .B2 (n_2328));
XNOR2_X1 i_78 (.ZN (n_53), .A (n_54), .B (n_64));
INV_X1 i_77 (.ZN (Res_imm[24]), .A (n_53));
NAND2_X1 i_76 (.ZN (n_52), .A1 (n_61), .A2 (n_2328));
XOR2_X1 i_75 (.Z (n_51), .A (n_52), .B (n_55));
INV_X1 i_74 (.ZN (Res_imm[23]), .A (n_51));
INV_X1 i_73 (.ZN (n_50), .A (n_2215));
NAND2_X1 i_72 (.ZN (n_49), .A1 (n_50), .A2 (n_59));
XNOR2_X1 i_71 (.ZN (n_48), .A (n_56), .B (n_49));
INV_X1 i_70 (.ZN (Res_imm[22]), .A (n_48));
INV_X1 i_69 (.ZN (n_47), .A (CLOCK_opt_ipo_n425));
NAND2_X1 i_68 (.ZN (n_46), .A1 (n_47), .A2 (n_1116));
XNOR2_X1 i_67 (.ZN (Res_imm[21]), .A (n_92), .B (n_46));
NAND3_X1 i_66 (.ZN (n_45), .A1 (n_1223), .A2 (n_1222), .A3 (n_1185));
NAND2_X1 i_65 (.ZN (n_44), .A1 (n_1129), .A2 (n_45));
NOR2_X1 i_64 (.ZN (n_43), .A1 (n_1185), .A2 (n_1133));
NAND2_X1 i_63 (.ZN (n_42), .A1 (n_43), .A2 (n_1161));
INV_X1 i_62 (.ZN (n_41), .A (n_42));
NAND3_X1 i_61 (.ZN (n_40), .A1 (n_1153), .A2 (n_1162), .A3 (n_1145));
INV_X1 i_60 (.ZN (n_39), .A (n_1140));
NAND2_X1 i_59 (.ZN (n_38), .A1 (n_1141), .A2 (n_1146));
INV_X1 i_58 (.ZN (n_37), .A (n_38));
NAND2_X1 i_57 (.ZN (n_36), .A1 (n_37), .A2 (n_1795));
INV_X1 i_56 (.ZN (n_35), .A (n_36));
OAI21_X1 i_55 (.ZN (n_34), .A (n_39), .B1 (n_1226), .B2 (n_35));
AOI21_X1 i_54 (.ZN (n_33), .A (n_1144), .B1 (n_34), .B2 (n_40));
OAI21_X1 i_53 (.ZN (n_32), .A (n_1128), .B1 (n_33), .B2 (n_41));
XOR2_X1 i_52 (.Z (Res_imm[20]), .A (n_44), .B (n_32));
NAND2_X1 i_51 (.ZN (n_31), .A1 (n_42), .A2 (n_1128));
XNOR2_X1 i_50 (.ZN (Res_imm[19]), .A (n_33), .B (n_31));
INV_X1 i_49 (.ZN (n_30), .A (n_1144));
NAND2_X1 i_48 (.ZN (n_29), .A1 (n_30), .A2 (n_40));
XNOR2_X1 i_47 (.ZN (n_28), .A (n_34), .B (n_29));
INV_X1 i_46 (.ZN (Res_imm[18]), .A (n_28));
NAND2_X1 i_45 (.ZN (n_27), .A1 (n_39), .A2 (n_36));
XNOR2_X1 i_44 (.ZN (Res_imm[17]), .A (n_1226), .B (n_27));
NAND2_X1 i_43 (.ZN (n_26), .A1 (n_1718), .A2 (n_1229));
AND2_X1 i_42 (.ZN (n_25), .A1 (n_1235), .A2 (n_1233));
XOR2_X2 i_41 (.Z (Res_imm[16]), .A (n_26), .B (n_25));
NAND2_X1 i_40 (.ZN (n_24), .A1 (n_1233), .A2 (n_1240));
NAND2_X1 i_39 (.ZN (n_23), .A1 (n_1243), .A2 (n_1238));
XOR2_X1 i_38 (.Z (Res_imm[15]), .A (n_24), .B (n_23));
OAI21_X1 i_37 (.ZN (n_22), .A (n_1537), .B1 (n_1244), .B2 (n_1534));
NAND2_X1 i_36 (.ZN (n_21), .A1 (n_1238), .A2 (n_1594));
XOR2_X1 i_35 (.Z (n_20), .A (n_21), .B (n_22));
INV_X1 i_34 (.ZN (Res_imm[14]), .A (n_20));
NAND2_X1 i_33 (.ZN (n_19), .A1 (n_1537), .A2 (n_1535));
XNOR2_X1 i_32 (.ZN (n_18), .A (n_1244), .B (n_19));
INV_X1 i_31 (.ZN (Res_imm[13]), .A (n_18));
NAND2_X1 i_30 (.ZN (n_17), .A1 (n_1530), .A2 (n_1488));
NAND2_X1 i_29 (.ZN (n_16), .A1 (n_1491), .A2 (n_17));
AOI21_X1 i_28 (.ZN (n_15), .A (n_1246), .B1 (n_1248), .B2 (n_1449));
XOR2_X1 i_27 (.Z (n_14), .A (n_16), .B (n_15));
INV_X1 i_26 (.ZN (Res_imm[12]), .A (n_14));
INV_X1 i_25 (.ZN (n_13), .A (n_1246));
NAND2_X1 i_24 (.ZN (n_12), .A1 (n_13), .A2 (n_1449));
XOR2_X1 i_23 (.Z (Res_imm[11]), .A (n_1248), .B (n_12));
NAND2_X1 i_22 (.ZN (n_11), .A1 (n_1339), .A2 (n_1334));
XNOR2_X1 i_21 (.ZN (Res_imm[10]), .A (n_11), .B (n_1249));
NAND2_X1 i_20 (.ZN (n_10), .A1 (n_1324), .A2 (n_1328));
XOR2_X1 i_19 (.Z (Res_imm[9]), .A (n_1250), .B (n_10));
NAND2_X1 i_18 (.ZN (n_9), .A1 (n_1315), .A2 (n_1314));
XNOR2_X1 i_17 (.ZN (Res_imm[8]), .A (n_9), .B (n_1251));
NAND2_X1 i_16 (.ZN (n_8), .A1 (n_1306), .A2 (n_1253));
XOR2_X1 i_15 (.Z (Res_imm[7]), .A (n_8), .B (n_1256));
NAND2_X1 i_14 (.ZN (n_7), .A1 (n_1297), .A2 (n_1296));
XOR2_X1 i_13 (.Z (Res_imm[6]), .A (n_1258), .B (n_7));
NAND2_X1 i_12 (.ZN (n_6), .A1 (n_1288), .A2 (n_1287));
XOR2_X1 i_11 (.Z (Res_imm[5]), .A (n_1260), .B (n_6));
NAND2_X1 i_10 (.ZN (n_5), .A1 (n_1281), .A2 (n_1280));
XOR2_X1 i_9 (.Z (Res_imm[4]), .A (n_1262), .B (n_5));
NAND2_X1 i_8 (.ZN (n_4), .A1 (n_1273), .A2 (n_1272));
XOR2_X1 i_7 (.Z (Res_imm[3]), .A (n_1264), .B (n_4));
NAND2_X1 i_6 (.ZN (n_3), .A1 (n_1270), .A2 (n_1268));
XNOR2_X1 i_5 (.ZN (Res_imm[2]), .A (n_3), .B (n_1265));
OAI22_X1 i_4 (.ZN (n_2), .A1 (n_6740), .A2 (n_6836), .B1 (n_4366), .B2 (n_3554));
NAND2_X1 i_3 (.ZN (n_1), .A1 (n_2), .A2 (n_1271));
INV_X1 i_2 (.ZN (Res_imm[1]), .A (n_1));
NAND2_X1 i_1 (.ZN (n_0), .A1 (A_imm[0]), .A2 (B_imm[0]));
INV_X1 i_0 (.ZN (Res_imm[0]), .A (n_0));
INV_X1 sgo__sro_c243 (.ZN (sgo__sro_n130), .A (n_144));
INV_X1 sgo__sro_c244 (.ZN (sgo__sro_n129), .A (n_971));
NAND2_X1 sgo__sro_c245 (.ZN (sgo__sro_n128), .A1 (sgo__sro_n130), .A2 (sgo__sro_n129));
OAI21_X1 sgo__sro_c246 (.ZN (n_131), .A (sgo__sro_n128), .B1 (n_132), .B2 (n_972));
INV_X1 sgo__sro_c301 (.ZN (sgo__sro_n157), .A (n_6817));
NAND2_X1 sgo__sro_c302 (.ZN (sgo__sro_n156), .A1 (sgo__sro_n158), .A2 (sgo__sro_n157));
INV_X1 sgo__sro_c156 (.ZN (sgo__sro_n83), .A (n_1038));
INV_X1 sgo__sro_c157 (.ZN (sgo__sro_n82), .A (n_1020));
NOR2_X1 sgo__sro_c158 (.ZN (sgo__sro_n81), .A1 (sgo__sro_n83), .A2 (sgo__sro_n82));
NAND3_X1 sgo__sro_c159 (.ZN (n_1007), .A1 (n_1008), .A2 (n_1010), .A3 (sgo__sro_n81));
INV_X2 CLOCK_opt_ipo_c546 (.ZN (CLOCK_opt_ipo_n324), .A (n_997));
INV_X2 CLOCK_opt_ipo_c548 (.ZN (CLOCK_opt_ipo_n326), .A (n_999));
INV_X4 CLOCK_opt_ipo_c555 (.ZN (CLOCK_opt_ipo_n333), .A (n_2630));
AND2_X2 sgo__c284 (.ZN (n_4221), .A1 (n_4222), .A2 (n_4229));
INV_X1 CLOCK_opt_ipo_c565 (.ZN (CLOCK_opt_ipo_n345), .A (n_238));
INV_X4 CLOCK_opt_ipo_c571 (.ZN (CLOCK_opt_ipo_n351), .A (n_5657));
INV_X2 CLOCK_opt_ipo_c579 (.ZN (Res_imm[41]), .A (CLOCK_opt_ipo_n363));
AND4_X4 sgo__c412 (.ZN (n_5109), .A1 (CLOCK_opt_ipo_n528), .A2 (CLOCK_opt_ipo_n351)
    , .A3 (n_6934), .A4 (n_5724));
INV_X4 CLOCK_opt_ipo_c634 (.ZN (CLOCK_opt_ipo_n418), .A (n_1136));
INV_X1 CLOCK_opt_ipo_c639 (.ZN (CLOCK_opt_ipo_n423), .A (n_2327));
BUF_X4 CLOCK_opt_ipo_c641 (.Z (CLOCK_opt_ipo_n425), .A (n_2105));
BUF_X4 CLOCK_opt_ipo_c649 (.Z (CLOCK_opt_ipo_n433), .A (n_9003));
INV_X4 CLOCK_opt_ipo_c666 (.ZN (Res_imm[57]), .A (CLOCK_opt_ipo_n452));
INV_X2 CLOCK_opt_ipo_c742 (.ZN (CLOCK_opt_ipo_n528), .A (n_5111));

endmodule //datapath__0_2

module datapath__0_0 (opt_ipoPP_0, A_in, p_0);

output [31:0] p_0;
input [31:0] A_in;
input opt_ipoPP_0;
wire n_6;
wire n_96;
wire n_15;
wire n_19;
wire n_0;
wire n_3;
wire n_2;
wire n_1;
wire n_12;
wire n_16;
wire n_11;
wire n_14;
wire n_7;
wire n_23;
wire n_8;
wire n_18;
wire n_13;
wire n_17;
wire n_32;
wire n_28;
wire n_52;
wire n_57;
wire n_54;
wire n_59;
wire n_65;
wire n_47;
wire n_48;
wire n_46;
wire n_66;
wire n_62;
wire n_51;
wire n_63;
wire n_69;
wire n_4;
wire n_5;
wire n_9;
wire n_10;
wire n_20;
wire n_22;
wire n_21;
wire n_24;
wire n_25;
wire n_27;
wire n_30;
wire n_31;
wire n_29;
wire n_33;
wire n_37;
wire n_34;
wire n_35;
wire n_36;
wire n_38;
wire n_40;
wire n_39;
wire n_42;
wire n_41;
wire n_43;
wire n_44;
wire n_45;
wire n_50;
wire n_49;
wire n_53;
wire n_55;
wire n_56;
wire n_58;
wire n_60;
wire n_61;
wire n_64;
wire n_67;
wire n_70;
wire n_68;
wire n_71;
wire n_72;
wire n_73;
wire n_75;
wire n_76;
wire n_78;
wire n_77;
wire n_80;
wire n_79;
wire n_82;
wire n_81;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_97;
wire CLOCK_opt_ipo_n46;
wire CLOCK_opt_ipo_n82;


NAND3_X1 i_128 (.ZN (n_97), .A1 (n_54), .A2 (n_88), .A3 (n_79));
NOR4_X2 i_127 (.ZN (n_96), .A1 (A_in[30]), .A2 (A_in[29]), .A3 (A_in[28]), .A4 (n_97));
AOI21_X1 i_126 (.ZN (p_0[30]), .A (n_96), .B1 (A_in[30]), .B2 (n_94));
INV_X1 i_125 (.ZN (n_95), .A (A_in[29]));
NAND4_X1 i_124 (.ZN (n_94), .A1 (n_95), .A2 (n_70), .A3 (n_92), .A4 (n_88));
INV_X1 i_123 (.ZN (n_93), .A (n_94));
AOI21_X1 i_122 (.ZN (p_0[29]), .A (n_93), .B1 (n_90), .B2 (A_in[29]));
INV_X1 i_121 (.ZN (n_92), .A (A_in[28]));
NAND3_X1 i_119 (.ZN (n_90), .A1 (n_92), .A2 (n_70), .A3 (n_88));
OAI21_X1 i_118 (.ZN (n_89), .A (n_90), .B1 (n_92), .B2 (n_85));
INV_X1 i_117 (.ZN (p_0[28]), .A (n_89));
INV_X1 i_116 (.ZN (n_88), .A (n_87));
NAND2_X1 i_115 (.ZN (n_87), .A1 (n_86), .A2 (n_82));
INV_X1 i_114 (.ZN (n_86), .A (A_in[27]));
AOI21_X1 i_113 (.ZN (p_0[27]), .A (n_85), .B1 (A_in[27]), .B2 (n_84));
NOR2_X1 i_112 (.ZN (n_85), .A1 (n_84), .A2 (A_in[27]));
NAND2_X1 i_111 (.ZN (n_84), .A1 (n_70), .A2 (n_82));
INV_X1 i_110 (.ZN (n_83), .A (n_78));
NOR2_X1 i_109 (.ZN (n_82), .A1 (n_83), .A2 (A_in[26]));
NAND3_X1 i_108 (.ZN (n_81), .A1 (n_78), .A2 (n_79), .A3 (n_54));
AOI22_X1 i_107 (.ZN (p_0[26]), .A1 (n_70), .A2 (n_82), .B1 (A_in[26]), .B2 (n_81));
INV_X1 i_106 (.ZN (n_80), .A (A_in[24]));
INV_X1 i_105 (.ZN (n_79), .A (n_71));
NOR2_X1 i_104 (.ZN (n_78), .A1 (A_in[25]), .A2 (A_in[24]));
NAND3_X1 i_103 (.ZN (n_77), .A1 (n_80), .A2 (n_54), .A3 (n_79));
AOI22_X1 i_102 (.ZN (p_0[25]), .A1 (n_70), .A2 (n_78), .B1 (A_in[25]), .B2 (n_77));
INV_X1 i_101 (.ZN (n_76), .A (n_70));
NOR3_X1 i_100 (.ZN (n_75), .A1 (A_in[24]), .A2 (n_71), .A3 (n_46));
AOI21_X1 i_99 (.ZN (p_0[24]), .A (n_75), .B1 (n_76), .B2 (A_in[24]));
NOR3_X1 i_97 (.ZN (n_73), .A1 (A_in[21]), .A2 (A_in[20]), .A3 (A_in[22]));
NOR2_X1 i_96 (.ZN (n_72), .A1 (A_in[23]), .A2 (n_56));
NAND4_X2 i_95 (.ZN (n_71), .A1 (n_67), .A2 (n_60), .A3 (n_72), .A4 (n_73));
NOR2_X2 i_94 (.ZN (n_70), .A1 (n_46), .A2 (n_71));
NOR4_X1 i_93 (.ZN (n_69), .A1 (A_in[22]), .A2 (A_in[21]), .A3 (A_in[20]), .A4 (n_66));
NAND2_X1 i_92 (.ZN (n_68), .A1 (n_54), .A2 (CLOCK_opt_ipo_n82));
AOI21_X1 i_91 (.ZN (p_0[23]), .A (n_70), .B1 (A_in[23]), .B2 (n_68));
INV_X1 i_90 (.ZN (n_67), .A (A_in[19]));
NAND2_X1 i_89 (.ZN (n_66), .A1 (n_67), .A2 (n_58));
INV_X1 i_88 (.ZN (n_65), .A (n_66));
NOR2_X1 i_87 (.ZN (n_64), .A1 (A_in[21]), .A2 (A_in[20]));
NAND4_X2 i_86 (.ZN (n_63), .A1 (n_33), .A2 (n_64), .A3 (n_65), .A4 (n_49));
INV_X1 i_85 (.ZN (n_62), .A (n_63));
AND2_X1 i_84 (.ZN (p_0[18]), .A1 (n_59), .A2 (n_61));
OAI21_X1 i_83 (.ZN (n_61), .A (A_in[18]), .B1 (n_56), .B2 (n_46));
INV_X1 i_82 (.ZN (n_60), .A (A_in[18]));
NAND2_X1 i_81 (.ZN (n_59), .A1 (n_58), .A2 (n_54));
NOR2_X1 i_80 (.ZN (n_58), .A1 (n_56), .A2 (A_in[18]));
INV_X1 i_79 (.ZN (n_57), .A (n_56));
NAND2_X2 i_78 (.ZN (n_56), .A1 (n_55), .A2 (n_53));
INV_X1 i_77 (.ZN (n_55), .A (A_in[17]));
INV_X4 i_76 (.ZN (n_54), .A (n_46));
INV_X2 i_75 (.ZN (n_53), .A (A_in[16]));
NAND2_X1 i_74 (.ZN (n_52), .A1 (n_54), .A2 (n_53));
AOI22_X1 i_73 (.ZN (p_0[16]), .A1 (n_54), .A2 (n_53), .B1 (n_46), .B2 (A_in[16]));
INV_X1 i_72 (.ZN (n_50), .A (A_in[15]));
AND4_X4 i_71 (.ZN (n_49), .A1 (n_50), .A2 (n_44), .A3 (n_41), .A4 (n_42));
NAND4_X4 i_70 (.ZN (n_46), .A1 (n_8), .A2 (n_49), .A3 (n_23), .A4 (n_36));
OAI21_X1 i_69 (.ZN (n_45), .A (n_46), .B1 (n_50), .B2 (n_43));
INV_X1 i_68 (.ZN (p_0[15]), .A (n_45));
INV_X1 i_66 (.ZN (n_44), .A (A_in[14]));
AND4_X1 i_65 (.ZN (n_43), .A1 (n_42), .A2 (n_41), .A3 (n_44), .A4 (n_33));
AOI21_X1 i_64 (.ZN (p_0[14]), .A (n_43), .B1 (A_in[14]), .B2 (n_40));
INV_X1 i_63 (.ZN (n_42), .A (A_in[13]));
INV_X1 i_62 (.ZN (n_41), .A (A_in[12]));
NAND3_X1 i_61 (.ZN (n_40), .A1 (n_42), .A2 (n_33), .A3 (n_41));
OAI21_X1 i_60 (.ZN (n_39), .A (A_in[13]), .B1 (A_in[12]), .B2 (n_34));
AND2_X1 i_59 (.ZN (p_0[13]), .A1 (n_40), .A2 (n_39));
XOR2_X1 i_58 (.Z (p_0[12]), .A (n_34), .B (A_in[12]));
INV_X1 i_57 (.ZN (n_38), .A (A_in[11]));
INV_X1 i_56 (.ZN (n_37), .A (A_in[10]));
AND4_X4 i_55 (.ZN (n_36), .A1 (n_38), .A2 (A_in[8]), .A3 (n_37), .A4 (n_31));
NOR2_X1 i_54 (.ZN (n_35), .A1 (A_in[3]), .A2 (A_in[0]));
NAND4_X2 i_53 (.ZN (n_34), .A1 (n_10), .A2 (n_23), .A3 (n_35), .A4 (n_36));
INV_X2 i_52 (.ZN (n_33), .A (n_34));
NAND4_X1 i_51 (.ZN (n_32), .A1 (n_37), .A2 (n_29), .A3 (n_31), .A4 (CLOCK_opt_ipo_n46));
AOI21_X1 i_50 (.ZN (p_0[11]), .A (n_33), .B1 (A_in[11]), .B2 (n_32));
INV_X2 i_49 (.ZN (n_31), .A (A_in[9]));
NAND2_X1 i_48 (.ZN (n_30), .A1 (n_8), .A2 (n_23));
INV_X1 i_47 (.ZN (n_29), .A (n_30));
NAND3_X1 i_46 (.ZN (n_28), .A1 (n_31), .A2 (n_29), .A3 (CLOCK_opt_ipo_n46));
OAI21_X1 i_45 (.ZN (n_27), .A (A_in[9]), .B1 (opt_ipoPP_0), .B2 (n_30));
AND2_X1 i_44 (.ZN (p_0[9]), .A1 (n_28), .A2 (n_27));
INV_X1 i_42 (.ZN (n_25), .A (A_in[7]));
NAND4_X4 i_41 (.ZN (n_24), .A1 (n_25), .A2 (n_20), .A3 (n_16), .A4 (n_19));
INV_X4 i_40 (.ZN (n_23), .A (n_24));
OR2_X1 i_39 (.ZN (n_22), .A1 (n_9), .A2 (n_24));
NOR2_X1 i_38 (.ZN (n_21), .A1 (opt_ipoPP_0), .A2 (n_24));
AOI22_X1 i_37 (.ZN (p_0[8]), .A1 (opt_ipoPP_0), .A2 (n_22), .B1 (n_8), .B2 (n_21));
INV_X2 i_36 (.ZN (n_20), .A (A_in[6]));
INV_X2 i_35 (.ZN (n_19), .A (A_in[5]));
AND3_X1 i_34 (.ZN (n_18), .A1 (n_19), .A2 (n_16), .A3 (n_20));
INV_X4 i_33 (.ZN (n_16), .A (A_in[4]));
NAND2_X1 i_32 (.ZN (n_15), .A1 (n_16), .A2 (n_8));
AOI22_X1 i_31 (.ZN (p_0[4]), .A1 (n_16), .A2 (n_8), .B1 (A_in[4]), .B2 (n_9));
INV_X2 i_30 (.ZN (n_14), .A (A_in[3]));
INV_X4 i_29 (.ZN (n_12), .A (A_in[1]));
INV_X4 i_28 (.ZN (n_11), .A (A_in[0]));
AND2_X4 i_27 (.ZN (n_10), .A1 (n_12), .A2 (n_7));
NAND3_X4 i_26 (.ZN (n_9), .A1 (n_14), .A2 (n_11), .A3 (n_10));
INV_X4 i_25 (.ZN (n_8), .A (n_9));
AOI21_X1 i_24 (.ZN (p_0[3]), .A (n_8), .B1 (A_in[3]), .B2 (n_5));
INV_X2 i_23 (.ZN (n_7), .A (A_in[2]));
NOR2_X1 i_22 (.ZN (n_6), .A1 (A_in[1]), .A2 (A_in[0]));
NAND2_X1 i_21 (.ZN (n_5), .A1 (n_7), .A2 (n_6));
OAI21_X1 i_20 (.ZN (n_4), .A (n_5), .B1 (n_7), .B2 (n_6));
INV_X1 i_19 (.ZN (p_0[2]), .A (n_4));
AOI22_X1 i_18 (.ZN (p_0[22]), .A1 (n_63), .A2 (A_in[22]), .B1 (CLOCK_opt_ipo_n82), .B2 (n_54));
INV_X1 i_17 (.ZN (n_51), .A (A_in[20]));
NAND3_X1 i_16 (.ZN (n_48), .A1 (n_54), .A2 (n_51), .A3 (n_65));
AOI21_X1 i_15 (.ZN (p_0[21]), .A (n_62), .B1 (n_48), .B2 (A_in[21]));
OAI21_X1 i_14 (.ZN (n_47), .A (A_in[20]), .B1 (n_46), .B2 (n_66));
AND2_X1 i_13 (.ZN (p_0[20]), .A1 (n_47), .A2 (n_48));
AOI22_X1 i_12 (.ZN (p_0[19]), .A1 (n_59), .A2 (A_in[19]), .B1 (n_65), .B2 (n_54));
AOI22_X1 i_11 (.ZN (p_0[17]), .A1 (n_52), .A2 (A_in[17]), .B1 (n_57), .B2 (n_54));
NAND2_X1 i_10 (.ZN (n_17), .A1 (n_28), .A2 (A_in[10]));
NAND2_X1 i_9 (.ZN (n_13), .A1 (n_17), .A2 (n_32));
INV_X1 i_8 (.ZN (p_0[10]), .A (n_13));
NAND2_X1 i_7 (.ZN (n_3), .A1 (n_8), .A2 (n_18));
AOI22_X1 i_6 (.ZN (p_0[7]), .A1 (A_in[7]), .A2 (n_3), .B1 (n_23), .B2 (n_8));
NAND3_X1 i_5 (.ZN (n_2), .A1 (n_11), .A2 (n_14), .A3 (n_7));
NAND3_X1 i_4 (.ZN (n_1), .A1 (n_12), .A2 (n_16), .A3 (n_19));
OAI21_X1 i_3 (.ZN (n_0), .A (A_in[6]), .B1 (n_2), .B2 (n_1));
AND2_X1 i_2 (.ZN (p_0[6]), .A1 (n_0), .A2 (n_3));
XNOR2_X1 i_1 (.ZN (p_0[5]), .A (n_15), .B (n_19));
XNOR2_X1 i_67 (.ZN (p_0[31]), .A (A_in[31]), .B (n_96));
AOI21_X1 i_0 (.ZN (p_0[1]), .A (n_6), .B1 (A_in[1]), .B2 (A_in[0]));
INV_X1 CLOCK_opt_ipo_c70 (.ZN (CLOCK_opt_ipo_n46), .A (opt_ipoPP_0));
BUF_X1 CLOCK_opt_ipo_c93 (.Z (CLOCK_opt_ipo_n82), .A (n_69));

endmodule //datapath__0_0

module datapath (opt_ipoPP_0, opt_ipoPP_2, B_in, p_0);

output [31:0] p_0;
input [31:0] B_in;
input opt_ipoPP_0;
input opt_ipoPP_2;
wire n_36;
wire n_17;
wire n_1;
wire n_8;
wire n_38;
wire n_0;
wire n_10;
wire n_7;
wire n_15;
wire n_6;
wire n_13;
wire n_34;
wire n_55;
wire n_50;
wire n_89;
wire n_85;
wire n_14;
wire n_29;
wire n_41;
wire n_24;
wire n_2;
wire n_5;
wire n_19;
wire n_9;
wire n_20;
wire n_22;
wire n_23;
wire n_21;
wire n_31;
wire n_30;
wire n_90;
wire n_93;
wire n_57;
wire n_46;
wire n_56;
wire n_54;
wire n_47;
wire n_64;
wire n_67;
wire n_62;
wire n_51;
wire n_81;
wire n_102;
wire n_88;
wire n_84;
wire n_92;
wire n_3;
wire n_4;
wire n_11;
wire n_18;
wire n_16;
wire n_25;
wire n_27;
wire n_26;
wire n_28;
wire n_32;
wire n_33;
wire n_35;
wire n_39;
wire n_40;
wire n_45;
wire n_42;
wire n_43;
wire n_44;
wire n_48;
wire n_49;
wire n_52;
wire n_53;
wire n_58;
wire n_60;
wire n_59;
wire n_65;
wire n_61;
wire n_63;
wire n_66;
wire sgo__n20;
wire n_69;
wire n_70;
wire n_72;
wire n_71;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_82;
wire n_83;
wire n_87;
wire n_91;
wire n_94;
wire n_96;
wire n_95;
wire n_98;
wire n_97;
wire n_99;
wire n_101;
wire n_100;
wire n_104;
wire n_103;
wire n_105;
wire sgo__n14;
wire sgo__sro_n28;
wire CLOCK_opt_ipo_n65;
wire CLOCK_opt_ipo_n66;


NAND2_X1 i_136 (.ZN (n_105), .A1 (n_102), .A2 (n_104));
XOR2_X1 i_135 (.Z (p_0[31]), .A (B_in[31]), .B (n_105));
NOR2_X1 i_134 (.ZN (n_104), .A1 (n_100), .A2 (B_in[30]));
NAND3_X1 i_133 (.ZN (n_103), .A1 (CLOCK_opt_ipo_n66), .A2 (n_97), .A3 (n_101));
AOI22_X1 i_132 (.ZN (p_0[30]), .A1 (n_102), .A2 (n_104), .B1 (B_in[30]), .B2 (n_103));
INV_X1 i_131 (.ZN (n_102), .A (n_96));
NOR2_X1 i_130 (.ZN (n_101), .A1 (B_in[29]), .A2 (B_in[28]));
INV_X1 i_129 (.ZN (n_100), .A (n_101));
NAND4_X1 i_128 (.ZN (n_99), .A1 (n_51), .A2 (n_38), .A3 (n_84), .A4 (n_95));
AOI22_X1 i_127 (.ZN (p_0[29]), .A1 (B_in[29]), .A2 (n_99), .B1 (n_102), .B2 (n_101));
INV_X1 i_126 (.ZN (n_98), .A (n_92));
NOR2_X1 i_125 (.ZN (n_97), .A1 (B_in[27]), .A2 (n_98));
NAND4_X1 i_124 (.ZN (n_96), .A1 (n_51), .A2 (n_38), .A3 (n_84), .A4 (n_97));
NOR3_X1 i_123 (.ZN (n_95), .A1 (B_in[28]), .A2 (n_98), .A3 (B_in[27]));
AOI22_X1 i_122 (.ZN (p_0[28]), .A1 (B_in[28]), .A2 (n_96), .B1 (CLOCK_opt_ipo_n66), .B2 (n_95));
NOR2_X1 i_121 (.ZN (n_94), .A1 (B_in[25]), .A2 (B_in[24]));
NAND4_X1 i_120 (.ZN (n_93), .A1 (n_51), .A2 (n_38), .A3 (n_94), .A4 (n_84));
NOR3_X1 i_119 (.ZN (n_92), .A1 (B_in[26]), .A2 (B_in[25]), .A3 (B_in[24]));
AOI22_X1 i_118 (.ZN (p_0[26]), .A1 (B_in[26]), .A2 (n_93), .B1 (CLOCK_opt_ipo_n66), .B2 (n_92));
NOR2_X1 i_117 (.ZN (n_91), .A1 (n_6), .A2 (B_in[24]));
NAND3_X1 i_116 (.ZN (n_90), .A1 (n_51), .A2 (n_84), .A3 (n_91));
INV_X1 i_115 (.ZN (n_89), .A (n_90));
AOI21_X1 i_114 (.ZN (p_0[23]), .A (CLOCK_opt_ipo_n66), .B1 (B_in[23]), .B2 (n_87));
NAND4_X1 i_113 (.ZN (n_87), .A1 (n_51), .A2 (n_38), .A3 (n_82), .A4 (n_71));
NAND3_X1 i_111 (.ZN (n_85), .A1 (n_84), .A2 (n_51), .A3 (n_38));
AND4_X1 i_110 (.ZN (n_84), .A1 (n_83), .A2 (n_66), .A3 (n_72), .A4 (n_82));
INV_X1 i_109 (.ZN (n_83), .A (B_in[23]));
NOR3_X4 i_108 (.ZN (n_82), .A1 (B_in[21]), .A2 (B_in[20]), .A3 (B_in[22]));
AOI22_X1 i_107 (.ZN (p_0[22]), .A1 (n_76), .A2 (n_82), .B1 (B_in[22]), .B2 (n_79));
NAND2_X1 i_106 (.ZN (n_81), .A1 (n_79), .A2 (n_80));
NAND2_X1 i_105 (.ZN (n_80), .A1 (n_75), .A2 (B_in[21]));
NAND4_X1 i_104 (.ZN (n_79), .A1 (n_78), .A2 (n_51), .A3 (n_38), .A4 (n_71));
NOR2_X1 i_103 (.ZN (n_78), .A1 (B_in[20]), .A2 (B_in[21]));
AOI21_X1 i_102 (.ZN (p_0[20]), .A (n_77), .B1 (B_in[20]), .B2 (n_70));
INV_X1 i_101 (.ZN (n_77), .A (n_75));
INV_X1 i_100 (.ZN (n_76), .A (n_70));
NAND4_X1 i_99 (.ZN (n_75), .A1 (n_74), .A2 (n_72), .A3 (n_51), .A4 (n_38));
NOR2_X1 i_98 (.ZN (n_74), .A1 (n_73), .A2 (B_in[20]));
INV_X1 i_97 (.ZN (n_73), .A (n_66));
INV_X1 i_96 (.ZN (n_72), .A (B_in[19]));
AND2_X1 i_95 (.ZN (n_71), .A1 (n_72), .A2 (n_66));
NAND3_X1 i_94 (.ZN (n_70), .A1 (n_51), .A2 (n_38), .A3 (n_71));
OAI21_X1 i_93 (.ZN (n_69), .A (n_70), .B1 (n_72), .B2 (n_65));
INV_X1 i_92 (.ZN (p_0[19]), .A (n_69));
OR2_X4 sgo__c30 (.ZN (sgo__n20), .A1 (n_40), .A2 (n_10));
INV_X2 i_90 (.ZN (n_67), .A (n_58));
NOR3_X2 i_89 (.ZN (n_66), .A1 (B_in[17]), .A2 (B_in[16]), .A3 (B_in[18]));
AND3_X1 i_88 (.ZN (n_65), .A1 (n_51), .A2 (n_66), .A3 (n_38));
NAND2_X1 i_87 (.ZN (n_63), .A1 (n_35), .A2 (n_53));
NOR2_X1 i_86 (.ZN (n_62), .A1 (B_in[17]), .A2 (n_63));
NAND2_X1 i_85 (.ZN (n_61), .A1 (n_67), .A2 (n_62));
AOI21_X1 i_84 (.ZN (p_0[18]), .A (n_65), .B1 (B_in[18]), .B2 (n_61));
INV_X1 i_83 (.ZN (n_60), .A (B_in[16]));
AND2_X4 sgo__sro_c45 (.ZN (sgo__sro_n28), .A1 (n_5), .A2 (n_11));
NAND4_X1 i_81 (.ZN (n_58), .A1 (n_60), .A2 (n_27), .A3 (n_11), .A4 (n_59));
NOR2_X1 i_80 (.ZN (n_55), .A1 (n_52), .A2 (n_58));
INV_X1 i_79 (.ZN (n_54), .A (B_in[15]));
AND4_X1 i_78 (.ZN (n_53), .A1 (n_54), .A2 (n_49), .A3 (n_44), .A4 (n_43));
NAND2_X2 i_77 (.ZN (n_52), .A1 (n_35), .A2 (n_53));
INV_X4 i_76 (.ZN (n_51), .A (n_52));
NAND2_X2 i_75 (.ZN (n_50), .A1 (n_38), .A2 (n_51));
INV_X1 i_74 (.ZN (n_49), .A (B_in[14]));
AND2_X1 i_73 (.ZN (n_48), .A1 (n_49), .A2 (n_44));
NAND4_X1 i_72 (.ZN (n_47), .A1 (n_43), .A2 (n_38), .A3 (n_35), .A4 (n_48));
NAND2_X1 i_71 (.ZN (n_46), .A1 (n_45), .A2 (n_42));
INV_X1 i_70 (.ZN (n_45), .A (n_34));
INV_X1 i_69 (.ZN (n_44), .A (B_in[13]));
INV_X1 i_68 (.ZN (n_43), .A (B_in[12]));
NOR2_X1 i_67 (.ZN (n_42), .A1 (B_in[13]), .A2 (B_in[12]));
NAND3_X1 i_66 (.ZN (n_41), .A1 (n_38), .A2 (n_35), .A3 (n_43));
AOI22_X1 i_65 (.ZN (p_0[13]), .A1 (B_in[13]), .A2 (n_41), .B1 (n_45), .B2 (n_42));
INV_X2 i_64 (.ZN (n_40), .A (n_27));
INV_X1 i_63 (.ZN (n_39), .A (B_in[11]));
INV_X8 sgo__c32 (.ZN (n_38), .A (sgo__n20));
AND4_X2 i_60 (.ZN (n_35), .A1 (n_39), .A2 (n_33), .A3 (n_32), .A4 (n_31));
NAND2_X1 i_59 (.ZN (n_34), .A1 (n_38), .A2 (n_35));
AOI22_X1 i_58 (.ZN (p_0[11]), .A1 (n_38), .A2 (n_35), .B1 (B_in[11]), .B2 (n_16));
INV_X1 i_57 (.ZN (n_33), .A (B_in[10]));
INV_X1 i_56 (.ZN (n_32), .A (B_in[9]));
INV_X1 i_55 (.ZN (n_31), .A (B_in[8]));
INV_X1 i_54 (.ZN (n_29), .A (B_in[6]));
NAND2_X4 i_53 (.ZN (n_28), .A1 (n_14), .A2 (B_in[4]));
NOR3_X4 i_52 (.ZN (n_27), .A1 (B_in[7]), .A2 (B_in[6]), .A3 (n_28));
NAND3_X1 i_51 (.ZN (n_26), .A1 (n_11), .A2 (n_4), .A3 (n_5));
NOR3_X1 i_50 (.ZN (n_25), .A1 (B_in[9]), .A2 (n_26), .A3 (B_in[8]));
NAND3_X1 i_49 (.ZN (n_21), .A1 (n_3), .A2 (n_25), .A3 (n_27));
NOR2_X2 i_48 (.ZN (n_18), .A1 (B_in[10]), .A2 (n_21));
INV_X1 i_47 (.ZN (n_16), .A (n_18));
AOI21_X1 i_46 (.ZN (p_0[10]), .A (n_18), .B1 (B_in[10]), .B2 (n_21));
INV_X4 i_45 (.ZN (n_14), .A (B_in[5]));
INV_X2 i_43 (.ZN (n_11), .A (B_in[3]));
OR2_X1 i_41 (.ZN (n_9), .A1 (opt_ipoPP_0), .A2 (n_10));
OR2_X1 i_40 (.ZN (n_8), .A1 (B_in[5]), .A2 (n_9));
INV_X2 i_39 (.ZN (n_5), .A (B_in[2]));
XNOR2_X1 i_38 (.ZN (p_0[2]), .A (B_in[2]), .B (n_2));
INV_X2 i_37 (.ZN (n_4), .A (B_in[1]));
INV_X2 i_36 (.ZN (n_3), .A (B_in[0]));
NOR2_X2 i_35 (.ZN (n_2), .A1 (B_in[1]), .A2 (B_in[0]));
AOI21_X1 i_34 (.ZN (p_0[1]), .A (n_2), .B1 (B_in[1]), .B2 (B_in[0]));
NAND4_X1 i_33 (.ZN (n_88), .A1 (n_51), .A2 (n_38), .A3 (n_84), .A4 (n_92));
AOI21_X1 i_32 (.ZN (p_0[27]), .A (n_102), .B1 (n_88), .B2 (B_in[27]));
INV_X1 i_31 (.ZN (p_0[21]), .A (n_81));
NAND2_X1 i_30 (.ZN (n_64), .A1 (n_67), .A2 (n_51));
AOI22_X1 i_29 (.ZN (p_0[17]), .A1 (n_64), .A2 (B_in[17]), .B1 (n_67), .B2 (n_62));
INV_X1 i_28 (.ZN (n_57), .A (n_47));
OAI21_X1 i_27 (.ZN (n_56), .A (n_50), .B1 (n_57), .B2 (n_54));
INV_X1 i_26 (.ZN (p_0[15]), .A (n_56));
AOI21_X1 i_25 (.ZN (p_0[14]), .A (n_57), .B1 (B_in[14]), .B2 (n_46));
INV_X1 i_24 (.ZN (n_36), .A (n_10));
INV_X1 i_22 (.ZN (n_30), .A (n_93));
AOI21_X1 i_21 (.ZN (p_0[25]), .A (n_30), .B1 (n_90), .B2 (B_in[25]));
NAND2_X1 i_20 (.ZN (n_24), .A1 (n_38), .A2 (n_31));
NAND2_X1 i_19 (.ZN (n_23), .A1 (n_24), .A2 (B_in[9]));
NAND2_X1 i_18 (.ZN (n_22), .A1 (n_23), .A2 (n_21));
INV_X1 i_17 (.ZN (p_0[9]), .A (n_22));
XNOR2_X1 i_16 (.ZN (p_0[5]), .A (n_9), .B (n_14));
NAND2_X1 i_15 (.ZN (n_20), .A1 (n_10), .A2 (opt_ipoPP_0));
NAND2_X1 i_14 (.ZN (n_19), .A1 (n_9), .A2 (n_20));
INV_X1 i_13 (.ZN (p_0[4]), .A (n_19));
NAND2_X1 i_12 (.ZN (n_17), .A1 (n_2), .A2 (n_5));
INV_X1 i_11 (.ZN (n_15), .A (n_24));
INV_X1 i_23 (.ZN (n_13), .A (n_41));
NAND3_X1 i_9 (.ZN (n_7), .A1 (n_14), .A2 (opt_ipoPP_2), .A3 (n_29));
INV_X1 i_8 (.ZN (n_6), .A (n_38));
AOI21_X1 i_7 (.ZN (p_0[24]), .A (n_89), .B1 (B_in[24]), .B2 (CLOCK_opt_ipo_n65));
AOI21_X1 i_6 (.ZN (p_0[16]), .A (n_55), .B1 (B_in[16]), .B2 (n_50));
AOI21_X1 i_10 (.ZN (p_0[12]), .A (n_13), .B1 (B_in[12]), .B2 (n_34));
AOI21_X1 i_5 (.ZN (p_0[8]), .A (n_15), .B1 (B_in[8]), .B2 (n_6));
NOR2_X1 i_4 (.ZN (n_1), .A1 (n_10), .A2 (n_7));
INV_X1 i_3 (.ZN (n_0), .A (n_1));
AOI21_X1 i_2 (.ZN (p_0[7]), .A (n_38), .B1 (B_in[7]), .B2 (n_0));
AOI21_X1 i_1 (.ZN (p_0[6]), .A (n_1), .B1 (B_in[6]), .B2 (n_8));
AOI21_X1 i_0 (.ZN (p_0[3]), .A (n_36), .B1 (B_in[3]), .B2 (n_17));
NAND3_X1 sgo__c17 (.ZN (sgo__n14), .A1 (n_3), .A2 (n_5), .A3 (n_4));
INV_X1 sgo__c19 (.ZN (n_59), .A (sgo__n14));
NAND3_X4 sgo__sro_c46 (.ZN (n_10), .A1 (n_3), .A2 (sgo__sro_n28), .A3 (n_4));
INV_X1 CLOCK_opt_ipo_c81 (.ZN (CLOCK_opt_ipo_n65), .A (CLOCK_opt_ipo_n66));
INV_X4 CLOCK_opt_ipo_c82 (.ZN (CLOCK_opt_ipo_n66), .A (n_85));

endmodule //datapath

module VM (Res, OVF, A, B, clk, reset, enable);

output OVF;
output [63:0] Res;
input [31:0] A;
input [31:0] B;
input clk;
input enable;
input reset;
wire CLOCK_sgo_n781;
wire CLOCK_slh__n1077;
wire CLOCK_slh_n1056;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire \Res_imm[63] ;
wire \Res_imm[62] ;
wire \Res_imm[61] ;
wire \Res_imm[60] ;
wire \Res_imm[59] ;
wire \Res_imm[58] ;
wire \Res_imm[57] ;
wire \Res_imm[56] ;
wire \Res_imm[55] ;
wire \Res_imm[54] ;
wire \Res_imm[53] ;
wire \Res_imm[52] ;
wire \Res_imm[51] ;
wire \Res_imm[50] ;
wire \Res_imm[49] ;
wire \Res_imm[48] ;
wire \Res_imm[47] ;
wire \Res_imm[46] ;
wire \Res_imm[45] ;
wire \Res_imm[44] ;
wire \Res_imm[43] ;
wire \Res_imm[42] ;
wire \Res_imm[41] ;
wire \Res_imm[40] ;
wire \Res_imm[39] ;
wire \Res_imm[38] ;
wire \Res_imm[37] ;
wire \Res_imm[36] ;
wire \Res_imm[35] ;
wire \Res_imm[34] ;
wire \Res_imm[33] ;
wire \Res_imm[32] ;
wire \Res_imm[31] ;
wire \Res_imm[30] ;
wire \Res_imm[29] ;
wire \Res_imm[28] ;
wire \Res_imm[27] ;
wire \Res_imm[26] ;
wire \Res_imm[25] ;
wire \Res_imm[24] ;
wire \Res_imm[23] ;
wire \Res_imm[22] ;
wire \Res_imm[21] ;
wire \Res_imm[20] ;
wire \Res_imm[19] ;
wire \Res_imm[18] ;
wire \Res_imm[17] ;
wire \Res_imm[16] ;
wire \Res_imm[15] ;
wire \Res_imm[14] ;
wire \Res_imm[13] ;
wire \Res_imm[12] ;
wire \Res_imm[11] ;
wire \Res_imm[10] ;
wire \Res_imm[9] ;
wire \Res_imm[8] ;
wire \Res_imm[7] ;
wire \Res_imm[6] ;
wire \Res_imm[5] ;
wire \Res_imm[4] ;
wire \Res_imm[3] ;
wire \Res_imm[2] ;
wire \Res_imm[1] ;
wire \Res_imm[0] ;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire B_in;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_288;
wire A_in;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_169;
wire n_0_170;
wire n_0_171;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_176;
wire n_0_177;
wire n_0_178;
wire n_0_179;
wire n_0_180;
wire n_0_181;
wire n_0_182;
wire n_0_183;
wire n_0_184;
wire n_0_185;
wire n_0_0;
wire n_0_186;
wire sph__n1165;
wire n_0_1_0;
wire sph__n1166;
wire n_0_1_1;
wire n_0_1_2;
wire n_0_190;
wire n_0_1_3;
wire n_0_191;
wire n_0_1_4;
wire n_0_192;
wire n_0_1_5;
wire CLOCK_slh__n1079;
wire n_0_1_6;
wire n_0_194;
wire n_0_1_7;
wire CLOCK_slh__n1078;
wire n_0_1_8;
wire n_0_196;
wire n_0_1_9;
wire n_0_197;
wire n_0_1_10;
wire n_0_198;
wire n_0_1_11;
wire CLOCK_slh__n1105;
wire n_0_1_12;
wire CLOCK_slh__n1107;
wire n_0_1_13;
wire n_0_201;
wire n_0_1_14;
wire n_0_202;
wire n_0_1_15;
wire n_0_203;
wire n_0_1_16;
wire n_0_204;
wire n_0_1_17;
wire n_0_205;
wire n_0_1_18;
wire n_0_206;
wire n_0_1_19;
wire n_0_207;
wire n_0_1_20;
wire n_0_208;
wire n_0_1_21;
wire n_0_209;
wire n_0_1_22;
wire n_0_210;
wire n_0_1_23;
wire n_0_211;
wire n_0_1_24;
wire n_0_212;
wire n_0_1_25;
wire n_0_213;
wire n_0_1_26;
wire n_0_214;
wire n_0_1_27;
wire n_0_215;
wire n_0_1_28;
wire n_0_216;
wire n_0_1_29;
wire n_0_217;
wire n_0_1_30;
wire n_0_218;
wire n_0_1_31;
wire n_0_219;
wire n_0_1_32;
wire n_0_220;
wire n_0_1_33;
wire n_0_221;
wire n_0_1_34;
wire n_0_222;
wire n_0_1_35;
wire n_0_223;
wire n_0_1_36;
wire n_0_224;
wire n_0_1_37;
wire n_0_225;
wire n_0_1_38;
wire n_0_226;
wire n_0_1_39;
wire n_0_227;
wire n_0_1_40;
wire n_0_228;
wire n_0_1_41;
wire n_0_229;
wire n_0_1_42;
wire n_0_230;
wire n_0_1_43;
wire n_0_231;
wire n_0_1_44;
wire n_0_232;
wire n_0_1_45;
wire n_0_233;
wire n_0_1_46;
wire n_0_234;
wire n_0_1_47;
wire n_0_235;
wire n_0_1_48;
wire n_0_236;
wire n_0_1_49;
wire n_0_237;
wire n_0_1_50;
wire n_0_238;
wire n_0_1_51;
wire n_0_239;
wire n_0_1_52;
wire n_0_240;
wire n_0_1_53;
wire n_0_241;
wire n_0_1_54;
wire n_0_242;
wire n_0_1_55;
wire n_0_243;
wire n_0_1_56;
wire n_0_244;
wire n_0_1_57;
wire n_0_245;
wire n_0_1_58;
wire n_0_246;
wire n_0_1_59;
wire n_0_247;
wire n_0_1_60;
wire n_0_248;
wire n_0_1_61;
wire n_0_249;
wire n_0_1_62;
wire n_0_1_63;
wire n_0_1_64;
wire n_0_1_65;
wire n_0_1_66;
wire n_0_1_67;
wire n_0_1_68;
wire n_0_1_69;
wire n_0_1_70;
wire n_0_1_71;
wire n_0_1_72;
wire n_0_1_73;
wire n_0_1_74;
wire n_0_1_75;
wire n_0_1_76;
wire n_0_1_77;
wire n_0_1_78;
wire sgo__n237;
wire n_0_1_80;
wire n_0_1_81;
wire n_0_1_82;
wire sgo__n270;
wire n_0_1_84;
wire n_0_1_85;
wire sgo__n274;
wire CTS_n769;
wire CTS_n770;
wire \A_imm[31] ;
wire \A_imm[30] ;
wire \A_imm[29] ;
wire \A_imm[28] ;
wire \A_imm[27] ;
wire \A_imm[26] ;
wire \A_imm[25] ;
wire \A_imm[24] ;
wire \A_imm[23] ;
wire \A_imm[22] ;
wire \A_imm[21] ;
wire \A_imm[20] ;
wire \A_imm[19] ;
wire \A_imm[18] ;
wire \A_imm[17] ;
wire \A_imm[16] ;
wire \A_imm[15] ;
wire \A_imm[14] ;
wire \A_imm[13] ;
wire \A_imm[12] ;
wire \A_imm[11] ;
wire \A_imm[10] ;
wire \A_imm[9] ;
wire \A_imm[8] ;
wire \A_imm[7] ;
wire \A_imm[6] ;
wire \A_imm[5] ;
wire \A_imm[4] ;
wire \A_imm[3] ;
wire \A_imm[2] ;
wire \A_imm[1] ;
wire \B_imm[31] ;
wire \B_imm[30] ;
wire \B_imm[29] ;
wire \B_imm[28] ;
wire \B_imm[27] ;
wire \B_imm[26] ;
wire \B_imm[25] ;
wire \B_imm[24] ;
wire \B_imm[23] ;
wire \B_imm[22] ;
wire \B_imm[21] ;
wire \B_imm[20] ;
wire \B_imm[19] ;
wire \B_imm[18] ;
wire \B_imm[17] ;
wire \B_imm[16] ;
wire \B_imm[15] ;
wire \B_imm[14] ;
wire \B_imm[13] ;
wire \B_imm[12] ;
wire \B_imm[11] ;
wire \B_imm[10] ;
wire \B_imm[9] ;
wire \B_imm[8] ;
wire \B_imm[7] ;
wire \B_imm[6] ;
wire \B_imm[5] ;
wire \B_imm[4] ;
wire \B_imm[3] ;
wire \B_imm[2] ;
wire \B_imm[1] ;
wire n_0_1_89;
wire n_0_250;
wire n_0_251;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_255;
wire n_0_256;
wire n_0_257;
wire n_0_258;
wire n_0_259;
wire n_0_260;
wire n_0_261;
wire n_0_262;
wire n_0_263;
wire n_0_264;
wire n_0_265;
wire n_0_266;
wire n_0_267;
wire n_0_268;
wire n_0_269;
wire n_0_270;
wire n_0_271;
wire n_0_272;
wire n_0_273;
wire n_0_274;
wire n_0_275;
wire n_0_276;
wire n_0_277;
wire n_0_278;
wire n_0_279;
wire n_0_280;
wire n_0_281;
wire n_0_283;
wire n_0_284;
wire n_0_285;
wire n_0_286;
wire n_0_287;
wire n_0_289;
wire n_0_290;
wire n_0_291;
wire n_0_292;
wire n_0_293;
wire n_0_294;
wire n_0_295;
wire n_0_296;
wire n_0_297;
wire n_0_298;
wire n_0_299;
wire n_0_300;
wire n_0_301;
wire n_0_302;
wire n_0_303;
wire n_0_304;
wire n_0_305;
wire n_0_306;
wire n_0_307;
wire n_0_308;
wire n_0_309;
wire n_0_310;
wire n_0_311;
wire n_0_312;
wire n_0_313;
wire n_0_314;
wire n_0_315;
wire n_0_316;
wire hfn_ipo_n121;
wire uc_0;
wire uc_1;
wire uc_2;
wire drc_ipo_n127;
wire drc_ipo_n128;
wire drc_ipo_n129;
wire drc_ipo_n130;
wire hfn_ipo_n120;
wire CLOCK_slh__n1106;
wire drc_ipo_n132;
wire drc_ipo_n149;
wire drc_ipo_n133;
wire drc_ipo_n131;
wire sgo__n175;
wire drc_ipo_n169;
wire drc_ipo_n168;
wire drc_ipo_n163;
wire drc_ipo_n159;
wire drc_ipo_n135;
wire drc_ipo_n134;
wire sgo__n220;
wire drc_ipo_n171;
wire drc_ipo_n170;
wire drc_ipo_n165;
wire drc_ipo_n164;
wire drc_ipo_n162;
wire drc_ipo_n161;
wire drc_ipo_n160;
wire drc_ipo_n150;
wire drc_ipo_n148;
wire drc_ipo_n144;
wire drc_ipo_n142;
wire drc_ipo_n141;
wire drc_ipo_n140;
wire drc_ipo_n139;
wire drc_ipo_n138;
wire drc_ipo_n136;
wire sgo__n172;
wire drc_ipo_n167;
wire drc_ipo_n166;
wire drc_ipo_n146;
wire drc_ipo_n145;
wire drc_ipo_n143;
wire drc_ipo_n137;
wire sgo__sro_n179;
wire sgo__n219;
wire drc_ipo_n154;
wire drc_ipo_n153;
wire drc_ipo_n152;
wire sgo__sro_n180;
wire drc_ipo_n156;
wire drc_ipo_n155;
wire drc_ipo_n151;
wire drc_ipo_n147;
wire sgo__sro_n181;
wire drc_ipo_n157;
wire sgo__sro_n182;
wire drc_ipo_n158;
wire drc_ipo_n126;
wire hfn_ipo_n125;
wire hfn_ipo_n123;
wire sgo__n238;
wire sgo__n269;
wire sgo__sro_n246;
wire sgo__sro_n247;
wire sgo__sro_n204;
wire sgo__sro_n205;
wire sgo__sro_n206;
wire sgo__sro_n207;
wire sgo__n291;
wire sgo__sro_n248;
wire sgo__n273;
wire sgo__sro_n256;
wire sgo__sro_n257;
wire sgo__sro_n258;
wire sgo__n292;
wire sgo__n307;
wire sgo__n308;
wire opt_ipo_n598;
wire slo__n360;
wire slo__n361;
wire slo__n366;
wire slo__n367;
wire slo__n383;
wire slo__n384;
wire CLOCK_opt_ipo_n651;
wire CLOCK_opt_ipo_n649;
wire CLOCK_slh__n1059;
wire CLOCK_slh__n1087;
wire CLOCK_slh__n1089;
wire CLOCK_slh__n1088;
wire CLOCK_opt_ipo_n661;
wire CLOCK_opt_ipo_n660;
wire CLOCK_opt_ipo_n663;
wire CLOCK_opt_ipo_n662;
wire CLOCK_slh__n1067;
wire CLOCK_opt_ipo_n664;
wire CLOCK_opt_ipo_n667;
wire CLOCK_opt_ipo_n666;
wire CLOCK_slh__n1058;
wire CLOCK_opt_ipo_n668;
wire CLOCK_slh__n1094;
wire CLOCK_slh__n1093;
wire CLOCK_slh__n1095;
wire CLOCK_slh__n1057;
wire CLOCK_opt_ipo_n679;
wire CLOCK_slh__n1099;
wire CLOCK_slh__n1101;
wire CLOCK_slh__n1100;
wire CLOCK_opt_ipo_n697;
wire CLOCK_opt_ipo_n695;
wire CLOCK_opt_ipo_n701;
wire CLOCK_opt_ipo_n699;
wire CLOCK_opt_ipo_n705;
wire CLOCK_opt_ipo_n703;
wire CLOCK_slh__n1068;
wire CLOCK_slh__n1069;
wire CLOCK_opt_ipo_n727;


BUF_X4 hfn_ipo_c121 (.Z (hfn_ipo_n121), .A (n_0_1_63));
INV_X1 slo__c380 (.ZN (slo__n361), .A (slo__n360));
NAND2_X4 i_0_1_218 (.ZN (n_0_316), .A1 (clk), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_217 (.ZN (n_0_315), .A1 (B[31]), .A2 (n_0_1_89));
AND2_X1 i_0_1_216 (.ZN (n_0_314), .A1 (B[30]), .A2 (n_0_1_89));
AND2_X1 i_0_1_215 (.ZN (n_0_313), .A1 (B[29]), .A2 (n_0_1_89));
AND2_X1 i_0_1_214 (.ZN (n_0_312), .A1 (B[28]), .A2 (n_0_1_89));
AND2_X1 i_0_1_213 (.ZN (n_0_311), .A1 (B[27]), .A2 (n_0_1_89));
AND2_X1 i_0_1_212 (.ZN (n_0_310), .A1 (B[26]), .A2 (n_0_1_89));
AND2_X1 i_0_1_211 (.ZN (n_0_309), .A1 (B[25]), .A2 (n_0_1_89));
AND2_X1 i_0_1_210 (.ZN (n_0_308), .A1 (B[24]), .A2 (n_0_1_89));
AND2_X1 i_0_1_209 (.ZN (n_0_307), .A1 (B[23]), .A2 (n_0_1_89));
AND2_X2 i_0_1_208 (.ZN (n_0_306), .A1 (B[22]), .A2 (n_0_1_89));
AND2_X1 i_0_1_207 (.ZN (n_0_305), .A1 (B[21]), .A2 (n_0_1_89));
AND2_X1 i_0_1_206 (.ZN (n_0_304), .A1 (B[20]), .A2 (n_0_1_89));
AND2_X1 i_0_1_205 (.ZN (n_0_303), .A1 (B[19]), .A2 (n_0_1_89));
AND2_X1 i_0_1_204 (.ZN (n_0_302), .A1 (B[18]), .A2 (n_0_1_89));
AND2_X1 i_0_1_203 (.ZN (n_0_301), .A1 (B[17]), .A2 (n_0_1_89));
AND2_X1 i_0_1_202 (.ZN (n_0_300), .A1 (B[16]), .A2 (n_0_1_89));
AND2_X1 i_0_1_201 (.ZN (n_0_299), .A1 (B[15]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_200 (.ZN (n_0_298), .A1 (B[14]), .A2 (n_0_1_89));
AND2_X1 i_0_1_199 (.ZN (n_0_297), .A1 (B[13]), .A2 (n_0_1_89));
AND2_X1 i_0_1_198 (.ZN (n_0_296), .A1 (B[12]), .A2 (n_0_1_89));
AND2_X1 i_0_1_197 (.ZN (n_0_295), .A1 (B[11]), .A2 (n_0_1_89));
AND2_X1 i_0_1_196 (.ZN (n_0_294), .A1 (B[10]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_195 (.ZN (n_0_293), .A1 (B[9]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_194 (.ZN (n_0_292), .A1 (B[8]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_193 (.ZN (n_0_291), .A1 (B[7]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_192 (.ZN (n_0_290), .A1 (B[6]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_191 (.ZN (n_0_289), .A1 (B[5]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_190 (.ZN (n_0_287), .A1 (B[4]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_189 (.ZN (n_0_286), .A1 (B[3]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_188 (.ZN (n_0_285), .A1 (B[2]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_187 (.ZN (n_0_284), .A1 (B[1]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_186 (.ZN (n_0_283), .A1 (B[0]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_185 (.ZN (n_0_281), .A1 (A[31]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_182 (.ZN (n_0_280), .A1 (A[30]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_181 (.ZN (n_0_279), .A1 (A[29]), .A2 (n_0_1_89));
AND2_X1 i_0_1_180 (.ZN (n_0_278), .A1 (A[28]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_179 (.ZN (n_0_277), .A1 (A[27]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_178 (.ZN (n_0_276), .A1 (A[26]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_177 (.ZN (n_0_275), .A1 (A[25]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_176 (.ZN (n_0_274), .A1 (A[24]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_175 (.ZN (n_0_273), .A1 (A[23]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_174 (.ZN (n_0_272), .A1 (A[22]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_173 (.ZN (n_0_271), .A1 (A[21]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_172 (.ZN (n_0_270), .A1 (A[20]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_171 (.ZN (n_0_269), .A1 (A[19]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_170 (.ZN (n_0_268), .A1 (A[18]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_169 (.ZN (n_0_267), .A1 (A[17]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_168 (.ZN (n_0_266), .A1 (A[16]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_167 (.ZN (n_0_265), .A1 (A[15]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_166 (.ZN (n_0_264), .A1 (A[14]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_165 (.ZN (n_0_263), .A1 (A[13]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_164 (.ZN (n_0_262), .A1 (A[12]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_163 (.ZN (n_0_261), .A1 (A[11]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_162 (.ZN (n_0_260), .A1 (A[10]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_161 (.ZN (n_0_259), .A1 (A[9]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_160 (.ZN (n_0_258), .A1 (A[8]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_159 (.ZN (n_0_257), .A1 (A[7]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_158 (.ZN (n_0_256), .A1 (A[6]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_157 (.ZN (n_0_255), .A1 (A[5]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_156 (.ZN (n_0_254), .A1 (A[4]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_155 (.ZN (n_0_253), .A1 (A[3]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_154 (.ZN (n_0_252), .A1 (A[2]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_153 (.ZN (n_0_251), .A1 (A[1]), .A2 (hfn_ipo_n125));
AND2_X1 i_0_1_152 (.ZN (n_0_250), .A1 (A[0]), .A2 (hfn_ipo_n125));
INV_X1 i_0_1_151 (.ZN (n_0_1_89), .A (reset));
AND2_X4 i_0_1_280 (.ZN (\B_imm[31] ), .A1 (drc_ipo_n167), .A2 (n_0_31));
MUX2_X1 i_0_1_279 (.Z (\B_imm[30] ), .A (n_0_126), .B (n_0_30), .S (drc_ipo_n167));
MUX2_X2 i_0_1_278 (.Z (\B_imm[29] ), .A (n_0_127), .B (n_0_29), .S (drc_ipo_n167));
MUX2_X1 i_0_1_277 (.Z (slo__n360), .A (n_0_128), .B (n_0_28), .S (drc_ipo_n167));
MUX2_X2 i_0_1_276 (.Z (\B_imm[27] ), .A (n_0_129), .B (n_0_27), .S (drc_ipo_n167));
MUX2_X1 i_0_1_275 (.Z (sgo__n273), .A (n_0_130), .B (n_0_26), .S (drc_ipo_n167));
MUX2_X1 i_0_1_274 (.Z (slo__n383), .A (n_0_131), .B (n_0_25), .S (drc_ipo_n167));
MUX2_X2 i_0_1_273 (.Z (\B_imm[24] ), .A (n_0_132), .B (n_0_24), .S (drc_ipo_n167));
MUX2_X1 i_0_1_272 (.Z (\B_imm[23] ), .A (n_0_133), .B (n_0_23), .S (drc_ipo_n167));
MUX2_X1 i_0_1_271 (.Z (\B_imm[22] ), .A (n_0_134), .B (n_0_22), .S (drc_ipo_n167));
MUX2_X1 i_0_1_270 (.Z (\B_imm[21] ), .A (n_0_135), .B (n_0_21), .S (drc_ipo_n167));
MUX2_X1 i_0_1_269 (.Z (\B_imm[20] ), .A (n_0_136), .B (n_0_20), .S (drc_ipo_n167));
MUX2_X1 i_0_1_268 (.Z (\B_imm[19] ), .A (n_0_137), .B (n_0_19), .S (drc_ipo_n167));
MUX2_X1 i_0_1_267 (.Z (\B_imm[18] ), .A (n_0_138), .B (n_0_18), .S (drc_ipo_n167));
MUX2_X1 i_0_1_266 (.Z (sgo__n219), .A (n_0_139), .B (n_0_17), .S (drc_ipo_n167));
MUX2_X1 i_0_1_265 (.Z (\B_imm[16] ), .A (n_0_140), .B (n_0_16), .S (drc_ipo_n167));
MUX2_X1 i_0_1_264 (.Z (\B_imm[15] ), .A (n_0_141), .B (n_0_15), .S (drc_ipo_n167));
MUX2_X1 i_0_1_263 (.Z (\B_imm[14] ), .A (n_0_142), .B (n_0_14), .S (drc_ipo_n167));
MUX2_X1 i_0_1_262 (.Z (\B_imm[13] ), .A (n_0_143), .B (n_0_13), .S (drc_ipo_n167));
MUX2_X1 i_0_1_261 (.Z (\B_imm[12] ), .A (n_0_144), .B (n_0_12), .S (drc_ipo_n167));
MUX2_X1 i_0_1_260 (.Z (\B_imm[11] ), .A (n_0_145), .B (n_0_11), .S (drc_ipo_n167));
MUX2_X2 i_0_1_259 (.Z (\B_imm[10] ), .A (n_0_146), .B (n_0_10), .S (drc_ipo_n167));
MUX2_X1 i_0_1_258 (.Z (\B_imm[9] ), .A (n_0_147), .B (n_0_9), .S (drc_ipo_n167));
MUX2_X1 i_0_1_257 (.Z (\B_imm[8] ), .A (n_0_148), .B (n_0_8), .S (drc_ipo_n167));
MUX2_X1 i_0_1_256 (.Z (\B_imm[7] ), .A (n_0_149), .B (n_0_7), .S (drc_ipo_n167));
MUX2_X1 i_0_1_255 (.Z (\B_imm[6] ), .A (n_0_150), .B (n_0_6), .S (drc_ipo_n167));
MUX2_X1 i_0_1_254 (.Z (sgo__n307), .A (n_0_151), .B (n_0_5), .S (drc_ipo_n167));
MUX2_X1 i_0_1_253 (.Z (\B_imm[4] ), .A (CLOCK_opt_ipo_n663), .B (n_0_4), .S (drc_ipo_n167));
MUX2_X1 i_0_1_252 (.Z (sgo__n237), .A (n_0_153), .B (n_0_3), .S (drc_ipo_n167));
MUX2_X2 i_0_1_251 (.Z (\B_imm[2] ), .A (n_0_154), .B (n_0_2), .S (drc_ipo_n167));
MUX2_X2 i_0_1_250 (.Z (\B_imm[1] ), .A (n_0_155), .B (n_0_1), .S (drc_ipo_n167));
AND2_X4 i_0_1_249 (.ZN (\A_imm[31] ), .A1 (drc_ipo_n165), .A2 (n_0_62));
MUX2_X1 i_0_1_248 (.Z (\A_imm[30] ), .A (n_0_156), .B (n_0_61), .S (drc_ipo_n165));
MUX2_X2 i_0_1_247 (.Z (\A_imm[29] ), .A (n_0_157), .B (n_0_60), .S (drc_ipo_n165));
MUX2_X1 i_0_1_246 (.Z (slo__n366), .A (n_0_158), .B (n_0_59), .S (drc_ipo_n165));
MUX2_X1 i_0_1_245 (.Z (\A_imm[27] ), .A (n_0_159), .B (n_0_58), .S (drc_ipo_n165));
MUX2_X1 i_0_1_244 (.Z (\A_imm[26] ), .A (n_0_160), .B (n_0_57), .S (drc_ipo_n165));
MUX2_X1 i_0_1_243 (.Z (sgo__n269), .A (n_0_161), .B (n_0_56), .S (drc_ipo_n165));
MUX2_X1 i_0_1_242 (.Z (sgo__n291), .A (n_0_162), .B (n_0_55), .S (drc_ipo_n165));
MUX2_X1 i_0_1_241 (.Z (\A_imm[23] ), .A (n_0_163), .B (n_0_54), .S (drc_ipo_n165));
MUX2_X1 i_0_1_240 (.Z (\A_imm[22] ), .A (n_0_164), .B (n_0_53), .S (drc_ipo_n165));
MUX2_X2 i_0_1_239 (.Z (\A_imm[21] ), .A (n_0_165), .B (n_0_52), .S (drc_ipo_n165));
MUX2_X1 i_0_1_238 (.Z (\A_imm[20] ), .A (n_0_166), .B (n_0_51), .S (drc_ipo_n165));
MUX2_X1 i_0_1_237 (.Z (\A_imm[19] ), .A (n_0_167), .B (n_0_50), .S (drc_ipo_n165));
MUX2_X1 i_0_1_236 (.Z (\A_imm[18] ), .A (n_0_168), .B (n_0_49), .S (drc_ipo_n165));
MUX2_X2 i_0_1_235 (.Z (sgo__n175), .A (n_0_169), .B (n_0_48), .S (drc_ipo_n165));
MUX2_X2 i_0_1_234 (.Z (\A_imm[16] ), .A (n_0_170), .B (n_0_47), .S (drc_ipo_n165));
MUX2_X2 i_0_1_233 (.Z (\A_imm[15] ), .A (n_0_171), .B (n_0_46), .S (drc_ipo_n165));
MUX2_X2 i_0_1_232 (.Z (\A_imm[14] ), .A (n_0_172), .B (n_0_45), .S (drc_ipo_n165));
MUX2_X1 i_0_1_231 (.Z (\A_imm[13] ), .A (n_0_173), .B (n_0_44), .S (drc_ipo_n165));
MUX2_X1 i_0_1_230 (.Z (\A_imm[12] ), .A (n_0_174), .B (n_0_43), .S (drc_ipo_n165));
MUX2_X1 i_0_1_229 (.Z (\A_imm[11] ), .A (n_0_175), .B (n_0_42), .S (drc_ipo_n165));
MUX2_X1 i_0_1_228 (.Z (\A_imm[10] ), .A (n_0_176), .B (n_0_41), .S (drc_ipo_n165));
MUX2_X1 i_0_1_227 (.Z (\A_imm[9] ), .A (n_0_177), .B (n_0_40), .S (drc_ipo_n165));
MUX2_X1 i_0_1_226 (.Z (\A_imm[8] ), .A (CLOCK_opt_ipo_n660), .B (n_0_39), .S (drc_ipo_n165));
MUX2_X1 i_0_1_225 (.Z (\A_imm[7] ), .A (n_0_179), .B (n_0_38), .S (drc_ipo_n165));
MUX2_X1 i_0_1_224 (.Z (\A_imm[6] ), .A (n_0_180), .B (n_0_37), .S (drc_ipo_n165));
MUX2_X1 i_0_1_223 (.Z (\A_imm[5] ), .A (n_0_181), .B (n_0_36), .S (drc_ipo_n165));
MUX2_X2 i_0_1_222 (.Z (\A_imm[4] ), .A (n_0_182), .B (n_0_35), .S (drc_ipo_n165));
MUX2_X1 i_0_1_221 (.Z (\A_imm[3] ), .A (n_0_183), .B (n_0_34), .S (drc_ipo_n165));
MUX2_X1 i_0_1_220 (.Z (\A_imm[2] ), .A (n_0_184), .B (n_0_33), .S (drc_ipo_n165));
MUX2_X2 i_0_1_219 (.Z (\A_imm[1] ), .A (n_0_185), .B (n_0_32), .S (drc_ipo_n165));
AOI21_X1 i_0_1_184 (.ZN (CTS_n770), .A (reset), .B1 (clk), .B2 (CLOCK_slh_n1056));
INV_X4 CTS_L2_remove_c626 (.ZN (CTS_n769), .A (CTS_n770));
INV_X4 sgo__c332 (.ZN (\A_imm[24] ), .A (sgo__n292));
NOR4_X2 i_0_1_149 (.ZN (n_0_1_85), .A1 (\Res_imm[52] ), .A2 (\Res_imm[53] ), .A3 (CLOCK_opt_ipo_n666), .A4 (\Res_imm[50] ));
NOR4_X2 i_0_1_148 (.ZN (n_0_1_84), .A1 (\Res_imm[63] ), .A2 (\Res_imm[62] ), .A3 (\Res_imm[57] ), .A4 (\Res_imm[32] ));
INV_X1 sgo__c303 (.ZN (sgo__n274), .A (sgo__n273));
INV_X1 sgo__c351 (.ZN (sgo__n308), .A (sgo__n307));
NOR4_X2 i_0_1_145 (.ZN (n_0_1_81), .A1 (\Res_imm[48] ), .A2 (\Res_imm[39] ), .A3 (\Res_imm[38] ), .A4 (\Res_imm[37] ));
NOR4_X2 i_0_1_144 (.ZN (n_0_1_80), .A1 (\Res_imm[36] ), .A2 (\Res_imm[35] ), .A3 (\Res_imm[34] ), .A4 (\Res_imm[33] ));
INV_X1 sgo__c299 (.ZN (sgo__n270), .A (sgo__n269));
NOR4_X4 i_0_1_142 (.ZN (n_0_1_78), .A1 (\Res_imm[44] ), .A2 (\Res_imm[43] ), .A3 (\Res_imm[42] ), .A4 (\Res_imm[41] ));
NAND4_X2 i_0_1_141 (.ZN (n_0_1_77), .A1 (n_0_1_81), .A2 (n_0_1_80), .A3 (sgo__sro_n179), .A4 (n_0_1_78));
NOR4_X2 i_0_1_140 (.ZN (n_0_1_76), .A1 (\Res_imm[23] ), .A2 (\Res_imm[22] ), .A3 (\Res_imm[21] ), .A4 (\Res_imm[16] ));
NOR4_X1 i_0_1_139 (.ZN (n_0_1_75), .A1 (\Res_imm[20] ), .A2 (\Res_imm[19] ), .A3 (\Res_imm[18] ), .A4 (\Res_imm[17] ));
NOR4_X1 i_0_1_138 (.ZN (n_0_1_74), .A1 (\Res_imm[31] ), .A2 (\Res_imm[30] ), .A3 (\Res_imm[29] ), .A4 (\Res_imm[24] ));
NOR4_X2 i_0_1_137 (.ZN (n_0_1_73), .A1 (\Res_imm[28] ), .A2 (\Res_imm[27] ), .A3 (\Res_imm[26] ), .A4 (\Res_imm[25] ));
NAND4_X1 i_0_1_136 (.ZN (n_0_1_72), .A1 (n_0_1_76), .A2 (n_0_1_75), .A3 (n_0_1_74), .A4 (n_0_1_73));
NOR4_X1 i_0_1_135 (.ZN (n_0_1_71), .A1 (\Res_imm[15] ), .A2 (\Res_imm[7] ), .A3 (\Res_imm[6] ), .A4 (\Res_imm[5] ));
NOR4_X1 i_0_1_134 (.ZN (n_0_1_70), .A1 (\Res_imm[4] ), .A2 (\Res_imm[3] ), .A3 (\Res_imm[2] ), .A4 (\Res_imm[1] ));
NOR4_X1 i_0_1_133 (.ZN (n_0_1_69), .A1 (\Res_imm[14] ), .A2 (\Res_imm[13] ), .A3 (\Res_imm[8] ), .A4 (\Res_imm[0] ));
NOR4_X1 i_0_1_132 (.ZN (n_0_1_68), .A1 (\Res_imm[12] ), .A2 (\Res_imm[11] ), .A3 (\Res_imm[10] ), .A4 (\Res_imm[9] ));
NAND4_X1 i_0_1_131 (.ZN (n_0_1_67), .A1 (n_0_1_71), .A2 (n_0_1_70), .A3 (n_0_1_69), .A4 (n_0_1_68));
NOR2_X1 sgo__sro_c283 (.ZN (sgo__sro_n257), .A1 (\Res_imm[55] ), .A2 (\Res_imm[56] ));
XOR2_X1 i_0_1_129 (.Z (n_0_1_65), .A (drc_ipo_n167), .B (drc_ipo_n165));
AND3_X4 i_0_1_128 (.ZN (n_0_1_64), .A1 (n_0_1_89), .A2 (n_0_1_66), .A3 (n_0_1_65));
AOI21_X2 i_0_1_127 (.ZN (n_0_1_63), .A (reset), .B1 (n_0_1_66), .B2 (n_0_1_65));
AOI22_X1 i_0_1_126 (.ZN (n_0_1_62), .A1 (n_0_125), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[63] ));
INV_X1 i_0_1_125 (.ZN (n_0_249), .A (n_0_1_62));
AOI22_X1 i_0_1_124 (.ZN (n_0_1_61), .A1 (n_0_124), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[62] ));
INV_X1 i_0_1_123 (.ZN (n_0_248), .A (n_0_1_61));
AOI22_X1 i_0_1_122 (.ZN (n_0_1_60), .A1 (n_0_123), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[61] ));
INV_X1 i_0_1_121 (.ZN (n_0_247), .A (n_0_1_60));
AOI22_X1 i_0_1_120 (.ZN (n_0_1_59), .A1 (n_0_122), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[60] ));
INV_X1 i_0_1_119 (.ZN (n_0_246), .A (n_0_1_59));
AOI22_X1 i_0_1_118 (.ZN (n_0_1_58), .A1 (n_0_121), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[59] ));
INV_X1 i_0_1_117 (.ZN (n_0_245), .A (n_0_1_58));
AOI22_X1 i_0_1_116 (.ZN (n_0_1_57), .A1 (n_0_120), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[58] ));
INV_X1 i_0_1_115 (.ZN (n_0_244), .A (n_0_1_57));
AOI22_X1 i_0_1_114 (.ZN (n_0_1_56), .A1 (n_0_119), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[57] ));
INV_X1 i_0_1_113 (.ZN (n_0_243), .A (n_0_1_56));
AOI22_X1 i_0_1_112 (.ZN (n_0_1_55), .A1 (n_0_118), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[56] ));
INV_X1 i_0_1_111 (.ZN (n_0_242), .A (n_0_1_55));
AOI22_X1 i_0_1_110 (.ZN (n_0_1_54), .A1 (n_0_117), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[55] ));
INV_X1 i_0_1_109 (.ZN (n_0_241), .A (n_0_1_54));
AOI22_X1 i_0_1_108 (.ZN (n_0_1_53), .A1 (n_0_116), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[54] ));
INV_X1 i_0_1_107 (.ZN (n_0_240), .A (n_0_1_53));
AOI22_X1 i_0_1_106 (.ZN (n_0_1_52), .A1 (n_0_115), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[53] ));
INV_X1 i_0_1_105 (.ZN (n_0_239), .A (n_0_1_52));
AOI22_X1 i_0_1_104 (.ZN (n_0_1_51), .A1 (n_0_114), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[52] ));
INV_X1 i_0_1_103 (.ZN (n_0_238), .A (n_0_1_51));
AOI22_X1 i_0_1_102 (.ZN (n_0_1_50), .A1 (n_0_113), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (CLOCK_opt_ipo_n666));
INV_X1 i_0_1_101 (.ZN (n_0_237), .A (n_0_1_50));
AOI22_X2 i_0_1_100 (.ZN (n_0_1_49), .A1 (n_0_112), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[50] ));
INV_X1 i_0_1_99 (.ZN (n_0_236), .A (n_0_1_49));
AOI22_X1 i_0_1_98 (.ZN (n_0_1_48), .A1 (n_0_111), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[49] ));
INV_X1 i_0_1_97 (.ZN (n_0_235), .A (n_0_1_48));
AOI22_X1 i_0_1_96 (.ZN (n_0_1_47), .A1 (n_0_110), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[48] ));
INV_X1 i_0_1_95 (.ZN (n_0_234), .A (n_0_1_47));
AOI22_X1 i_0_1_94 (.ZN (n_0_1_46), .A1 (n_0_109), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[47] ));
INV_X1 i_0_1_93 (.ZN (n_0_233), .A (n_0_1_46));
AOI22_X1 i_0_1_92 (.ZN (n_0_1_45), .A1 (n_0_108), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[46] ));
INV_X1 i_0_1_91 (.ZN (n_0_232), .A (n_0_1_45));
AOI22_X1 i_0_1_90 (.ZN (n_0_1_44), .A1 (n_0_107), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[45] ));
INV_X1 i_0_1_89 (.ZN (n_0_231), .A (n_0_1_44));
AOI22_X1 i_0_1_88 (.ZN (n_0_1_43), .A1 (n_0_106), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[44] ));
INV_X1 i_0_1_87 (.ZN (n_0_230), .A (n_0_1_43));
AOI22_X1 i_0_1_86 (.ZN (n_0_1_42), .A1 (n_0_105), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[43] ));
INV_X1 i_0_1_85 (.ZN (n_0_229), .A (n_0_1_42));
AOI22_X1 i_0_1_84 (.ZN (n_0_1_41), .A1 (n_0_104), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[42] ));
INV_X1 i_0_1_83 (.ZN (n_0_228), .A (n_0_1_41));
AOI22_X1 i_0_1_82 (.ZN (n_0_1_40), .A1 (n_0_103), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[41] ));
INV_X1 i_0_1_81 (.ZN (n_0_227), .A (n_0_1_40));
AOI22_X1 i_0_1_80 (.ZN (n_0_1_39), .A1 (n_0_102), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[40] ));
INV_X1 i_0_1_79 (.ZN (n_0_226), .A (n_0_1_39));
AOI22_X1 i_0_1_78 (.ZN (n_0_1_38), .A1 (n_0_101), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[39] ));
INV_X1 i_0_1_77 (.ZN (n_0_225), .A (n_0_1_38));
AOI22_X1 i_0_1_76 (.ZN (n_0_1_37), .A1 (n_0_100), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[38] ));
INV_X1 i_0_1_75 (.ZN (n_0_224), .A (n_0_1_37));
AOI22_X1 i_0_1_74 (.ZN (n_0_1_36), .A1 (n_0_99), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[37] ));
INV_X1 i_0_1_73 (.ZN (n_0_223), .A (n_0_1_36));
AOI22_X1 i_0_1_72 (.ZN (n_0_1_35), .A1 (n_0_98), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[36] ));
INV_X1 i_0_1_71 (.ZN (n_0_222), .A (n_0_1_35));
AOI22_X1 i_0_1_70 (.ZN (n_0_1_34), .A1 (n_0_97), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[35] ));
INV_X1 i_0_1_69 (.ZN (n_0_221), .A (n_0_1_34));
AOI22_X2 i_0_1_68 (.ZN (n_0_1_33), .A1 (n_0_96), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[34] ));
INV_X1 i_0_1_67 (.ZN (n_0_220), .A (n_0_1_33));
AOI22_X1 i_0_1_66 (.ZN (n_0_1_32), .A1 (n_0_95), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[33] ));
INV_X1 i_0_1_65 (.ZN (n_0_219), .A (n_0_1_32));
AOI22_X1 i_0_1_64 (.ZN (n_0_1_31), .A1 (n_0_94), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[32] ));
INV_X1 i_0_1_63 (.ZN (n_0_218), .A (n_0_1_31));
AOI22_X1 i_0_1_62 (.ZN (n_0_1_30), .A1 (n_0_93), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[31] ));
INV_X1 i_0_1_61 (.ZN (n_0_217), .A (n_0_1_30));
AOI22_X1 i_0_1_60 (.ZN (n_0_1_29), .A1 (n_0_92), .A2 (hfn_ipo_n123), .B1 (hfn_ipo_n121), .B2 (\Res_imm[30] ));
INV_X1 i_0_1_59 (.ZN (n_0_216), .A (n_0_1_29));
AOI22_X1 i_0_1_58 (.ZN (n_0_1_28), .A1 (n_0_91), .A2 (n_0_1_64), .B1 (hfn_ipo_n120), .B2 (\Res_imm[29] ));
INV_X1 i_0_1_57 (.ZN (n_0_215), .A (n_0_1_28));
AOI22_X1 i_0_1_56 (.ZN (n_0_1_27), .A1 (n_0_90), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[28] ));
INV_X1 i_0_1_55 (.ZN (n_0_214), .A (n_0_1_27));
AOI22_X1 i_0_1_54 (.ZN (n_0_1_26), .A1 (n_0_89), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[27] ));
INV_X1 i_0_1_53 (.ZN (n_0_213), .A (n_0_1_26));
AOI22_X1 i_0_1_52 (.ZN (n_0_1_25), .A1 (n_0_88), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[26] ));
INV_X1 i_0_1_51 (.ZN (n_0_212), .A (n_0_1_25));
AOI22_X1 i_0_1_50 (.ZN (n_0_1_24), .A1 (n_0_87), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[25] ));
INV_X1 i_0_1_49 (.ZN (n_0_211), .A (n_0_1_24));
AOI22_X1 i_0_1_48 (.ZN (n_0_1_23), .A1 (n_0_86), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[24] ));
INV_X1 i_0_1_47 (.ZN (n_0_210), .A (n_0_1_23));
AOI22_X1 i_0_1_46 (.ZN (n_0_1_22), .A1 (n_0_85), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[23] ));
INV_X1 i_0_1_45 (.ZN (n_0_209), .A (n_0_1_22));
AOI22_X1 i_0_1_44 (.ZN (n_0_1_21), .A1 (n_0_84), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[22] ));
INV_X1 i_0_1_43 (.ZN (n_0_208), .A (n_0_1_21));
AOI22_X1 i_0_1_42 (.ZN (n_0_1_20), .A1 (n_0_83), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[21] ));
INV_X1 i_0_1_41 (.ZN (n_0_207), .A (n_0_1_20));
AOI22_X1 i_0_1_40 (.ZN (n_0_1_19), .A1 (n_0_82), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[20] ));
INV_X1 i_0_1_39 (.ZN (n_0_206), .A (n_0_1_19));
AOI22_X1 i_0_1_38 (.ZN (n_0_1_18), .A1 (n_0_81), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[19] ));
INV_X1 i_0_1_37 (.ZN (n_0_205), .A (n_0_1_18));
AOI22_X1 i_0_1_36 (.ZN (n_0_1_17), .A1 (n_0_80), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[18] ));
INV_X1 i_0_1_35 (.ZN (n_0_204), .A (n_0_1_17));
AOI22_X1 i_0_1_34 (.ZN (n_0_1_16), .A1 (n_0_79), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[17] ));
INV_X1 i_0_1_33 (.ZN (n_0_203), .A (n_0_1_16));
AOI22_X1 i_0_1_32 (.ZN (n_0_1_15), .A1 (n_0_78), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[16] ));
INV_X1 i_0_1_31 (.ZN (n_0_202), .A (n_0_1_15));
AOI22_X1 i_0_1_30 (.ZN (n_0_1_14), .A1 (n_0_77), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[15] ));
INV_X1 i_0_1_29 (.ZN (n_0_201), .A (n_0_1_14));
AOI22_X4 i_0_1_28 (.ZN (n_0_1_13), .A1 (n_0_76), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[14] ));
CLKBUF_X1 CLOCK_slh__c813 (.Z (sph__n1165), .A (CLOCK_slh__n1107));
AOI22_X4 i_0_1_26 (.ZN (n_0_1_12), .A1 (n_0_75), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[13] ));
CLKBUF_X1 CLOCK_slh__c811 (.Z (CLOCK_slh__n1106), .A (CLOCK_slh__n1105));
AOI22_X1 i_0_1_24 (.ZN (n_0_1_11), .A1 (CLOCK_opt_ipo_n697), .A2 (n_0_74), .B1 (hfn_ipo_n120), .B2 (\Res_imm[12] ));
INV_X1 i_0_1_23 (.ZN (n_0_198), .A (n_0_1_11));
AOI22_X2 i_0_1_22 (.ZN (n_0_1_10), .A1 (n_0_73), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[11] ));
INV_X1 i_0_1_21 (.ZN (n_0_197), .A (n_0_1_10));
AOI22_X2 i_0_1_20 (.ZN (n_0_1_9), .A1 (n_0_72), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[10] ));
INV_X1 i_0_1_19 (.ZN (n_0_196), .A (n_0_1_9));
AOI22_X4 i_0_1_18 (.ZN (n_0_1_8), .A1 (n_0_71), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[9] ));
CLKBUF_X1 CLOCK_slh__c784 (.Z (CLOCK_slh__n1079), .A (CLOCK_slh__n1078));
AOI22_X2 i_0_1_16 (.ZN (n_0_1_7), .A1 (n_0_70), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[8] ));
INV_X1 i_0_1_15 (.ZN (n_0_194), .A (n_0_1_7));
AOI22_X4 i_0_1_14 (.ZN (n_0_1_6), .A1 (n_0_69), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[7] ));
CLKBUF_X1 CLOCK_slh__c785 (.Z (CLOCK_slh__n1087), .A (CLOCK_slh__n1079));
AOI22_X2 i_0_1_12 (.ZN (n_0_1_5), .A1 (n_0_68), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[6] ));
INV_X1 i_0_1_11 (.ZN (n_0_192), .A (n_0_1_5));
AOI22_X2 i_0_1_10 (.ZN (n_0_1_4), .A1 (n_0_67), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[5] ));
INV_X1 i_0_1_9 (.ZN (n_0_191), .A (n_0_1_4));
AOI22_X2 i_0_1_8 (.ZN (n_0_1_3), .A1 (n_0_66), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[4] ));
INV_X1 i_0_1_7 (.ZN (n_0_190), .A (n_0_1_3));
AOI22_X4 i_0_1_6 (.ZN (n_0_1_2), .A1 (n_0_65), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[3] ));
AOI22_X4 i_0_1_4 (.ZN (n_0_1_1), .A1 (n_0_64), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[2] ));
CLKBUF_X1 sph__c872 (.Z (CLOCK_slh_n1056), .A (sph__n1166));
AOI22_X4 i_0_1_2 (.ZN (n_0_1_0), .A1 (n_0_63), .A2 (CLOCK_opt_ipo_n697), .B1 (hfn_ipo_n120), .B2 (\Res_imm[1] ));
CLKBUF_X1 sph__c871 (.Z (sph__n1166), .A (sph__n1165));
AND2_X1 i_0_1_0 (.ZN (n_0_186), .A1 (hfn_ipo_n125), .A2 (\Res_imm[0] ));
DLH_X2 \A_in_reg[0]  (.Q (n_0_0), .D (n_0_250), .G (CTS_n769));
DLH_X2 \A_in_reg[1]  (.Q (n_0_185), .D (n_0_251), .G (CTS_n769));
DLH_X1 \A_in_reg[2]  (.Q (n_0_184), .D (n_0_252), .G (CTS_n769));
DLH_X1 \A_in_reg[3]  (.Q (n_0_183), .D (n_0_253), .G (CTS_n769));
DLH_X2 \A_in_reg[4]  (.Q (n_0_182), .D (n_0_254), .G (CTS_n769));
DLH_X1 \A_in_reg[5]  (.Q (n_0_181), .D (n_0_255), .G (CTS_n769));
DLH_X1 \A_in_reg[6]  (.Q (n_0_180), .D (n_0_256), .G (CTS_n769));
DLH_X1 \A_in_reg[7]  (.Q (n_0_179), .D (n_0_257), .G (CTS_n769));
DLH_X1 \A_in_reg[8]  (.Q (n_0_178), .D (n_0_258), .G (CTS_n769));
DLH_X1 \A_in_reg[9]  (.Q (n_0_177), .D (n_0_259), .G (CTS_n769));
DLH_X1 \A_in_reg[10]  (.Q (n_0_176), .D (n_0_260), .G (CTS_n769));
DLH_X1 \A_in_reg[11]  (.Q (n_0_175), .D (n_0_261), .G (CTS_n769));
DLH_X1 \A_in_reg[12]  (.Q (n_0_174), .D (n_0_262), .G (CTS_n769));
DLH_X1 \A_in_reg[13]  (.Q (n_0_173), .D (n_0_263), .G (CTS_n769));
DLH_X1 \A_in_reg[14]  (.Q (n_0_172), .D (n_0_264), .G (CTS_n769));
DLH_X1 \A_in_reg[15]  (.Q (n_0_171), .D (n_0_265), .G (CTS_n769));
DLH_X1 \A_in_reg[16]  (.Q (n_0_170), .D (n_0_266), .G (CTS_n769));
DLH_X1 \A_in_reg[17]  (.Q (n_0_169), .D (n_0_267), .G (CTS_n769));
DLH_X1 \A_in_reg[18]  (.Q (n_0_168), .D (n_0_268), .G (CTS_n769));
DLH_X1 \A_in_reg[19]  (.Q (n_0_167), .D (n_0_269), .G (CTS_n769));
DLH_X1 \A_in_reg[20]  (.Q (n_0_166), .D (n_0_270), .G (CTS_n769));
DLH_X1 \A_in_reg[21]  (.Q (n_0_165), .D (n_0_271), .G (CTS_n769));
DLH_X1 \A_in_reg[22]  (.Q (n_0_164), .D (n_0_272), .G (CTS_n769));
DLH_X1 \A_in_reg[23]  (.Q (n_0_163), .D (n_0_273), .G (CTS_n769));
DLH_X1 \A_in_reg[24]  (.Q (n_0_162), .D (n_0_274), .G (CTS_n769));
DLH_X1 \A_in_reg[25]  (.Q (n_0_161), .D (n_0_275), .G (CTS_n769));
DLH_X1 \A_in_reg[26]  (.Q (n_0_160), .D (n_0_276), .G (CTS_n769));
DLH_X1 \A_in_reg[27]  (.Q (n_0_159), .D (n_0_277), .G (CTS_n769));
DLH_X1 \A_in_reg[28]  (.Q (n_0_158), .D (n_0_278), .G (CTS_n769));
DLH_X1 \A_in_reg[29]  (.Q (n_0_157), .D (n_0_279), .G (CTS_n769));
DLH_X1 \A_in_reg[30]  (.Q (n_0_156), .D (n_0_280), .G (CTS_n769));
DLH_X1 \A_in_reg[31]  (.Q (A_in), .D (n_0_281), .G (CTS_n769));
DLH_X2 \B_in_reg[0]  (.Q (n_0_288), .D (n_0_283), .G (CTS_n769));
DLH_X1 \B_in_reg[1]  (.Q (n_0_155), .D (n_0_284), .G (CTS_n769));
DLH_X1 \B_in_reg[2]  (.Q (n_0_154), .D (n_0_285), .G (CTS_n769));
DLH_X1 \B_in_reg[3]  (.Q (n_0_153), .D (n_0_286), .G (CTS_n769));
DLH_X1 \B_in_reg[4]  (.Q (n_0_152), .D (n_0_287), .G (CTS_n769));
DLH_X2 \B_in_reg[5]  (.Q (n_0_151), .D (n_0_289), .G (CTS_n769));
DLH_X1 \B_in_reg[6]  (.Q (n_0_150), .D (n_0_290), .G (CTS_n769));
DLH_X1 \B_in_reg[7]  (.Q (n_0_149), .D (n_0_291), .G (CTS_n769));
DLH_X1 \B_in_reg[8]  (.Q (n_0_148), .D (n_0_292), .G (CTS_n769));
DLH_X1 \B_in_reg[9]  (.Q (n_0_147), .D (n_0_293), .G (CTS_n769));
DLH_X1 \B_in_reg[10]  (.Q (n_0_146), .D (n_0_294), .G (CTS_n769));
DLH_X1 \B_in_reg[11]  (.Q (n_0_145), .D (n_0_295), .G (CTS_n769));
DLH_X1 \B_in_reg[12]  (.Q (n_0_144), .D (n_0_296), .G (CTS_n769));
DLH_X1 \B_in_reg[13]  (.Q (n_0_143), .D (n_0_297), .G (CTS_n769));
DLH_X1 \B_in_reg[14]  (.Q (n_0_142), .D (n_0_298), .G (CTS_n769));
DLH_X1 \B_in_reg[15]  (.Q (n_0_141), .D (n_0_299), .G (CTS_n769));
DLH_X1 \B_in_reg[16]  (.Q (n_0_140), .D (n_0_300), .G (CTS_n769));
DLH_X1 \B_in_reg[17]  (.Q (n_0_139), .D (n_0_301), .G (CTS_n769));
DLH_X1 \B_in_reg[18]  (.Q (n_0_138), .D (n_0_302), .G (CTS_n769));
DLH_X1 \B_in_reg[19]  (.Q (n_0_137), .D (n_0_303), .G (CTS_n769));
DLH_X1 \B_in_reg[20]  (.Q (n_0_136), .D (n_0_304), .G (CTS_n769));
DLH_X1 \B_in_reg[21]  (.Q (n_0_135), .D (n_0_305), .G (CTS_n769));
DLH_X1 \B_in_reg[22]  (.Q (n_0_134), .D (n_0_306), .G (CTS_n769));
DLH_X1 \B_in_reg[23]  (.Q (n_0_133), .D (n_0_307), .G (CTS_n769));
DLH_X1 \B_in_reg[24]  (.Q (n_0_132), .D (n_0_308), .G (CTS_n769));
DLH_X1 \B_in_reg[25]  (.Q (n_0_131), .D (n_0_309), .G (CTS_n769));
DLH_X1 \B_in_reg[26]  (.Q (n_0_130), .D (n_0_310), .G (CTS_n769));
DLH_X1 \B_in_reg[27]  (.Q (n_0_129), .D (n_0_311), .G (CTS_n769));
DLH_X1 \B_in_reg[28]  (.Q (n_0_128), .D (n_0_312), .G (CTS_n769));
DLH_X1 \B_in_reg[29]  (.Q (n_0_127), .D (n_0_313), .G (CTS_n769));
DLH_X1 \B_in_reg[30]  (.Q (n_0_126), .D (n_0_314), .G (CTS_n769));
DLH_X1 \B_in_reg[31]  (.Q (B_in), .D (n_0_315), .G (CTS_n769));
DLH_X1 \Res_reg[0]  (.Q (Res[0]), .D (n_0_186), .G (n_0_316));
DLH_X1 \Res_reg[1]  (.Q (Res[1]), .D (CLOCK_opt_ipo_n701), .G (n_0_316));
DLH_X1 \Res_reg[2]  (.Q (Res[2]), .D (CLOCK_opt_ipo_n703), .G (n_0_316));
DLH_X1 \Res_reg[3]  (.Q (Res[3]), .D (CLOCK_opt_ipo_n705), .G (n_0_316));
DLH_X1 \Res_reg[4]  (.Q (Res[4]), .D (n_0_190), .G (n_0_316));
DLH_X1 \Res_reg[5]  (.Q (Res[5]), .D (n_0_191), .G (n_0_316));
DLH_X1 \Res_reg[6]  (.Q (Res[6]), .D (n_0_192), .G (n_0_316));
DLH_X1 \Res_reg[7]  (.Q (Res[7]), .D (CLOCK_opt_ipo_n651), .G (n_0_316));
DLH_X1 \Res_reg[8]  (.Q (Res[8]), .D (n_0_194), .G (n_0_316));
DLH_X1 \Res_reg[9]  (.Q (Res[9]), .D (CLOCK_opt_ipo_n649), .G (n_0_316));
DLH_X1 \Res_reg[10]  (.Q (Res[10]), .D (n_0_196), .G (n_0_316));
DLH_X1 \Res_reg[11]  (.Q (Res[11]), .D (n_0_197), .G (n_0_316));
DLH_X1 \Res_reg[12]  (.Q (Res[12]), .D (n_0_198), .G (n_0_316));
DLH_X1 \Res_reg[13]  (.Q (Res[13]), .D (CLOCK_opt_ipo_n695), .G (n_0_316));
DLH_X1 \Res_reg[14]  (.Q (Res[14]), .D (CLOCK_opt_ipo_n699), .G (n_0_316));
DLH_X1 \Res_reg[15]  (.Q (Res[15]), .D (n_0_201), .G (n_0_316));
DLH_X1 \Res_reg[16]  (.Q (Res[16]), .D (n_0_202), .G (n_0_316));
DLH_X1 \Res_reg[17]  (.Q (Res[17]), .D (n_0_203), .G (n_0_316));
DLH_X1 \Res_reg[18]  (.Q (Res[18]), .D (n_0_204), .G (n_0_316));
DLH_X1 \Res_reg[19]  (.Q (Res[19]), .D (n_0_205), .G (n_0_316));
DLH_X1 \Res_reg[20]  (.Q (Res[20]), .D (n_0_206), .G (n_0_316));
DLH_X1 \Res_reg[21]  (.Q (Res[21]), .D (n_0_207), .G (n_0_316));
DLH_X1 \Res_reg[22]  (.Q (Res[22]), .D (n_0_208), .G (n_0_316));
DLH_X1 \Res_reg[23]  (.Q (Res[23]), .D (n_0_209), .G (n_0_316));
DLH_X1 \Res_reg[24]  (.Q (Res[24]), .D (n_0_210), .G (n_0_316));
DLH_X1 \Res_reg[25]  (.Q (Res[25]), .D (n_0_211), .G (n_0_316));
DLH_X1 \Res_reg[26]  (.Q (Res[26]), .D (n_0_212), .G (n_0_316));
DLH_X1 \Res_reg[27]  (.Q (Res[27]), .D (n_0_213), .G (n_0_316));
DLH_X1 \Res_reg[28]  (.Q (Res[28]), .D (n_0_214), .G (n_0_316));
DLH_X1 \Res_reg[29]  (.Q (Res[29]), .D (n_0_215), .G (n_0_316));
DLH_X1 \Res_reg[30]  (.Q (Res[30]), .D (n_0_216), .G (n_0_316));
DLH_X1 \Res_reg[31]  (.Q (Res[31]), .D (n_0_217), .G (n_0_316));
DLH_X1 \Res_reg[32]  (.Q (Res[32]), .D (n_0_218), .G (n_0_316));
DLH_X1 \Res_reg[33]  (.Q (Res[33]), .D (n_0_219), .G (n_0_316));
DLH_X1 \Res_reg[34]  (.Q (Res[34]), .D (n_0_220), .G (n_0_316));
DLH_X1 \Res_reg[35]  (.Q (Res[35]), .D (n_0_221), .G (n_0_316));
DLH_X1 \Res_reg[36]  (.Q (Res[36]), .D (n_0_222), .G (n_0_316));
DLH_X1 \Res_reg[37]  (.Q (Res[37]), .D (n_0_223), .G (n_0_316));
DLH_X1 \Res_reg[38]  (.Q (Res[38]), .D (n_0_224), .G (n_0_316));
DLH_X1 \Res_reg[39]  (.Q (Res[39]), .D (n_0_225), .G (n_0_316));
DLH_X1 \Res_reg[40]  (.Q (Res[40]), .D (n_0_226), .G (n_0_316));
DLH_X1 \Res_reg[41]  (.Q (Res[41]), .D (n_0_227), .G (n_0_316));
DLH_X1 \Res_reg[42]  (.Q (Res[42]), .D (n_0_228), .G (n_0_316));
DLH_X1 \Res_reg[43]  (.Q (Res[43]), .D (n_0_229), .G (n_0_316));
DLH_X1 \Res_reg[44]  (.Q (Res[44]), .D (n_0_230), .G (n_0_316));
DLH_X1 \Res_reg[45]  (.Q (Res[45]), .D (n_0_231), .G (n_0_316));
DLH_X1 \Res_reg[46]  (.Q (Res[46]), .D (n_0_232), .G (n_0_316));
DLH_X1 \Res_reg[47]  (.Q (Res[47]), .D (n_0_233), .G (n_0_316));
DLH_X1 \Res_reg[48]  (.Q (Res[48]), .D (n_0_234), .G (n_0_316));
DLH_X1 \Res_reg[49]  (.Q (Res[49]), .D (n_0_235), .G (n_0_316));
DLH_X1 \Res_reg[50]  (.Q (Res[50]), .D (n_0_236), .G (n_0_316));
DLH_X1 \Res_reg[51]  (.Q (Res[51]), .D (n_0_237), .G (n_0_316));
DLH_X1 \Res_reg[52]  (.Q (Res[52]), .D (n_0_238), .G (n_0_316));
DLH_X1 \Res_reg[53]  (.Q (Res[53]), .D (n_0_239), .G (n_0_316));
DLH_X1 \Res_reg[54]  (.Q (Res[54]), .D (n_0_240), .G (n_0_316));
DLH_X1 \Res_reg[55]  (.Q (Res[55]), .D (n_0_241), .G (n_0_316));
DLH_X1 \Res_reg[56]  (.Q (Res[56]), .D (n_0_242), .G (n_0_316));
DLH_X1 \Res_reg[57]  (.Q (Res[57]), .D (n_0_243), .G (n_0_316));
DLH_X1 \Res_reg[58]  (.Q (Res[58]), .D (n_0_244), .G (n_0_316));
DLH_X1 \Res_reg[59]  (.Q (Res[59]), .D (n_0_245), .G (n_0_316));
DLH_X1 \Res_reg[60]  (.Q (Res[60]), .D (n_0_246), .G (n_0_316));
DLH_X1 \Res_reg[61]  (.Q (Res[61]), .D (n_0_247), .G (n_0_316));
DLH_X1 \Res_reg[62]  (.Q (Res[62]), .D (n_0_248), .G (n_0_316));
DLH_X1 \Res_reg[63]  (.Q (sgo__n172), .D (n_0_249), .G (n_0_316));
datapath__0_3 i_0_5 (.p_0 ({n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, 
    n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, 
    n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, 
    n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, 
    n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, 
    n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, 
    n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, uc_2})
    , .Res_imm ({\Res_imm[63] , \Res_imm[62] , \Res_imm[61] , \Res_imm[60] , \Res_imm[59] , 
    \Res_imm[58] , \Res_imm[57] , \Res_imm[56] , \Res_imm[55] , \Res_imm[54] , \Res_imm[53] , 
    \Res_imm[52] , CLOCK_opt_ipo_n666, \Res_imm[50] , \Res_imm[49] , \Res_imm[48] , 
    \Res_imm[47] , \Res_imm[46] , \Res_imm[45] , \Res_imm[44] , \Res_imm[43] , \Res_imm[42] , 
    \Res_imm[41] , \Res_imm[40] , \Res_imm[39] , \Res_imm[38] , \Res_imm[37] , \Res_imm[36] , 
    \Res_imm[35] , \Res_imm[34] , \Res_imm[33] , \Res_imm[32] , \Res_imm[31] , \Res_imm[30] , 
    \Res_imm[29] , \Res_imm[28] , \Res_imm[27] , \Res_imm[26] , \Res_imm[25] , \Res_imm[24] , 
    \Res_imm[23] , \Res_imm[22] , \Res_imm[21] , \Res_imm[20] , \Res_imm[19] , \Res_imm[18] , 
    \Res_imm[17] , \Res_imm[16] , \Res_imm[15] , \Res_imm[14] , \Res_imm[13] , \Res_imm[12] , 
    \Res_imm[11] , \Res_imm[10] , \Res_imm[9] , \Res_imm[8] , \Res_imm[7] , \Res_imm[6] , 
    \Res_imm[5] , \Res_imm[4] , \Res_imm[3] , \Res_imm[2] , \Res_imm[1] , \Res_imm[0] })
    , .opt_ipoPP_2 (\Res_imm[41] ), .opt_ipoPP_6 (\Res_imm[57] ), .opt_ipoPP_7 (\Res_imm[52] ));
datapath__0_2 i_0_4 (.Res_imm ({\Res_imm[63] , \Res_imm[62] , \Res_imm[61] , \Res_imm[60] , 
    \Res_imm[59] , \Res_imm[58] , \Res_imm[57] , \Res_imm[56] , \Res_imm[55] , \Res_imm[54] , 
    \Res_imm[53] , \Res_imm[52] , \Res_imm[51] , \Res_imm[50] , \Res_imm[49] , \Res_imm[48] , 
    \Res_imm[47] , \Res_imm[46] , \Res_imm[45] , \Res_imm[44] , \Res_imm[43] , \Res_imm[42] , 
    \Res_imm[41] , \Res_imm[40] , \Res_imm[39] , \Res_imm[38] , \Res_imm[37] , \Res_imm[36] , 
    \Res_imm[35] , \Res_imm[34] , \Res_imm[33] , \Res_imm[32] , \Res_imm[31] , \Res_imm[30] , 
    \Res_imm[29] , \Res_imm[28] , \Res_imm[27] , \Res_imm[26] , \Res_imm[25] , \Res_imm[24] , 
    \Res_imm[23] , \Res_imm[22] , \Res_imm[21] , \Res_imm[20] , \Res_imm[19] , \Res_imm[18] , 
    \Res_imm[17] , \Res_imm[16] , \Res_imm[15] , \Res_imm[14] , \Res_imm[13] , \Res_imm[12] , 
    \Res_imm[11] , \Res_imm[10] , \Res_imm[9] , \Res_imm[8] , \Res_imm[7] , \Res_imm[6] , 
    \Res_imm[5] , \Res_imm[4] , \Res_imm[3] , \Res_imm[2] , \Res_imm[1] , \Res_imm[0] })
    , .A_imm ({CLOCK_opt_ipo_n667, drc_ipo_n133, \A_imm[29] , \A_imm[28] , drc_ipo_n132, 
    drc_ipo_n149, \A_imm[25] , \A_imm[24] , drc_ipo_n148, drc_ipo_n153, drc_ipo_n147, 
    drc_ipo_n146, drc_ipo_n145, drc_ipo_n144, \A_imm[17] , drc_ipo_n169, drc_ipo_n143, 
    drc_ipo_n152, drc_ipo_n151, drc_ipo_n162, drc_ipo_n142, drc_ipo_n126, drc_ipo_n141, 
    drc_ipo_n161, drc_ipo_n157, drc_ipo_n156, drc_ipo_n155, drc_ipo_n171, drc_ipo_n160, 
    drc_ipo_n163, \A_imm[1] , drc_ipo_n164}), .B_imm ({\B_imm[31] , drc_ipo_n131, 
    \B_imm[29] , \B_imm[28] , \B_imm[27] , \B_imm[26] , \B_imm[25] , CLOCK_opt_ipo_n679, 
    drc_ipo_n140, drc_ipo_n139, drc_ipo_n130, drc_ipo_n138, drc_ipo_n137, CLOCK_opt_ipo_n662, 
    \B_imm[17] , drc_ipo_n168, drc_ipo_n129, drc_ipo_n128, drc_ipo_n136, drc_ipo_n135, 
    drc_ipo_n150, drc_ipo_n170, drc_ipo_n127, drc_ipo_n134, drc_ipo_n154, drc_ipo_n159, 
    \B_imm[5] , drc_ipo_n158, \B_imm[3] , CLOCK_opt_ipo_n727, \B_imm[1] , drc_ipo_n166}), .opt_ipoPP_0 (CLOCK_opt_ipo_n668));
datapath__0_0 i_0_2 (.p_0 ({n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, 
    n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, 
    n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, 
    n_0_35, n_0_34, n_0_33, n_0_32, uc_1}), .A_in ({drc_ipo_n165, n_0_156, n_0_157, 
    n_0_158, n_0_159, n_0_160, n_0_161, n_0_162, n_0_163, n_0_164, n_0_165, n_0_166, 
    n_0_167, n_0_168, n_0_169, n_0_170, n_0_171, n_0_172, n_0_173, n_0_174, n_0_175, 
    n_0_176, n_0_177, CLOCK_opt_ipo_n661, n_0_179, n_0_180, n_0_181, n_0_182, n_0_183, 
    n_0_184, n_0_185, drc_ipo_n164}), .opt_ipoPP_0 (CLOCK_opt_ipo_n660));
datapath i_0_0 (.p_0 ({n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, 
    n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, 
    n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, 
    n_0_2, n_0_1, uc_0}), .B_in ({drc_ipo_n167, n_0_126, n_0_127, n_0_128, n_0_129, 
    n_0_130, n_0_131, n_0_132, n_0_133, n_0_134, n_0_135, n_0_136, n_0_137, n_0_138, 
    n_0_139, n_0_140, n_0_141, n_0_142, n_0_143, n_0_144, n_0_145, n_0_146, n_0_147, 
    n_0_148, n_0_149, n_0_150, n_0_151, CLOCK_opt_ipo_n664, n_0_153, n_0_154, n_0_155, 
    drc_ipo_n166}), .opt_ipoPP_0 (CLOCK_opt_ipo_n663), .opt_ipoPP_2 (CLOCK_opt_ipo_n664));
BUF_X32 drc_ipo_c127 (.Z (drc_ipo_n127), .A (\B_imm[9] ));
BUF_X32 drc_ipo_c128 (.Z (drc_ipo_n128), .A (\B_imm[14] ));
BUF_X32 drc_ipo_c129 (.Z (drc_ipo_n129), .A (\B_imm[15] ));
BUF_X8 drc_ipo_c130 (.Z (drc_ipo_n130), .A (\B_imm[21] ));
BUF_X8 hfn_ipo_c120 (.Z (hfn_ipo_n120), .A (n_0_1_63));
CLKBUF_X1 CLOCK_slh__c812 (.Z (CLOCK_slh__n1107), .A (CLOCK_slh__n1106));
BUF_X4 drc_ipo_c132 (.Z (drc_ipo_n132), .A (\A_imm[27] ));
BUF_X4 drc_ipo_c149 (.Z (drc_ipo_n149), .A (\A_imm[26] ));
BUF_X32 drc_ipo_c133 (.Z (drc_ipo_n133), .A (\A_imm[30] ));
BUF_X4 drc_ipo_c131 (.Z (drc_ipo_n131), .A (\B_imm[30] ));
INV_X8 sgo__c240 (.ZN (\B_imm[17] ), .A (sgo__n220));
BUF_X4 drc_ipo_c169 (.Z (drc_ipo_n169), .A (\A_imm[16] ));
BUF_X8 drc_ipo_c168 (.Z (drc_ipo_n168), .A (\B_imm[16] ));
BUF_X4 drc_ipo_c163 (.Z (drc_ipo_n163), .A (\A_imm[2] ));
BUF_X16 drc_ipo_c159 (.Z (drc_ipo_n159), .A (\B_imm[6] ));
BUF_X32 drc_ipo_c135 (.Z (drc_ipo_n135), .A (\B_imm[12] ));
BUF_X32 drc_ipo_c134 (.Z (drc_ipo_n134), .A (\B_imm[8] ));
BUF_X16 sgo__c178 (.Z (\A_imm[17] ), .A (sgo__n175));
BUF_X4 drc_ipo_c171 (.Z (drc_ipo_n171), .A (\A_imm[4] ));
BUF_X4 drc_ipo_c170 (.Z (drc_ipo_n170), .A (\B_imm[10] ));
BUF_X16 drc_ipo_c165 (.Z (drc_ipo_n165), .A (A_in));
BUF_X8 drc_ipo_c164 (.Z (drc_ipo_n164), .A (n_0_0));
BUF_X4 drc_ipo_c162 (.Z (drc_ipo_n162), .A (\A_imm[12] ));
BUF_X4 drc_ipo_c161 (.Z (drc_ipo_n161), .A (\A_imm[8] ));
BUF_X4 drc_ipo_c160 (.Z (drc_ipo_n160), .A (\A_imm[3] ));
BUF_X4 drc_ipo_c150 (.Z (drc_ipo_n150), .A (\B_imm[11] ));
BUF_X16 drc_ipo_c148 (.Z (drc_ipo_n148), .A (\A_imm[23] ));
BUF_X4 drc_ipo_c144 (.Z (drc_ipo_n144), .A (\A_imm[18] ));
BUF_X8 drc_ipo_c142 (.Z (drc_ipo_n142), .A (\A_imm[11] ));
BUF_X8 drc_ipo_c141 (.Z (drc_ipo_n141), .A (\A_imm[9] ));
BUF_X4 drc_ipo_c140 (.Z (drc_ipo_n140), .A (\B_imm[23] ));
BUF_X16 drc_ipo_c139 (.Z (drc_ipo_n139), .A (\B_imm[22] ));
BUF_X4 drc_ipo_c138 (.Z (drc_ipo_n138), .A (\B_imm[20] ));
BUF_X16 drc_ipo_c136 (.Z (drc_ipo_n136), .A (\B_imm[13] ));
BUF_X4 sgo__c172 (.Z (CLOCK_sgo_n781), .A (sgo__n172));
BUF_X16 drc_ipo_c167 (.Z (drc_ipo_n167), .A (B_in));
BUF_X8 drc_ipo_c166 (.Z (drc_ipo_n166), .A (n_0_288));
BUF_X4 drc_ipo_c146 (.Z (drc_ipo_n146), .A (\A_imm[20] ));
BUF_X8 drc_ipo_c145 (.Z (drc_ipo_n145), .A (\A_imm[19] ));
BUF_X8 drc_ipo_c143 (.Z (drc_ipo_n143), .A (\A_imm[15] ));
BUF_X8 drc_ipo_c137 (.Z (drc_ipo_n137), .A (\B_imm[19] ));
INV_X1 sgo__c257 (.ZN (sgo__n238), .A (sgo__n237));
INV_X2 sgo__c239 (.ZN (sgo__n220), .A (sgo__n219));
BUF_X32 drc_ipo_c154 (.Z (drc_ipo_n154), .A (\B_imm[7] ));
BUF_X4 drc_ipo_c153 (.Z (drc_ipo_n153), .A (\A_imm[22] ));
BUF_X8 drc_ipo_c152 (.Z (drc_ipo_n152), .A (\A_imm[14] ));
INV_X8 sgo__c258 (.ZN (\B_imm[3] ), .A (sgo__n238));
BUF_X4 drc_ipo_c156 (.Z (drc_ipo_n156), .A (\A_imm[6] ));
BUF_X4 drc_ipo_c155 (.Z (drc_ipo_n155), .A (\A_imm[5] ));
BUF_X4 drc_ipo_c151 (.Z (drc_ipo_n151), .A (\A_imm[13] ));
BUF_X8 drc_ipo_c147 (.Z (drc_ipo_n147), .A (\A_imm[21] ));
INV_X1 sgo__sro_c185 (.ZN (sgo__sro_n182), .A (\Res_imm[46] ));
BUF_X8 drc_ipo_c157 (.Z (drc_ipo_n157), .A (\A_imm[7] ));
INV_X1 sgo__sro_c186 (.ZN (sgo__sro_n181), .A (\Res_imm[45] ));
BUF_X16 drc_ipo_c158 (.Z (drc_ipo_n158), .A (\B_imm[4] ));
BUF_X16 drc_ipo_c126 (.Z (drc_ipo_n126), .A (\A_imm[10] ));
BUF_X2 hfn_ipo_c125 (.Z (hfn_ipo_n125), .A (n_0_1_89));
CLKBUF_X1 CLOCK_slh__c759 (.Z (CLOCK_slh__n1057), .A (enable));
BUF_X16 hfn_ipo_c123 (.Z (hfn_ipo_n123), .A (n_0_1_64));
NAND2_X1 sgo__sro_c187 (.ZN (sgo__sro_n180), .A1 (sgo__sro_n181), .A2 (sgo__sro_n182));
NOR3_X1 sgo__sro_c188 (.ZN (sgo__sro_n179), .A1 (sgo__sro_n180), .A2 (\Res_imm[47] ), .A3 (\Res_imm[40] ));
INV_X4 sgo__c300 (.ZN (\A_imm[25] ), .A (sgo__n270));
NOR2_X1 sgo__sro_c269 (.ZN (sgo__sro_n248), .A1 (\Res_imm[60] ), .A2 (\Res_imm[59] ));
NOR2_X1 sgo__sro_c270 (.ZN (sgo__sro_n247), .A1 (\Res_imm[61] ), .A2 (\Res_imm[58] ));
AND2_X1 sgo__sro_c271 (.ZN (sgo__sro_n246), .A1 (sgo__sro_n247), .A2 (sgo__sro_n248));
INV_X16 sgo__c304 (.ZN (\B_imm[26] ), .A (sgo__n274));
INV_X1 sgo__c331 (.ZN (sgo__n292), .A (sgo__n291));
NOR2_X1 sgo__sro_c282 (.ZN (sgo__sro_n258), .A1 (\Res_imm[54] ), .A2 (\Res_imm[49] ));
INV_X4 sgo__c352 (.ZN (\B_imm[5] ), .A (sgo__n308));
INV_X1 sgo__sro_c221 (.ZN (sgo__sro_n207), .A (n_0_1_72));
INV_X1 sgo__sro_c222 (.ZN (sgo__sro_n206), .A (n_0_1_67));
NAND2_X1 sgo__sro_c223 (.ZN (sgo__sro_n205), .A1 (sgo__sro_n206), .A2 (sgo__sro_n207));
NOR2_X2 sgo__sro_c224 (.ZN (sgo__sro_n204), .A1 (n_0_1_77), .A2 (sgo__sro_n205));
NAND2_X2 sgo__sro_c225 (.ZN (n_0_1_66), .A1 (n_0_1_82), .A2 (sgo__sro_n204));
AND2_X2 sgo__sro_c284 (.ZN (sgo__sro_n256), .A1 (sgo__sro_n257), .A2 (sgo__sro_n258));
AND4_X2 sgo__c293 (.ZN (n_0_1_82), .A1 (n_0_1_84), .A2 (sgo__sro_n256), .A3 (n_0_1_85), .A4 (sgo__sro_n246));
NOR2_X4 sgo__c361 (.ZN (opt_ipo_n598), .A1 (CLOCK_sgo_n781), .A2 (drc_ipo_n165));
CLKBUF_X1 CLOCK_slh__c783 (.Z (CLOCK_slh__n1078), .A (CLOCK_slh__n1077));
INV_X4 slo__c381 (.ZN (\B_imm[28] ), .A (slo__n361));
INV_X1 slo__c386 (.ZN (slo__n367), .A (slo__n366));
INV_X4 slo__c387 (.ZN (\A_imm[28] ), .A (slo__n367));
INV_X1 slo__c403 (.ZN (slo__n384), .A (slo__n383));
INV_X4 slo__c404 (.ZN (\B_imm[25] ), .A (slo__n384));
BUF_X4 CLOCK_sgo__L1_c639 (.Z (Res[63]), .A (CLOCK_sgo_n781));
INV_X2 CLOCK_opt_ipo_c529 (.ZN (CLOCK_opt_ipo_n651), .A (n_0_1_6));
INV_X2 CLOCK_opt_ipo_c527 (.ZN (CLOCK_opt_ipo_n649), .A (n_0_1_8));
CLKBUF_X1 CLOCK_slh__c765 (.Z (CLOCK_slh__n1067), .A (CLOCK_slh__n1059));
CLKBUF_X1 CLOCK_slh__c793 (.Z (CLOCK_slh__n1088), .A (CLOCK_slh__n1087));
CLKBUF_X1 CLOCK_slh__c795 (.Z (CLOCK_slh__n1093), .A (CLOCK_slh__n1089));
CLKBUF_X1 CLOCK_slh__c794 (.Z (CLOCK_slh__n1089), .A (CLOCK_slh__n1088));
INV_X2 CLOCK_opt_ipo_c539 (.ZN (CLOCK_opt_ipo_n661), .A (n_0_178));
INV_X1 CLOCK_opt_ipo_c538 (.ZN (CLOCK_opt_ipo_n660), .A (CLOCK_opt_ipo_n661));
INV_X1 CLOCK_opt_ipo_c541 (.ZN (CLOCK_opt_ipo_n663), .A (CLOCK_opt_ipo_n664));
BUF_X8 CLOCK_opt_ipo_c540 (.Z (CLOCK_opt_ipo_n662), .A (\B_imm[18] ));
CLKBUF_X1 CLOCK_slh__c773 (.Z (CLOCK_slh__n1068), .A (CLOCK_slh__n1067));
INV_X4 CLOCK_opt_ipo_c542 (.ZN (CLOCK_opt_ipo_n664), .A (n_0_152));
BUF_X8 CLOCK_opt_ipo_c545 (.Z (CLOCK_opt_ipo_n667), .A (\A_imm[31] ));
INV_X4 CLOCK_opt_ipo_c544 (.ZN (CLOCK_opt_ipo_n666), .A (\Res_imm[51] ));
CLKBUF_X1 CLOCK_slh__c764 (.Z (CLOCK_slh__n1059), .A (CLOCK_slh__n1058));
CLKBUF_X2 CLOCK_opt_ipo_c546 (.Z (CLOCK_opt_ipo_n668), .A (\A_imm[31] ));
CLKBUF_X1 CLOCK_slh__c800 (.Z (CLOCK_slh__n1095), .A (CLOCK_slh__n1094));
CLKBUF_X1 CLOCK_slh__c799 (.Z (CLOCK_slh__n1094), .A (CLOCK_slh__n1093));
CLKBUF_X1 CLOCK_slh__c801 (.Z (CLOCK_slh__n1099), .A (CLOCK_slh__n1095));
CLKBUF_X1 CLOCK_slh__c763 (.Z (CLOCK_slh__n1058), .A (CLOCK_slh__n1057));
BUF_X8 CLOCK_opt_ipo_c557 (.Z (CLOCK_opt_ipo_n679), .A (\B_imm[24] ));
CLKBUF_X1 CLOCK_slh__c805 (.Z (CLOCK_slh__n1100), .A (CLOCK_slh__n1099));
CLKBUF_X1 CLOCK_slh__c807 (.Z (CLOCK_slh__n1105), .A (CLOCK_slh__n1101));
CLKBUF_X1 CLOCK_slh__c806 (.Z (CLOCK_slh__n1101), .A (CLOCK_slh__n1100));
BUF_X16 CLOCK_opt_ipo_c567 (.Z (CLOCK_opt_ipo_n697), .A (n_0_1_64));
INV_X2 CLOCK_opt_ipo_c565 (.ZN (CLOCK_opt_ipo_n695), .A (n_0_1_12));
INV_X2 CLOCK_opt_ipo_c571 (.ZN (CLOCK_opt_ipo_n701), .A (n_0_1_0));
INV_X2 CLOCK_opt_ipo_c569 (.ZN (CLOCK_opt_ipo_n699), .A (n_0_1_13));
INV_X2 CLOCK_opt_ipo_c575 (.ZN (CLOCK_opt_ipo_n705), .A (n_0_1_2));
INV_X2 CLOCK_opt_ipo_c573 (.ZN (CLOCK_opt_ipo_n703), .A (n_0_1_1));
INV_X2 opt_ipo_c504 (.ZN (OVF), .A (opt_ipo_n598));
CLKBUF_X1 CLOCK_slh__c774 (.Z (CLOCK_slh__n1069), .A (CLOCK_slh__n1068));
CLKBUF_X1 CLOCK_slh__c775 (.Z (CLOCK_slh__n1077), .A (CLOCK_slh__n1069));
BUF_X8 CLOCK_opt_ipo_c597 (.Z (CLOCK_opt_ipo_n727), .A (\B_imm[2] ));

endmodule //VM


