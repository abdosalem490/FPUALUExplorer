/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 16 22:57:54 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2030762560 */

module datapath(B, p_0);
   input [31:0]B;
   output [31:0]p_0;

   XOR2_X1 i_0 (.A(B[1]), .B(B[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(B[2]), .B1(B[1]), .B2(B[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(B[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(B[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(B[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(B[6]), .B1(n_27), .B2(B[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(B[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(B[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(B[9]), .B1(n_25), .B2(B[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(B[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(B[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(B[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(B[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(B[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(B[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(B[16]), .B1(n_19), .B2(B[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(B[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(B[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(B[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(B[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(B[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(B[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(B[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(B[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(B[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(B[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(B[27]), .B1(n_9), .B2(B[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(B[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(B[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(B[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(B[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(B[28]), .A3(B[29]), .A4(B[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(B[28]), .A3(B[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(B[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(B[26]), .A3(B[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(B[23]), .A3(B[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(B[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(B[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(B[18]), .A3(B[19]), .A4(B[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(B[18]), .A3(B[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(B[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(B[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(B[15]), .A3(B[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(B[12]), .A3(B[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(B[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(B[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(B[8]), .A3(B[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(B[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(B[5]), .A3(B[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(B[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(B[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(B[2]), .A2(B[1]), .A3(B[0]), .ZN(n_29));
   INV_X1 i_61 (.A(B[11]), .ZN(n_30));
   INV_X1 i_62 (.A(B[14]), .ZN(n_31));
   INV_X1 i_63 (.A(B[21]), .ZN(n_32));
   INV_X1 i_64 (.A(B[25]), .ZN(n_33));
endmodule

module datapath__0_0(A, p_0);
   input [31:0]A;
   output [31:0]p_0;

   XOR2_X1 i_0 (.A(A[1]), .B(A[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(A[2]), .B1(A[1]), .B2(A[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(A[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(A[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(A[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(A[6]), .B1(n_27), .B2(A[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(A[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(A[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(A[9]), .B1(n_25), .B2(A[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(A[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(A[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(A[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(A[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(A[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(A[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(A[16]), .B1(n_19), .B2(A[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(A[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(A[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(A[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(A[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(A[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(A[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(A[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(A[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(A[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(A[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(A[27]), .B1(n_9), .B2(A[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(A[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(A[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(A[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(A[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(A[28]), .A3(A[29]), .A4(A[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(A[28]), .A3(A[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(A[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(A[26]), .A3(A[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(A[23]), .A3(A[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(A[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(A[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(A[18]), .A3(A[19]), .A4(A[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(A[18]), .A3(A[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(A[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(A[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(A[15]), .A3(A[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(A[12]), .A3(A[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(A[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(A[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(A[8]), .A3(A[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(A[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(A[5]), .A3(A[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(A[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(A[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(A[2]), .A2(A[1]), .A3(A[0]), .ZN(n_29));
   INV_X1 i_61 (.A(A[11]), .ZN(n_30));
   INV_X1 i_62 (.A(A[14]), .ZN(n_31));
   INV_X1 i_63 (.A(A[21]), .ZN(n_32));
   INV_X1 i_64 (.A(A[25]), .ZN(n_33));
endmodule

module datapath__0_18(p_0, p_1);
   input [63:0]p_0;
   output [63:0]p_1;

   XOR2_X1 i_0 (.A(p_0[1]), .B(p_0[0]), .Z(p_1[1]));
   AND2_X1 i_1 (.A1(n_61), .A2(n_0), .ZN(p_1[2]));
   OAI21_X1 i_2 (.A(p_0[2]), .B1(p_0[1]), .B2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_0[3]), .B(n_61), .Z(p_1[3]));
   XOR2_X1 i_4 (.A(p_0[4]), .B(n_60), .Z(p_1[4]));
   XOR2_X1 i_5 (.A(p_0[5]), .B(n_59), .Z(p_1[5]));
   AND2_X1 i_6 (.A1(n_58), .A2(n_1), .ZN(p_1[6]));
   OAI21_X1 i_7 (.A(p_0[6]), .B1(n_59), .B2(p_0[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_0[7]), .B(n_58), .Z(p_1[7]));
   XOR2_X1 i_9 (.A(p_0[8]), .B(n_57), .Z(p_1[8]));
   AND2_X1 i_10 (.A1(n_56), .A2(n_2), .ZN(p_1[9]));
   OAI21_X1 i_11 (.A(p_0[9]), .B1(n_57), .B2(p_0[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_0[10]), .B(n_56), .Z(p_1[10]));
   XNOR2_X1 i_13 (.A(p_0[11]), .B(n_55), .ZN(p_1[11]));
   XOR2_X1 i_14 (.A(p_0[12]), .B(n_54), .Z(p_1[12]));
   XNOR2_X1 i_15 (.A(p_0[13]), .B(n_53), .ZN(p_1[13]));
   XOR2_X1 i_16 (.A(p_0[14]), .B(n_52), .Z(p_1[14]));
   AND2_X1 i_17 (.A1(n_51), .A2(n_3), .ZN(p_1[15]));
   OAI21_X1 i_18 (.A(p_0[15]), .B1(n_52), .B2(p_0[14]), .ZN(n_3));
   XOR2_X1 i_19 (.A(p_0[16]), .B(n_51), .Z(p_1[16]));
   XOR2_X1 i_20 (.A(p_0[17]), .B(n_50), .Z(p_1[17]));
   XOR2_X1 i_21 (.A(p_0[18]), .B(n_49), .Z(p_1[18]));
   XNOR2_X1 i_22 (.A(p_0[19]), .B(n_48), .ZN(p_1[19]));
   XNOR2_X1 i_23 (.A(p_0[20]), .B(n_47), .ZN(p_1[20]));
   XNOR2_X1 i_24 (.A(p_0[21]), .B(n_46), .ZN(p_1[21]));
   XOR2_X1 i_25 (.A(p_0[22]), .B(n_45), .Z(p_1[22]));
   XOR2_X1 i_26 (.A(p_0[23]), .B(n_44), .Z(p_1[23]));
   XNOR2_X1 i_27 (.A(p_0[24]), .B(n_43), .ZN(p_1[24]));
   XNOR2_X1 i_28 (.A(p_0[25]), .B(n_42), .ZN(p_1[25]));
   XNOR2_X1 i_29 (.A(p_0[26]), .B(n_41), .ZN(p_1[26]));
   XOR2_X1 i_30 (.A(p_0[27]), .B(n_40), .Z(p_1[27]));
   XOR2_X1 i_31 (.A(p_0[28]), .B(n_39), .Z(p_1[28]));
   XNOR2_X1 i_32 (.A(p_0[29]), .B(n_38), .ZN(p_1[29]));
   XNOR2_X1 i_33 (.A(p_0[30]), .B(n_37), .ZN(p_1[30]));
   XNOR2_X1 i_34 (.A(p_0[31]), .B(n_36), .ZN(p_1[31]));
   XOR2_X1 i_35 (.A(p_0[32]), .B(n_35), .Z(p_1[32]));
   XOR2_X1 i_36 (.A(p_0[33]), .B(n_34), .Z(p_1[33]));
   XNOR2_X1 i_37 (.A(p_0[34]), .B(n_33), .ZN(p_1[34]));
   XNOR2_X1 i_38 (.A(p_0[35]), .B(n_32), .ZN(p_1[35]));
   XNOR2_X1 i_39 (.A(p_0[36]), .B(n_31), .ZN(p_1[36]));
   XOR2_X1 i_40 (.A(p_0[37]), .B(n_30), .Z(p_1[37]));
   XOR2_X1 i_41 (.A(p_0[38]), .B(n_29), .Z(p_1[38]));
   XNOR2_X1 i_42 (.A(p_0[39]), .B(n_28), .ZN(p_1[39]));
   XNOR2_X1 i_43 (.A(p_0[40]), .B(n_27), .ZN(p_1[40]));
   XOR2_X1 i_44 (.A(p_0[41]), .B(n_26), .Z(p_1[41]));
   XNOR2_X1 i_45 (.A(p_0[42]), .B(n_25), .ZN(p_1[42]));
   XOR2_X1 i_46 (.A(p_0[43]), .B(n_24), .Z(p_1[43]));
   AND2_X1 i_47 (.A1(n_23), .A2(n_4), .ZN(p_1[44]));
   OAI21_X1 i_48 (.A(p_0[44]), .B1(n_24), .B2(p_0[43]), .ZN(n_4));
   XOR2_X1 i_49 (.A(p_0[45]), .B(n_23), .Z(p_1[45]));
   XOR2_X1 i_50 (.A(p_0[46]), .B(n_22), .Z(p_1[46]));
   XOR2_X1 i_51 (.A(p_0[47]), .B(n_21), .Z(p_1[47]));
   XOR2_X1 i_52 (.A(p_0[48]), .B(n_20), .Z(p_1[48]));
   XNOR2_X1 i_53 (.A(p_0[49]), .B(n_19), .ZN(p_1[49]));
   XNOR2_X1 i_54 (.A(p_0[50]), .B(n_18), .ZN(p_1[50]));
   XNOR2_X1 i_55 (.A(p_0[51]), .B(n_17), .ZN(p_1[51]));
   XOR2_X1 i_56 (.A(p_0[52]), .B(n_16), .Z(p_1[52]));
   XNOR2_X1 i_57 (.A(p_0[53]), .B(n_15), .ZN(p_1[53]));
   XNOR2_X1 i_58 (.A(p_0[54]), .B(n_14), .ZN(p_1[54]));
   XNOR2_X1 i_59 (.A(p_0[55]), .B(n_13), .ZN(p_1[55]));
   XOR2_X1 i_60 (.A(p_0[56]), .B(n_12), .Z(p_1[56]));
   AND2_X1 i_61 (.A1(n_11), .A2(n_5), .ZN(p_1[57]));
   OAI21_X1 i_62 (.A(p_0[57]), .B1(n_12), .B2(p_0[56]), .ZN(n_5));
   XOR2_X1 i_63 (.A(p_0[58]), .B(n_11), .Z(p_1[58]));
   XNOR2_X1 i_64 (.A(p_0[59]), .B(n_10), .ZN(p_1[59]));
   XNOR2_X1 i_65 (.A(p_0[60]), .B(n_9), .ZN(p_1[60]));
   XOR2_X1 i_66 (.A(p_0[61]), .B(n_8), .Z(p_1[61]));
   XNOR2_X1 i_67 (.A(p_0[62]), .B(n_7), .ZN(p_1[62]));
   XNOR2_X1 i_68 (.A(p_0[63]), .B(n_6), .ZN(p_1[63]));
   NOR3_X1 i_69 (.A1(n_8), .A2(p_0[61]), .A3(p_0[62]), .ZN(n_6));
   NOR2_X1 i_70 (.A1(n_8), .A2(p_0[61]), .ZN(n_7));
   NAND2_X1 i_71 (.A1(n_9), .A2(n_72), .ZN(n_8));
   NOR3_X1 i_72 (.A1(n_11), .A2(p_0[58]), .A3(p_0[59]), .ZN(n_9));
   NOR2_X1 i_73 (.A1(n_11), .A2(p_0[58]), .ZN(n_10));
   OR3_X1 i_74 (.A1(n_12), .A2(p_0[56]), .A3(p_0[57]), .ZN(n_11));
   NAND2_X1 i_75 (.A1(n_13), .A2(n_71), .ZN(n_12));
   NOR4_X1 i_76 (.A1(n_16), .A2(p_0[52]), .A3(p_0[53]), .A4(p_0[54]), .ZN(n_13));
   NOR3_X1 i_77 (.A1(n_16), .A2(p_0[52]), .A3(p_0[53]), .ZN(n_14));
   NOR2_X1 i_78 (.A1(n_16), .A2(p_0[52]), .ZN(n_15));
   NAND2_X1 i_79 (.A1(n_17), .A2(n_70), .ZN(n_16));
   NOR4_X1 i_80 (.A1(n_20), .A2(p_0[48]), .A3(p_0[49]), .A4(p_0[50]), .ZN(n_17));
   NOR3_X1 i_81 (.A1(n_20), .A2(p_0[48]), .A3(p_0[49]), .ZN(n_18));
   NOR2_X1 i_82 (.A1(n_20), .A2(p_0[48]), .ZN(n_19));
   OR2_X1 i_83 (.A1(n_21), .A2(p_0[47]), .ZN(n_20));
   OR2_X1 i_84 (.A1(n_22), .A2(p_0[46]), .ZN(n_21));
   OR2_X1 i_85 (.A1(n_23), .A2(p_0[45]), .ZN(n_22));
   OR3_X1 i_86 (.A1(n_24), .A2(p_0[43]), .A3(p_0[44]), .ZN(n_23));
   NAND2_X1 i_87 (.A1(n_25), .A2(n_69), .ZN(n_24));
   NOR2_X1 i_88 (.A1(n_26), .A2(p_0[41]), .ZN(n_25));
   NAND2_X1 i_89 (.A1(n_27), .A2(n_68), .ZN(n_26));
   NOR3_X1 i_90 (.A1(n_29), .A2(p_0[38]), .A3(p_0[39]), .ZN(n_27));
   NOR2_X1 i_91 (.A1(n_29), .A2(p_0[38]), .ZN(n_28));
   OR2_X1 i_92 (.A1(n_30), .A2(p_0[37]), .ZN(n_29));
   NAND2_X1 i_93 (.A1(n_31), .A2(n_67), .ZN(n_30));
   NOR4_X1 i_94 (.A1(n_34), .A2(p_0[33]), .A3(p_0[34]), .A4(p_0[35]), .ZN(n_31));
   NOR3_X1 i_95 (.A1(n_34), .A2(p_0[33]), .A3(p_0[34]), .ZN(n_32));
   NOR2_X1 i_96 (.A1(n_34), .A2(p_0[33]), .ZN(n_33));
   OR2_X1 i_97 (.A1(n_35), .A2(p_0[32]), .ZN(n_34));
   NAND2_X1 i_98 (.A1(n_36), .A2(n_66), .ZN(n_35));
   NOR4_X1 i_99 (.A1(n_39), .A2(p_0[28]), .A3(p_0[29]), .A4(p_0[30]), .ZN(n_36));
   NOR3_X1 i_100 (.A1(n_39), .A2(p_0[28]), .A3(p_0[29]), .ZN(n_37));
   NOR2_X1 i_101 (.A1(n_39), .A2(p_0[28]), .ZN(n_38));
   OR2_X1 i_102 (.A1(n_40), .A2(p_0[27]), .ZN(n_39));
   NAND2_X1 i_103 (.A1(n_41), .A2(n_65), .ZN(n_40));
   NOR4_X1 i_104 (.A1(n_44), .A2(p_0[23]), .A3(p_0[24]), .A4(p_0[25]), .ZN(n_41));
   NOR3_X1 i_105 (.A1(n_44), .A2(p_0[23]), .A3(p_0[24]), .ZN(n_42));
   NOR2_X1 i_106 (.A1(n_44), .A2(p_0[23]), .ZN(n_43));
   OR2_X1 i_107 (.A1(n_45), .A2(p_0[22]), .ZN(n_44));
   NAND2_X1 i_108 (.A1(n_46), .A2(n_64), .ZN(n_45));
   NOR4_X1 i_109 (.A1(n_49), .A2(p_0[18]), .A3(p_0[19]), .A4(p_0[20]), .ZN(n_46));
   NOR3_X1 i_110 (.A1(n_49), .A2(p_0[18]), .A3(p_0[19]), .ZN(n_47));
   NOR2_X1 i_111 (.A1(n_49), .A2(p_0[18]), .ZN(n_48));
   OR2_X1 i_112 (.A1(n_50), .A2(p_0[17]), .ZN(n_49));
   OR2_X1 i_113 (.A1(n_51), .A2(p_0[16]), .ZN(n_50));
   OR3_X1 i_114 (.A1(n_52), .A2(p_0[14]), .A3(p_0[15]), .ZN(n_51));
   NAND2_X1 i_115 (.A1(n_53), .A2(n_63), .ZN(n_52));
   NOR2_X1 i_116 (.A1(n_54), .A2(p_0[12]), .ZN(n_53));
   NAND2_X1 i_117 (.A1(n_55), .A2(n_62), .ZN(n_54));
   NOR2_X1 i_118 (.A1(n_56), .A2(p_0[10]), .ZN(n_55));
   OR3_X1 i_119 (.A1(n_57), .A2(p_0[8]), .A3(p_0[9]), .ZN(n_56));
   OR2_X1 i_120 (.A1(n_58), .A2(p_0[7]), .ZN(n_57));
   OR3_X1 i_121 (.A1(n_59), .A2(p_0[5]), .A3(p_0[6]), .ZN(n_58));
   OR2_X1 i_122 (.A1(n_60), .A2(p_0[4]), .ZN(n_59));
   OR2_X1 i_123 (.A1(n_61), .A2(p_0[3]), .ZN(n_60));
   OR3_X1 i_124 (.A1(p_0[2]), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_61));
   INV_X1 i_125 (.A(p_0[11]), .ZN(n_62));
   INV_X1 i_126 (.A(p_0[13]), .ZN(n_63));
   INV_X1 i_127 (.A(p_0[21]), .ZN(n_64));
   INV_X1 i_128 (.A(p_0[26]), .ZN(n_65));
   INV_X1 i_129 (.A(p_0[31]), .ZN(n_66));
   INV_X1 i_130 (.A(p_0[36]), .ZN(n_67));
   INV_X1 i_131 (.A(p_0[40]), .ZN(n_68));
   INV_X1 i_132 (.A(p_0[42]), .ZN(n_69));
   INV_X1 i_133 (.A(p_0[51]), .ZN(n_70));
   INV_X1 i_134 (.A(p_0[55]), .ZN(n_71));
   INV_X1 i_135 (.A(p_0[60]), .ZN(n_72));
endmodule

module datapath__0_5(multiplier, accumulator, p_0);
   input [31:0]multiplier;
   input [31:0]accumulator;
   output [32:0]p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0[0]));
   OAI21_X1 i_1 (.A(n_146), .B1(multiplier[0]), .B2(accumulator[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_146), .B(n_1), .Z(p_0[1]));
   OAI21_X1 i_3 (.A(n_145), .B1(multiplier[1]), .B2(accumulator[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_144), .B(n_2), .ZN(p_0[2]));
   OAI21_X1 i_5 (.A(n_149), .B1(multiplier[2]), .B2(accumulator[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_143), .B(n_3), .Z(p_0[3]));
   OAI21_X1 i_7 (.A(n_150), .B1(n_179), .B2(n_176), .ZN(n_3));
   XOR2_X1 i_8 (.A(n_141), .B(n_10), .Z(p_0[4]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_0[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_0[6]));
   NOR2_X1 i_11 (.A1(n_138), .A2(n_129), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_0[7]));
   OAI22_X1 i_13 (.A1(multiplier[6]), .A2(accumulator[6]), .B1(n_129), .B2(n_7), 
      .ZN(n_5));
   AOI21_X1 i_14 (.A(n_139), .B1(multiplier[5]), .B2(accumulator[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_139), .B1(n_133), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_136), .B1(n_141), .B2(n_134), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_134), .B1(multiplier[4]), .B2(accumulator[4]), .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_140), .A2(n_131), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_127), .B(n_18), .ZN(p_0[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_0[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_0[10]));
   NOR2_X1 i_23 (.A1(n_124), .A2(n_115), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_0[11]));
   OAI22_X1 i_25 (.A1(multiplier[10]), .A2(accumulator[10]), .B1(n_115), 
      .B2(n_15), .ZN(n_13));
   AOI21_X1 i_26 (.A(n_125), .B1(multiplier[9]), .B2(accumulator[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_125), .B1(n_119), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_122), .B1(n_127), .B2(n_120), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_122), .B1(multiplier[8]), .B2(accumulator[8]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_126), .A2(n_117), .ZN(n_19));
   XOR2_X1 i_32 (.A(n_113), .B(n_26), .Z(p_0[12]));
   XOR2_X1 i_33 (.A(n_25), .B(n_22), .Z(p_0[13]));
   XOR2_X1 i_34 (.A(n_23), .B(n_20), .Z(p_0[14]));
   NOR2_X1 i_35 (.A1(n_110), .A2(n_101), .ZN(n_20));
   XNOR2_X1 i_36 (.A(n_27), .B(n_21), .ZN(p_0[15]));
   OAI22_X1 i_37 (.A1(multiplier[14]), .A2(accumulator[14]), .B1(n_101), 
      .B2(n_23), .ZN(n_21));
   AOI21_X1 i_38 (.A(n_111), .B1(multiplier[13]), .B2(accumulator[13]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_111), .B1(n_105), .B2(n_24), .ZN(n_23));
   INV_X1 i_40 (.A(n_25), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_108), .B1(n_113), .B2(n_106), .ZN(n_25));
   OAI21_X1 i_42 (.A(n_106), .B1(multiplier[12]), .B2(accumulator[12]), .ZN(n_26));
   NOR2_X1 i_43 (.A1(n_112), .A2(n_103), .ZN(n_27));
   XOR2_X1 i_44 (.A(n_99), .B(n_34), .Z(p_0[16]));
   XOR2_X1 i_45 (.A(n_33), .B(n_30), .Z(p_0[17]));
   XOR2_X1 i_46 (.A(n_31), .B(n_28), .Z(p_0[18]));
   NOR2_X1 i_47 (.A1(n_159), .A2(n_152), .ZN(n_28));
   XNOR2_X1 i_48 (.A(n_35), .B(n_29), .ZN(p_0[19]));
   OAI21_X1 i_49 (.A(n_158), .B1(n_152), .B2(n_31), .ZN(n_29));
   NOR2_X1 i_50 (.A1(n_161), .A2(n_155), .ZN(n_30));
   INV_X1 i_51 (.A(n_32), .ZN(n_31));
   OAI21_X1 i_52 (.A(n_160), .B1(n_155), .B2(n_33), .ZN(n_32));
   AOI21_X1 i_53 (.A(n_97), .B1(n_156), .B2(n_99), .ZN(n_33));
   OAI21_X1 i_54 (.A(n_156), .B1(multiplier[16]), .B2(accumulator[16]), .ZN(n_34));
   AOI21_X1 i_55 (.A(n_162), .B1(multiplier[19]), .B2(accumulator[19]), .ZN(n_35));
   XOR2_X1 i_56 (.A(n_95), .B(n_42), .Z(p_0[20]));
   XOR2_X1 i_57 (.A(n_41), .B(n_38), .Z(p_0[21]));
   XOR2_X1 i_58 (.A(n_39), .B(n_36), .Z(p_0[22]));
   NOR2_X1 i_59 (.A1(n_85), .A2(n_68), .ZN(n_36));
   XNOR2_X1 i_60 (.A(n_43), .B(n_37), .ZN(p_0[23]));
   OAI21_X1 i_61 (.A(n_84), .B1(n_68), .B2(n_39), .ZN(n_37));
   NOR2_X1 i_62 (.A1(n_87), .A2(n_70), .ZN(n_38));
   INV_X1 i_63 (.A(n_40), .ZN(n_39));
   OAI21_X1 i_64 (.A(n_86), .B1(n_70), .B2(n_41), .ZN(n_40));
   AOI21_X1 i_65 (.A(n_82), .B1(n_95), .B2(n_72), .ZN(n_41));
   OAI21_X1 i_66 (.A(n_72), .B1(multiplier[20]), .B2(accumulator[20]), .ZN(n_42));
   AOI21_X1 i_67 (.A(n_89), .B1(multiplier[23]), .B2(accumulator[23]), .ZN(n_43));
   XNOR2_X1 i_68 (.A(n_53), .B(n_52), .ZN(p_0[24]));
   AOI22_X1 i_69 (.A1(n_51), .A2(n_48), .B1(n_50), .B2(n_49), .ZN(p_0[25]));
   XNOR2_X1 i_70 (.A(n_45), .B(n_44), .ZN(p_0[26]));
   OAI22_X1 i_71 (.A1(multiplier[25]), .A2(accumulator[25]), .B1(n_77), .B2(n_50), 
      .ZN(n_44));
   NOR2_X1 i_72 (.A1(n_92), .A2(n_74), .ZN(n_45));
   XNOR2_X1 i_73 (.A(n_54), .B(n_46), .ZN(p_0[27]));
   AOI221_X1 i_74 (.A(n_92), .B1(n_93), .B2(n_75), .C1(n_51), .C2(n_47), 
      .ZN(n_46));
   NOR2_X1 i_75 (.A1(n_74), .A2(n_48), .ZN(n_47));
   INV_X1 i_76 (.A(n_49), .ZN(n_48));
   NOR2_X1 i_77 (.A1(n_93), .A2(n_77), .ZN(n_49));
   INV_X1 i_78 (.A(n_51), .ZN(n_50));
   OAI22_X1 i_79 (.A1(multiplier[24]), .A2(accumulator[24]), .B1(n_78), .B2(n_53), 
      .ZN(n_51));
   OAI21_X1 i_80 (.A(n_79), .B1(multiplier[24]), .B2(accumulator[24]), .ZN(n_52));
   OAI21_X1 i_81 (.A(n_67), .B1(n_95), .B2(n_81), .ZN(n_53));
   OAI22_X1 i_82 (.A1(multiplier[27]), .A2(accumulator[27]), .B1(n_180), 
      .B2(n_177), .ZN(n_54));
   XOR2_X1 i_83 (.A(n_65), .B(n_63), .Z(p_0[28]));
   AOI22_X1 i_84 (.A1(n_61), .A2(n_59), .B1(n_62), .B2(n_60), .ZN(p_0[29]));
   XNOR2_X1 i_85 (.A(n_56), .B(n_55), .ZN(p_0[30]));
   OAI22_X1 i_86 (.A1(multiplier[29]), .A2(accumulator[29]), .B1(n_169), 
      .B2(n_62), .ZN(n_55));
   NOR2_X1 i_87 (.A1(n_173), .A2(n_166), .ZN(n_56));
   XNOR2_X1 i_88 (.A(n_64), .B(n_57), .ZN(p_0[31]));
   AOI221_X1 i_89 (.A(n_173), .B1(n_174), .B2(n_167), .C1(n_61), .C2(n_58), 
      .ZN(n_57));
   NOR2_X1 i_90 (.A1(n_166), .A2(n_59), .ZN(n_58));
   INV_X1 i_91 (.A(n_60), .ZN(n_59));
   NOR2_X1 i_92 (.A1(n_174), .A2(n_169), .ZN(n_60));
   INV_X1 i_93 (.A(n_62), .ZN(n_61));
   AOI21_X1 i_94 (.A(n_164), .B1(n_171), .B2(n_65), .ZN(n_62));
   OR2_X1 i_95 (.A1(n_170), .A2(n_164), .ZN(n_63));
   OAI21_X1 i_96 (.A(n_175), .B1(n_181), .B2(n_178), .ZN(n_64));
   OAI221_X1 i_97 (.A(n_165), .B1(n_172), .B2(n_168), .C1(n_163), .C2(n_65), 
      .ZN(p_0[32]));
   NOR3_X1 i_98 (.A1(n_73), .A2(n_66), .A3(n_80), .ZN(n_65));
   NOR2_X1 i_99 (.A1(n_90), .A2(n_67), .ZN(n_66));
   AOI221_X1 i_100 (.A(n_69), .B1(multiplier[23]), .B2(accumulator[23]), 
      .C1(n_88), .C2(n_68), .ZN(n_67));
   AND2_X1 i_101 (.A1(multiplier[22]), .A2(accumulator[22]), .ZN(n_68));
   AOI21_X1 i_102 (.A(n_83), .B1(n_72), .B2(n_71), .ZN(n_69));
   INV_X1 i_103 (.A(n_71), .ZN(n_70));
   NAND2_X1 i_104 (.A1(multiplier[21]), .A2(accumulator[21]), .ZN(n_71));
   NAND2_X1 i_105 (.A1(multiplier[20]), .A2(accumulator[20]), .ZN(n_72));
   OAI221_X1 i_106 (.A(n_76), .B1(n_180), .B2(n_177), .C1(n_94), .C2(n_75), 
      .ZN(n_73));
   INV_X1 i_107 (.A(n_75), .ZN(n_74));
   NAND2_X1 i_108 (.A1(multiplier[26]), .A2(accumulator[26]), .ZN(n_75));
   OAI21_X1 i_109 (.A(n_91), .B1(n_78), .B2(n_77), .ZN(n_76));
   AND2_X1 i_110 (.A1(multiplier[25]), .A2(accumulator[25]), .ZN(n_77));
   INV_X1 i_111 (.A(n_79), .ZN(n_78));
   NAND2_X1 i_112 (.A1(multiplier[24]), .A2(accumulator[24]), .ZN(n_79));
   NOR3_X1 i_113 (.A1(n_90), .A2(n_81), .A3(n_95), .ZN(n_80));
   OR2_X1 i_114 (.A1(n_83), .A2(n_82), .ZN(n_81));
   NOR2_X1 i_115 (.A1(multiplier[20]), .A2(accumulator[20]), .ZN(n_82));
   NAND3_X1 i_116 (.A1(n_88), .A2(n_84), .A3(n_86), .ZN(n_83));
   INV_X1 i_117 (.A(n_85), .ZN(n_84));
   NOR2_X1 i_118 (.A1(multiplier[22]), .A2(accumulator[22]), .ZN(n_85));
   INV_X1 i_119 (.A(n_87), .ZN(n_86));
   NOR2_X1 i_120 (.A1(multiplier[21]), .A2(accumulator[21]), .ZN(n_87));
   INV_X1 i_121 (.A(n_89), .ZN(n_88));
   NOR2_X1 i_122 (.A1(multiplier[23]), .A2(accumulator[23]), .ZN(n_89));
   OAI21_X1 i_123 (.A(n_91), .B1(multiplier[24]), .B2(accumulator[24]), .ZN(n_90));
   NOR3_X1 i_124 (.A1(n_94), .A2(n_92), .A3(n_93), .ZN(n_91));
   NOR2_X1 i_125 (.A1(multiplier[26]), .A2(accumulator[26]), .ZN(n_92));
   NOR2_X1 i_126 (.A1(multiplier[25]), .A2(accumulator[25]), .ZN(n_93));
   NOR2_X1 i_127 (.A1(multiplier[27]), .A2(accumulator[27]), .ZN(n_94));
   AOI221_X1 i_128 (.A(n_151), .B1(multiplier[19]), .B2(accumulator[19]), 
      .C1(n_98), .C2(n_96), .ZN(n_95));
   NOR2_X1 i_129 (.A1(n_157), .A2(n_97), .ZN(n_96));
   NOR2_X1 i_130 (.A1(multiplier[16]), .A2(accumulator[16]), .ZN(n_97));
   INV_X1 i_131 (.A(n_99), .ZN(n_98));
   NOR4_X1 i_132 (.A1(n_103), .A2(n_100), .A3(n_104), .A4(n_107), .ZN(n_99));
   NOR2_X1 i_133 (.A1(n_112), .A2(n_102), .ZN(n_100));
   INV_X1 i_134 (.A(n_102), .ZN(n_101));
   NAND2_X1 i_135 (.A1(multiplier[14]), .A2(accumulator[14]), .ZN(n_102));
   AND2_X1 i_136 (.A1(multiplier[15]), .A2(accumulator[15]), .ZN(n_103));
   AOI21_X1 i_137 (.A(n_109), .B1(n_106), .B2(n_105), .ZN(n_104));
   NAND2_X1 i_138 (.A1(multiplier[13]), .A2(accumulator[13]), .ZN(n_105));
   NAND2_X1 i_139 (.A1(multiplier[12]), .A2(accumulator[12]), .ZN(n_106));
   NOR3_X1 i_140 (.A1(n_109), .A2(n_108), .A3(n_113), .ZN(n_107));
   NOR2_X1 i_141 (.A1(multiplier[12]), .A2(accumulator[12]), .ZN(n_108));
   OR3_X1 i_142 (.A1(n_112), .A2(n_110), .A3(n_111), .ZN(n_109));
   NOR2_X1 i_143 (.A1(multiplier[14]), .A2(accumulator[14]), .ZN(n_110));
   NOR2_X1 i_144 (.A1(multiplier[13]), .A2(accumulator[13]), .ZN(n_111));
   NOR2_X1 i_145 (.A1(multiplier[15]), .A2(accumulator[15]), .ZN(n_112));
   NOR4_X1 i_146 (.A1(n_117), .A2(n_114), .A3(n_118), .A4(n_121), .ZN(n_113));
   NOR2_X1 i_147 (.A1(n_126), .A2(n_116), .ZN(n_114));
   INV_X1 i_148 (.A(n_116), .ZN(n_115));
   NAND2_X1 i_149 (.A1(multiplier[10]), .A2(accumulator[10]), .ZN(n_116));
   AND2_X1 i_150 (.A1(multiplier[11]), .A2(accumulator[11]), .ZN(n_117));
   AOI21_X1 i_151 (.A(n_123), .B1(n_120), .B2(n_119), .ZN(n_118));
   NAND2_X1 i_152 (.A1(multiplier[9]), .A2(accumulator[9]), .ZN(n_119));
   NAND2_X1 i_153 (.A1(multiplier[8]), .A2(accumulator[8]), .ZN(n_120));
   NOR3_X1 i_154 (.A1(n_123), .A2(n_122), .A3(n_127), .ZN(n_121));
   NOR2_X1 i_155 (.A1(multiplier[8]), .A2(accumulator[8]), .ZN(n_122));
   OR3_X1 i_156 (.A1(n_126), .A2(n_124), .A3(n_125), .ZN(n_123));
   NOR2_X1 i_157 (.A1(multiplier[10]), .A2(accumulator[10]), .ZN(n_124));
   NOR2_X1 i_158 (.A1(multiplier[9]), .A2(accumulator[9]), .ZN(n_125));
   NOR2_X1 i_159 (.A1(multiplier[11]), .A2(accumulator[11]), .ZN(n_126));
   NOR4_X1 i_160 (.A1(n_131), .A2(n_128), .A3(n_132), .A4(n_135), .ZN(n_127));
   NOR2_X1 i_161 (.A1(n_140), .A2(n_130), .ZN(n_128));
   INV_X1 i_162 (.A(n_130), .ZN(n_129));
   NAND2_X1 i_163 (.A1(multiplier[6]), .A2(accumulator[6]), .ZN(n_130));
   AND2_X1 i_164 (.A1(multiplier[7]), .A2(accumulator[7]), .ZN(n_131));
   AOI21_X1 i_165 (.A(n_137), .B1(n_134), .B2(n_133), .ZN(n_132));
   NAND2_X1 i_166 (.A1(multiplier[5]), .A2(accumulator[5]), .ZN(n_133));
   NAND2_X1 i_167 (.A1(multiplier[4]), .A2(accumulator[4]), .ZN(n_134));
   NOR3_X1 i_168 (.A1(n_137), .A2(n_136), .A3(n_141), .ZN(n_135));
   NOR2_X1 i_169 (.A1(multiplier[4]), .A2(accumulator[4]), .ZN(n_136));
   OR3_X1 i_170 (.A1(n_140), .A2(n_138), .A3(n_139), .ZN(n_137));
   NOR2_X1 i_171 (.A1(multiplier[6]), .A2(accumulator[6]), .ZN(n_138));
   NOR2_X1 i_172 (.A1(multiplier[5]), .A2(accumulator[5]), .ZN(n_139));
   NOR2_X1 i_173 (.A1(multiplier[7]), .A2(accumulator[7]), .ZN(n_140));
   NAND2_X1 i_174 (.A1(n_150), .A2(n_142), .ZN(n_141));
   OAI21_X1 i_175 (.A(n_143), .B1(n_179), .B2(n_176), .ZN(n_142));
   OAI22_X1 i_176 (.A1(multiplier[2]), .A2(accumulator[2]), .B1(n_148), .B2(
      n_144), .ZN(n_143));
   AOI21_X1 i_177 (.A(n_147), .B1(n_146), .B2(n_145), .ZN(n_144));
   NAND2_X1 i_178 (.A1(multiplier[1]), .A2(accumulator[1]), .ZN(n_145));
   NAND2_X1 i_179 (.A1(multiplier[0]), .A2(accumulator[0]), .ZN(n_146));
   NOR2_X1 i_180 (.A1(multiplier[1]), .A2(accumulator[1]), .ZN(n_147));
   INV_X1 i_181 (.A(n_149), .ZN(n_148));
   NAND2_X1 i_182 (.A1(multiplier[2]), .A2(accumulator[2]), .ZN(n_149));
   NAND2_X1 i_183 (.A1(n_179), .A2(n_176), .ZN(n_150));
   OAI22_X1 i_184 (.A1(n_157), .A2(n_154), .B1(n_162), .B2(n_153), .ZN(n_151));
   INV_X1 i_185 (.A(n_153), .ZN(n_152));
   NAND2_X1 i_186 (.A1(multiplier[18]), .A2(accumulator[18]), .ZN(n_153));
   AOI21_X1 i_187 (.A(n_155), .B1(multiplier[16]), .B2(accumulator[16]), 
      .ZN(n_154));
   AND2_X1 i_188 (.A1(multiplier[17]), .A2(accumulator[17]), .ZN(n_155));
   NAND2_X1 i_189 (.A1(multiplier[16]), .A2(accumulator[16]), .ZN(n_156));
   OAI211_X1 i_190 (.A(n_158), .B(n_160), .C1(multiplier[19]), .C2(
      accumulator[19]), .ZN(n_157));
   INV_X1 i_191 (.A(n_159), .ZN(n_158));
   NOR2_X1 i_192 (.A1(multiplier[18]), .A2(accumulator[18]), .ZN(n_159));
   INV_X1 i_193 (.A(n_161), .ZN(n_160));
   NOR2_X1 i_194 (.A1(multiplier[17]), .A2(accumulator[17]), .ZN(n_161));
   NOR2_X1 i_195 (.A1(multiplier[19]), .A2(accumulator[19]), .ZN(n_162));
   OR2_X1 i_196 (.A1(n_172), .A2(n_164), .ZN(n_163));
   NOR2_X1 i_197 (.A1(multiplier[28]), .A2(accumulator[28]), .ZN(n_164));
   AOI22_X1 i_198 (.A1(multiplier[31]), .A2(accumulator[31]), .B1(n_175), 
      .B2(n_166), .ZN(n_165));
   INV_X1 i_199 (.A(n_167), .ZN(n_166));
   NAND2_X1 i_200 (.A1(multiplier[30]), .A2(accumulator[30]), .ZN(n_167));
   NOR2_X1 i_201 (.A1(n_170), .A2(n_169), .ZN(n_168));
   AND2_X1 i_202 (.A1(multiplier[29]), .A2(accumulator[29]), .ZN(n_169));
   INV_X1 i_203 (.A(n_171), .ZN(n_170));
   NAND2_X1 i_204 (.A1(multiplier[28]), .A2(accumulator[28]), .ZN(n_171));
   OAI221_X1 i_205 (.A(n_175), .B1(multiplier[29]), .B2(accumulator[29]), 
      .C1(multiplier[30]), .C2(accumulator[30]), .ZN(n_172));
   NOR2_X1 i_206 (.A1(multiplier[30]), .A2(accumulator[30]), .ZN(n_173));
   NOR2_X1 i_207 (.A1(multiplier[29]), .A2(accumulator[29]), .ZN(n_174));
   NAND2_X1 i_208 (.A1(n_181), .A2(n_178), .ZN(n_175));
   INV_X1 i_209 (.A(accumulator[3]), .ZN(n_176));
   INV_X1 i_210 (.A(accumulator[27]), .ZN(n_177));
   INV_X1 i_211 (.A(accumulator[31]), .ZN(n_178));
   INV_X1 i_212 (.A(multiplier[3]), .ZN(n_179));
   INV_X1 i_213 (.A(multiplier[27]), .ZN(n_180));
   INV_X1 i_214 (.A(multiplier[31]), .ZN(n_181));
endmodule

module sequentialMultiplier(Res, OVF, A, B, clk, reset, enable);
   output [63:0]Res;
   output OVF;
   input [31:0]A;
   input [31:0]B;
   input clk;
   input reset;
   input enable;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire [1:0]isNeg;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire [31:0]accumulator;
   wire [31:0]multiplicand;
   wire ready;
   wire [31:0]multiplier;
   wire carry;
   wire [4:0]counter;
   wire n_0_158;
   wire n_0_159;
   wire n_0_1_0;
   wire n_0_160;
   wire n_0_161;
   wire n_0_1_1;
   wire n_0_162;
   wire n_0_1_2;
   wire n_0_163;
   wire n_0_1_3;
   wire n_0_164;
   wire n_0_1_4;
   wire n_0_1_5;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_165;
   wire n_0_1_8;
   wire n_0_166;
   wire n_0_1_9;
   wire n_0_167;
   wire n_0_1_10;
   wire n_0_168;
   wire n_0_1_11;
   wire n_0_169;
   wire n_0_1_12;
   wire n_0_170;
   wire n_0_1_13;
   wire n_0_171;
   wire n_0_1_14;
   wire n_0_172;
   wire n_0_1_15;
   wire n_0_173;
   wire n_0_1_16;
   wire n_0_174;
   wire n_0_1_17;
   wire n_0_175;
   wire n_0_1_18;
   wire n_0_176;
   wire n_0_1_19;
   wire n_0_177;
   wire n_0_1_20;
   wire n_0_178;
   wire n_0_1_21;
   wire n_0_179;
   wire n_0_1_22;
   wire n_0_180;
   wire n_0_1_23;
   wire n_0_181;
   wire n_0_1_24;
   wire n_0_182;
   wire n_0_1_25;
   wire n_0_183;
   wire n_0_1_26;
   wire n_0_184;
   wire n_0_1_27;
   wire n_0_185;
   wire n_0_1_28;
   wire n_0_186;
   wire n_0_1_29;
   wire n_0_187;
   wire n_0_1_30;
   wire n_0_188;
   wire n_0_1_31;
   wire n_0_189;
   wire n_0_1_32;
   wire n_0_190;
   wire n_0_1_33;
   wire n_0_191;
   wire n_0_1_34;
   wire n_0_192;
   wire n_0_1_35;
   wire n_0_193;
   wire n_0_1_36;
   wire n_0_194;
   wire n_0_1_37;
   wire n_0_195;
   wire n_0_1_38;
   wire n_0_196;
   wire n_0_1_39;
   wire n_0_197;
   wire n_0_1_40;
   wire n_0_1_41;
   wire n_0_1_42;
   wire n_0_198;
   wire n_0_1_43;
   wire n_0_199;
   wire n_0_1_44;
   wire n_0_200;
   wire n_0_1_45;
   wire n_0_201;
   wire n_0_1_46;
   wire n_0_202;
   wire n_0_1_47;
   wire n_0_203;
   wire n_0_1_48;
   wire n_0_204;
   wire n_0_1_49;
   wire n_0_205;
   wire n_0_1_50;
   wire n_0_206;
   wire n_0_1_51;
   wire n_0_207;
   wire n_0_1_52;
   wire n_0_208;
   wire n_0_1_53;
   wire n_0_209;
   wire n_0_1_54;
   wire n_0_210;
   wire n_0_1_55;
   wire n_0_211;
   wire n_0_1_56;
   wire n_0_212;
   wire n_0_1_57;
   wire n_0_213;
   wire n_0_1_58;
   wire n_0_214;
   wire n_0_1_59;
   wire n_0_215;
   wire n_0_1_60;
   wire n_0_216;
   wire n_0_1_61;
   wire n_0_217;
   wire n_0_1_62;
   wire n_0_218;
   wire n_0_1_63;
   wire n_0_219;
   wire n_0_1_64;
   wire n_0_220;
   wire n_0_1_65;
   wire n_0_221;
   wire n_0_1_66;
   wire n_0_222;
   wire n_0_1_67;
   wire n_0_223;
   wire n_0_1_68;
   wire n_0_224;
   wire n_0_1_69;
   wire n_0_225;
   wire n_0_1_70;
   wire n_0_226;
   wire n_0_1_71;
   wire n_0_227;
   wire n_0_1_72;
   wire n_0_228;
   wire n_0_1_73;
   wire n_0_1_74;
   wire n_0_229;
   wire n_0_1_75;
   wire n_0_1_76;
   wire n_0_1_77;
   wire n_0_1_78;
   wire n_0_230;
   wire n_0_231;
   wire n_0_1_79;
   wire n_0_232;
   wire n_0_1_80;
   wire n_0_233;
   wire n_0_1_81;
   wire n_0_234;
   wire n_0_1_82;
   wire n_0_235;
   wire n_0_1_83;
   wire n_0_236;
   wire n_0_1_84;
   wire n_0_237;
   wire n_0_1_85;
   wire n_0_238;
   wire n_0_1_86;
   wire n_0_239;
   wire n_0_1_87;
   wire n_0_240;
   wire n_0_1_88;
   wire n_0_241;
   wire n_0_1_89;
   wire n_0_242;
   wire n_0_1_90;
   wire n_0_243;
   wire n_0_1_91;
   wire n_0_244;
   wire n_0_1_92;
   wire n_0_245;
   wire n_0_1_93;
   wire n_0_246;
   wire n_0_1_94;
   wire n_0_247;
   wire n_0_1_95;
   wire n_0_248;
   wire n_0_1_96;
   wire n_0_249;
   wire n_0_1_97;
   wire n_0_250;
   wire n_0_1_98;
   wire n_0_251;
   wire n_0_1_99;
   wire n_0_252;
   wire n_0_1_100;
   wire n_0_253;
   wire n_0_1_101;
   wire n_0_254;
   wire n_0_1_102;
   wire n_0_255;
   wire n_0_1_103;
   wire n_0_256;
   wire n_0_1_104;
   wire n_0_257;
   wire n_0_1_105;
   wire n_0_258;
   wire n_0_1_106;
   wire n_0_259;
   wire n_0_1_107;
   wire n_0_260;
   wire n_0_1_108;
   wire n_0_1_109;
   wire n_0_261;
   wire n_0_263;
   wire n_0_264;
   wire n_0_1_110;
   wire n_0_1_111;
   wire n_0_262;
   wire n_0_1_112;
   wire n_0_1_113;
   wire n_0_1_114;
   wire n_0_265;
   wire n_0_266;
   wire n_0_1_115;
   wire n_0_1_116;
   wire n_0_1_117;
   wire n_0_1_118;
   wire n_0_1_119;
   wire n_0_1_120;
   wire n_0_1_121;
   wire n_0_1_122;
   wire n_0_1_123;
   wire n_0_1_124;
   wire n_0_1_125;
   wire n_0_1_126;
   wire n_0_1_127;
   wire n_0_1_128;
   wire n_0_1_129;
   wire n_0_1_130;
   wire n_0_1_131;
   wire n_0_1_132;
   wire n_0_1_133;
   wire n_0_1_134;
   wire n_0_1_135;
   wire n_0_1_136;
   wire n_0_1_137;
   wire n_0_1_138;
   wire n_0_1_139;
   wire n_0_1_140;
   wire n_0_1_141;
   wire n_0_1_142;

   datapath i_0_0 (.B(B), .p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, uc_0}));
   datapath__0_0 i_0_2 (.A(A), .p_0({n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, 
      n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, 
      n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, 
      n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, uc_1}));
   datapath__0_18 i_0_4 (.p_0({accumulator[31], accumulator[30], accumulator[29], 
      accumulator[28], accumulator[27], accumulator[26], accumulator[25], 
      accumulator[24], accumulator[23], accumulator[22], accumulator[21], 
      accumulator[20], accumulator[19], accumulator[18], accumulator[17], 
      accumulator[16], accumulator[15], accumulator[14], accumulator[13], 
      accumulator[12], accumulator[11], accumulator[10], accumulator[9], 
      accumulator[8], accumulator[7], accumulator[6], accumulator[5], 
      accumulator[4], accumulator[3], accumulator[2], accumulator[1], 
      accumulator[0], multiplicand[31], multiplicand[30], multiplicand[29], 
      multiplicand[28], multiplicand[27], multiplicand[26], multiplicand[25], 
      multiplicand[24], multiplicand[23], multiplicand[22], multiplicand[21], 
      multiplicand[20], multiplicand[19], multiplicand[18], multiplicand[17], 
      multiplicand[16], multiplicand[15], multiplicand[14], multiplicand[13], 
      multiplicand[12], multiplicand[11], multiplicand[10], multiplicand[9], 
      multiplicand[8], multiplicand[7], multiplicand[6], multiplicand[5], 
      multiplicand[4], multiplicand[3], multiplicand[2], multiplicand[1], Res[0]}), 
      .p_1({n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, 
      n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, 
      n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, 
      n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, 
      n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, 
      n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, 
      n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, 
      n_0_65, n_0_64, n_0_63, n_0_62, uc_2}));
   DLH_X1 \isNeg_reg[1]  (.D(n_0_266), .G(n_0_262), .Q(isNeg[1]));
   DLH_X1 \isNeg_reg[0]  (.D(n_0_265), .G(n_0_262), .Q(isNeg[0]));
   datapath__0_5 i_0_13 (.multiplier(multiplier), .accumulator(accumulator), 
      .p_0({n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, n_0_151, 
      n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, n_0_143, 
      n_0_142, n_0_141, n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, 
      n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, 
      n_0_126, n_0_125}));
   DLH_X1 \accumulator_reg[31]  (.D(n_0_197), .G(n_0_165), .Q(accumulator[31]));
   DLH_X1 \accumulator_reg[30]  (.D(n_0_196), .G(n_0_165), .Q(accumulator[30]));
   DLH_X1 \accumulator_reg[29]  (.D(n_0_195), .G(n_0_165), .Q(accumulator[29]));
   DLH_X1 \accumulator_reg[28]  (.D(n_0_194), .G(n_0_165), .Q(accumulator[28]));
   DLH_X1 \accumulator_reg[27]  (.D(n_0_193), .G(n_0_165), .Q(accumulator[27]));
   DLH_X1 \accumulator_reg[26]  (.D(n_0_192), .G(n_0_165), .Q(accumulator[26]));
   DLH_X1 \accumulator_reg[25]  (.D(n_0_191), .G(n_0_165), .Q(accumulator[25]));
   DLH_X1 \accumulator_reg[24]  (.D(n_0_190), .G(n_0_165), .Q(accumulator[24]));
   DLH_X1 \accumulator_reg[23]  (.D(n_0_189), .G(n_0_165), .Q(accumulator[23]));
   DLH_X1 \accumulator_reg[22]  (.D(n_0_188), .G(n_0_165), .Q(accumulator[22]));
   DLH_X1 \accumulator_reg[21]  (.D(n_0_187), .G(n_0_165), .Q(accumulator[21]));
   DLH_X1 \accumulator_reg[20]  (.D(n_0_186), .G(n_0_165), .Q(accumulator[20]));
   DLH_X1 \accumulator_reg[19]  (.D(n_0_185), .G(n_0_165), .Q(accumulator[19]));
   DLH_X1 \accumulator_reg[18]  (.D(n_0_184), .G(n_0_165), .Q(accumulator[18]));
   DLH_X1 \accumulator_reg[17]  (.D(n_0_183), .G(n_0_165), .Q(accumulator[17]));
   DLH_X1 \accumulator_reg[16]  (.D(n_0_182), .G(n_0_165), .Q(accumulator[16]));
   DLH_X1 \accumulator_reg[15]  (.D(n_0_181), .G(n_0_165), .Q(accumulator[15]));
   DLH_X1 \accumulator_reg[14]  (.D(n_0_180), .G(n_0_165), .Q(accumulator[14]));
   DLH_X1 \accumulator_reg[13]  (.D(n_0_179), .G(n_0_165), .Q(accumulator[13]));
   DLH_X1 \accumulator_reg[12]  (.D(n_0_178), .G(n_0_165), .Q(accumulator[12]));
   DLH_X1 \accumulator_reg[11]  (.D(n_0_177), .G(n_0_165), .Q(accumulator[11]));
   DLH_X1 \accumulator_reg[10]  (.D(n_0_176), .G(n_0_165), .Q(accumulator[10]));
   DLH_X1 \accumulator_reg[9]  (.D(n_0_175), .G(n_0_165), .Q(accumulator[9]));
   DLH_X1 \accumulator_reg[8]  (.D(n_0_174), .G(n_0_165), .Q(accumulator[8]));
   DLH_X1 \accumulator_reg[7]  (.D(n_0_173), .G(n_0_165), .Q(accumulator[7]));
   DLH_X1 \accumulator_reg[6]  (.D(n_0_172), .G(n_0_165), .Q(accumulator[6]));
   DLH_X1 \accumulator_reg[5]  (.D(n_0_171), .G(n_0_165), .Q(accumulator[5]));
   DLH_X1 \accumulator_reg[4]  (.D(n_0_170), .G(n_0_165), .Q(accumulator[4]));
   DLH_X1 \accumulator_reg[3]  (.D(n_0_169), .G(n_0_165), .Q(accumulator[3]));
   DLH_X1 \accumulator_reg[2]  (.D(n_0_168), .G(n_0_165), .Q(accumulator[2]));
   DLH_X1 \accumulator_reg[1]  (.D(n_0_167), .G(n_0_165), .Q(accumulator[1]));
   DLH_X1 \accumulator_reg[0]  (.D(n_0_166), .G(n_0_165), .Q(accumulator[0]));
   DLH_X1 \multiplicand_reg[31]  (.D(n_0_229), .G(n_0_165), .Q(multiplicand[31]));
   DLH_X1 \multiplicand_reg[30]  (.D(n_0_228), .G(n_0_165), .Q(multiplicand[30]));
   DLH_X1 \multiplicand_reg[29]  (.D(n_0_227), .G(n_0_165), .Q(multiplicand[29]));
   DLH_X1 \multiplicand_reg[28]  (.D(n_0_226), .G(n_0_165), .Q(multiplicand[28]));
   DLH_X1 \multiplicand_reg[27]  (.D(n_0_225), .G(n_0_165), .Q(multiplicand[27]));
   DLH_X1 \multiplicand_reg[26]  (.D(n_0_224), .G(n_0_165), .Q(multiplicand[26]));
   DLH_X1 \multiplicand_reg[25]  (.D(n_0_223), .G(n_0_165), .Q(multiplicand[25]));
   DLH_X1 \multiplicand_reg[24]  (.D(n_0_222), .G(n_0_165), .Q(multiplicand[24]));
   DLH_X1 \multiplicand_reg[23]  (.D(n_0_221), .G(n_0_165), .Q(multiplicand[23]));
   DLH_X1 \multiplicand_reg[22]  (.D(n_0_220), .G(n_0_165), .Q(multiplicand[22]));
   DLH_X1 \multiplicand_reg[21]  (.D(n_0_219), .G(n_0_165), .Q(multiplicand[21]));
   DLH_X1 \multiplicand_reg[20]  (.D(n_0_218), .G(n_0_165), .Q(multiplicand[20]));
   DLH_X1 \multiplicand_reg[19]  (.D(n_0_217), .G(n_0_165), .Q(multiplicand[19]));
   DLH_X1 \multiplicand_reg[18]  (.D(n_0_216), .G(n_0_165), .Q(multiplicand[18]));
   DLH_X1 \multiplicand_reg[17]  (.D(n_0_215), .G(n_0_165), .Q(multiplicand[17]));
   DLH_X1 \multiplicand_reg[16]  (.D(n_0_214), .G(n_0_165), .Q(multiplicand[16]));
   DLH_X1 \multiplicand_reg[15]  (.D(n_0_213), .G(n_0_165), .Q(multiplicand[15]));
   DLH_X1 \multiplicand_reg[14]  (.D(n_0_212), .G(n_0_165), .Q(multiplicand[14]));
   DLH_X1 \multiplicand_reg[13]  (.D(n_0_211), .G(n_0_165), .Q(multiplicand[13]));
   DLH_X1 \multiplicand_reg[12]  (.D(n_0_210), .G(n_0_165), .Q(multiplicand[12]));
   DLH_X1 \multiplicand_reg[11]  (.D(n_0_209), .G(n_0_165), .Q(multiplicand[11]));
   DLH_X1 \multiplicand_reg[10]  (.D(n_0_208), .G(n_0_165), .Q(multiplicand[10]));
   DLH_X1 \multiplicand_reg[9]  (.D(n_0_207), .G(n_0_165), .Q(multiplicand[9]));
   DLH_X1 \multiplicand_reg[8]  (.D(n_0_206), .G(n_0_165), .Q(multiplicand[8]));
   DLH_X1 \multiplicand_reg[7]  (.D(n_0_205), .G(n_0_165), .Q(multiplicand[7]));
   DLH_X1 \multiplicand_reg[6]  (.D(n_0_204), .G(n_0_165), .Q(multiplicand[6]));
   DLH_X1 \multiplicand_reg[5]  (.D(n_0_203), .G(n_0_165), .Q(multiplicand[5]));
   DLH_X1 \multiplicand_reg[4]  (.D(n_0_202), .G(n_0_165), .Q(multiplicand[4]));
   DLH_X1 \multiplicand_reg[3]  (.D(n_0_201), .G(n_0_165), .Q(multiplicand[3]));
   DLH_X1 \multiplicand_reg[2]  (.D(n_0_200), .G(n_0_165), .Q(multiplicand[2]));
   DLH_X1 \multiplicand_reg[1]  (.D(n_0_199), .G(n_0_165), .Q(multiplicand[1]));
   DLH_X1 \multiplicand_reg[0]  (.D(n_0_198), .G(n_0_165), .Q(Res[0]));
   DLH_X1 ready_reg (.D(n_0_158), .G(n_0_159), .Q(ready));
   DLH_X1 \multiplier_reg[31]  (.D(n_0_261), .G(n_0_262), .Q(multiplier[31]));
   DLH_X1 \multiplier_reg[30]  (.D(n_0_260), .G(n_0_262), .Q(multiplier[30]));
   DLH_X1 \multiplier_reg[29]  (.D(n_0_259), .G(n_0_262), .Q(multiplier[29]));
   DLH_X1 \multiplier_reg[28]  (.D(n_0_258), .G(n_0_262), .Q(multiplier[28]));
   DLH_X1 \multiplier_reg[27]  (.D(n_0_257), .G(n_0_262), .Q(multiplier[27]));
   DLH_X1 \multiplier_reg[26]  (.D(n_0_256), .G(n_0_262), .Q(multiplier[26]));
   DLH_X1 \multiplier_reg[25]  (.D(n_0_255), .G(n_0_262), .Q(multiplier[25]));
   DLH_X1 \multiplier_reg[24]  (.D(n_0_254), .G(n_0_262), .Q(multiplier[24]));
   DLH_X1 \multiplier_reg[23]  (.D(n_0_253), .G(n_0_262), .Q(multiplier[23]));
   DLH_X1 \multiplier_reg[22]  (.D(n_0_252), .G(n_0_262), .Q(multiplier[22]));
   DLH_X1 \multiplier_reg[21]  (.D(n_0_251), .G(n_0_262), .Q(multiplier[21]));
   DLH_X1 \multiplier_reg[20]  (.D(n_0_250), .G(n_0_262), .Q(multiplier[20]));
   DLH_X1 \multiplier_reg[19]  (.D(n_0_249), .G(n_0_262), .Q(multiplier[19]));
   DLH_X1 \multiplier_reg[18]  (.D(n_0_248), .G(n_0_262), .Q(multiplier[18]));
   DLH_X1 \multiplier_reg[17]  (.D(n_0_247), .G(n_0_262), .Q(multiplier[17]));
   DLH_X1 \multiplier_reg[16]  (.D(n_0_246), .G(n_0_262), .Q(multiplier[16]));
   DLH_X1 \multiplier_reg[15]  (.D(n_0_245), .G(n_0_262), .Q(multiplier[15]));
   DLH_X1 \multiplier_reg[14]  (.D(n_0_244), .G(n_0_262), .Q(multiplier[14]));
   DLH_X1 \multiplier_reg[13]  (.D(n_0_243), .G(n_0_262), .Q(multiplier[13]));
   DLH_X1 \multiplier_reg[12]  (.D(n_0_242), .G(n_0_262), .Q(multiplier[12]));
   DLH_X1 \multiplier_reg[11]  (.D(n_0_241), .G(n_0_262), .Q(multiplier[11]));
   DLH_X1 \multiplier_reg[10]  (.D(n_0_240), .G(n_0_262), .Q(multiplier[10]));
   DLH_X1 \multiplier_reg[9]  (.D(n_0_239), .G(n_0_262), .Q(multiplier[9]));
   DLH_X1 \multiplier_reg[8]  (.D(n_0_238), .G(n_0_262), .Q(multiplier[8]));
   DLH_X1 \multiplier_reg[7]  (.D(n_0_237), .G(n_0_262), .Q(multiplier[7]));
   DLH_X1 \multiplier_reg[6]  (.D(n_0_236), .G(n_0_262), .Q(multiplier[6]));
   DLH_X1 \multiplier_reg[5]  (.D(n_0_235), .G(n_0_262), .Q(multiplier[5]));
   DLH_X1 \multiplier_reg[4]  (.D(n_0_234), .G(n_0_262), .Q(multiplier[4]));
   DLH_X1 \multiplier_reg[3]  (.D(n_0_233), .G(n_0_262), .Q(multiplier[3]));
   DLH_X1 \multiplier_reg[2]  (.D(n_0_232), .G(n_0_262), .Q(multiplier[2]));
   DLH_X1 \multiplier_reg[1]  (.D(n_0_231), .G(n_0_262), .Q(multiplier[1]));
   DLH_X1 \multiplier_reg[0]  (.D(n_0_230), .G(n_0_262), .Q(multiplier[0]));
   DLH_X1 carry_reg (.D(n_0_263), .G(n_0_264), .Q(carry));
   DLH_X1 \counter_reg[4]  (.D(n_0_164), .G(n_0_165), .Q(counter[4]));
   DLH_X1 \counter_reg[3]  (.D(n_0_163), .G(n_0_165), .Q(counter[3]));
   DLH_X1 \counter_reg[2]  (.D(n_0_162), .G(n_0_165), .Q(counter[2]));
   DLH_X1 \counter_reg[1]  (.D(n_0_161), .G(n_0_165), .Q(counter[1]));
   DLH_X1 \counter_reg[0]  (.D(n_0_160), .G(n_0_165), .Q(counter[0]));
   OAI211_X1 i_0_1_0 (.A(n_0_1_139), .B(clk), .C1(ready), .C2(enable), .ZN(
      n_0_158));
   OAI21_X1 i_0_1_1 (.A(n_0_1_112), .B1(n_0_1_7), .B2(n_0_1_0), .ZN(n_0_159));
   NAND3_X1 i_0_1_2 (.A1(n_0_1_111), .A2(n_0_1_142), .A3(counter[0]), .ZN(
      n_0_1_0));
   NOR2_X1 i_0_1_3 (.A1(n_0_262), .A2(counter[0]), .ZN(n_0_160));
   NOR2_X1 i_0_1_4 (.A1(n_0_1_1), .A2(n_0_262), .ZN(n_0_161));
   XOR2_X1 i_0_1_5 (.A(counter[1]), .B(counter[0]), .Z(n_0_1_1));
   AOI21_X1 i_0_1_6 (.A(n_0_262), .B1(n_0_1_6), .B2(n_0_1_2), .ZN(n_0_162));
   OAI21_X1 i_0_1_7 (.A(counter[2]), .B1(counter[1]), .B2(counter[0]), .ZN(
      n_0_1_2));
   NOR2_X1 i_0_1_8 (.A1(n_0_1_3), .A2(n_0_262), .ZN(n_0_163));
   XOR2_X1 i_0_1_9 (.A(counter[3]), .B(n_0_1_6), .Z(n_0_1_3));
   AOI21_X1 i_0_1_10 (.A(n_0_262), .B1(n_0_1_5), .B2(n_0_1_4), .ZN(n_0_164));
   OR3_X1 i_0_1_11 (.A1(n_0_1_7), .A2(counter[0]), .A3(counter[4]), .ZN(n_0_1_4));
   OAI21_X1 i_0_1_12 (.A(counter[4]), .B1(n_0_1_7), .B2(counter[0]), .ZN(n_0_1_5));
   OR3_X1 i_0_1_13 (.A1(counter[2]), .A2(counter[1]), .A3(counter[0]), .ZN(
      n_0_1_6));
   OR3_X1 i_0_1_14 (.A1(counter[3]), .A2(counter[2]), .A3(counter[1]), .ZN(
      n_0_1_7));
   NAND2_X1 i_0_1_15 (.A1(n_0_1_139), .A2(n_0_1_8), .ZN(n_0_165));
   XNOR2_X1 i_0_1_16 (.A(ready), .B(n_0_1_114), .ZN(n_0_1_8));
   INV_X1 i_0_1_17 (.A(n_0_1_9), .ZN(n_0_166));
   AOI22_X1 i_0_1_18 (.A1(n_0_126), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[1]), .ZN(n_0_1_9));
   INV_X1 i_0_1_19 (.A(n_0_1_10), .ZN(n_0_167));
   AOI22_X1 i_0_1_20 (.A1(n_0_127), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[2]), .ZN(n_0_1_10));
   INV_X1 i_0_1_21 (.A(n_0_1_11), .ZN(n_0_168));
   AOI22_X1 i_0_1_22 (.A1(n_0_128), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[3]), .ZN(n_0_1_11));
   INV_X1 i_0_1_23 (.A(n_0_1_12), .ZN(n_0_169));
   AOI22_X1 i_0_1_24 (.A1(n_0_129), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[4]), .ZN(n_0_1_12));
   INV_X1 i_0_1_25 (.A(n_0_1_13), .ZN(n_0_170));
   AOI22_X1 i_0_1_26 (.A1(n_0_130), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[5]), .ZN(n_0_1_13));
   INV_X1 i_0_1_27 (.A(n_0_1_14), .ZN(n_0_171));
   AOI22_X1 i_0_1_28 (.A1(n_0_131), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[6]), .ZN(n_0_1_14));
   INV_X1 i_0_1_29 (.A(n_0_1_15), .ZN(n_0_172));
   AOI22_X1 i_0_1_30 (.A1(n_0_132), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[7]), .ZN(n_0_1_15));
   INV_X1 i_0_1_31 (.A(n_0_1_16), .ZN(n_0_173));
   AOI22_X1 i_0_1_32 (.A1(n_0_133), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[8]), .ZN(n_0_1_16));
   INV_X1 i_0_1_33 (.A(n_0_1_17), .ZN(n_0_174));
   AOI22_X1 i_0_1_34 (.A1(n_0_134), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[9]), .ZN(n_0_1_17));
   INV_X1 i_0_1_35 (.A(n_0_1_18), .ZN(n_0_175));
   AOI22_X1 i_0_1_36 (.A1(n_0_135), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[10]), .ZN(n_0_1_18));
   INV_X1 i_0_1_37 (.A(n_0_1_19), .ZN(n_0_176));
   AOI22_X1 i_0_1_38 (.A1(n_0_136), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[11]), .ZN(n_0_1_19));
   INV_X1 i_0_1_39 (.A(n_0_1_20), .ZN(n_0_177));
   AOI22_X1 i_0_1_40 (.A1(n_0_137), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[12]), .ZN(n_0_1_20));
   INV_X1 i_0_1_41 (.A(n_0_1_21), .ZN(n_0_178));
   AOI22_X1 i_0_1_42 (.A1(n_0_138), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[13]), .ZN(n_0_1_21));
   INV_X1 i_0_1_43 (.A(n_0_1_22), .ZN(n_0_179));
   AOI22_X1 i_0_1_44 (.A1(n_0_139), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[14]), .ZN(n_0_1_22));
   INV_X1 i_0_1_45 (.A(n_0_1_23), .ZN(n_0_180));
   AOI22_X1 i_0_1_46 (.A1(n_0_140), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[15]), .ZN(n_0_1_23));
   INV_X1 i_0_1_47 (.A(n_0_1_24), .ZN(n_0_181));
   AOI22_X1 i_0_1_48 (.A1(n_0_141), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[16]), .ZN(n_0_1_24));
   INV_X1 i_0_1_49 (.A(n_0_1_25), .ZN(n_0_182));
   AOI22_X1 i_0_1_50 (.A1(n_0_142), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[17]), .ZN(n_0_1_25));
   INV_X1 i_0_1_51 (.A(n_0_1_26), .ZN(n_0_183));
   AOI22_X1 i_0_1_52 (.A1(n_0_143), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[18]), .ZN(n_0_1_26));
   INV_X1 i_0_1_53 (.A(n_0_1_27), .ZN(n_0_184));
   AOI22_X1 i_0_1_54 (.A1(n_0_144), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[19]), .ZN(n_0_1_27));
   INV_X1 i_0_1_55 (.A(n_0_1_28), .ZN(n_0_185));
   AOI22_X1 i_0_1_56 (.A1(n_0_145), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[20]), .ZN(n_0_1_28));
   INV_X1 i_0_1_57 (.A(n_0_1_29), .ZN(n_0_186));
   AOI22_X1 i_0_1_58 (.A1(n_0_146), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[21]), .ZN(n_0_1_29));
   INV_X1 i_0_1_59 (.A(n_0_1_30), .ZN(n_0_187));
   AOI22_X1 i_0_1_60 (.A1(n_0_147), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[22]), .ZN(n_0_1_30));
   INV_X1 i_0_1_61 (.A(n_0_1_31), .ZN(n_0_188));
   AOI22_X1 i_0_1_62 (.A1(n_0_148), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[23]), .ZN(n_0_1_31));
   INV_X1 i_0_1_63 (.A(n_0_1_32), .ZN(n_0_189));
   AOI22_X1 i_0_1_64 (.A1(n_0_149), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[24]), .ZN(n_0_1_32));
   INV_X1 i_0_1_65 (.A(n_0_1_33), .ZN(n_0_190));
   AOI22_X1 i_0_1_66 (.A1(n_0_150), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[25]), .ZN(n_0_1_33));
   INV_X1 i_0_1_67 (.A(n_0_1_34), .ZN(n_0_191));
   AOI22_X1 i_0_1_68 (.A1(n_0_151), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[26]), .ZN(n_0_1_34));
   INV_X1 i_0_1_69 (.A(n_0_1_35), .ZN(n_0_192));
   AOI22_X1 i_0_1_70 (.A1(n_0_152), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[27]), .ZN(n_0_1_35));
   INV_X1 i_0_1_71 (.A(n_0_1_36), .ZN(n_0_193));
   AOI22_X1 i_0_1_72 (.A1(n_0_153), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[28]), .ZN(n_0_1_36));
   INV_X1 i_0_1_73 (.A(n_0_1_37), .ZN(n_0_194));
   AOI22_X1 i_0_1_74 (.A1(n_0_154), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[29]), .ZN(n_0_1_37));
   INV_X1 i_0_1_75 (.A(n_0_1_38), .ZN(n_0_195));
   AOI22_X1 i_0_1_76 (.A1(n_0_155), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[30]), .ZN(n_0_1_38));
   INV_X1 i_0_1_77 (.A(n_0_1_39), .ZN(n_0_196));
   AOI22_X1 i_0_1_78 (.A1(n_0_156), .A2(n_0_1_42), .B1(n_0_1_41), .B2(
      accumulator[31]), .ZN(n_0_1_39));
   INV_X1 i_0_1_79 (.A(n_0_1_40), .ZN(n_0_197));
   AOI22_X1 i_0_1_80 (.A1(n_0_157), .A2(n_0_1_42), .B1(n_0_1_41), .B2(carry), 
      .ZN(n_0_1_40));
   NOR2_X1 i_0_1_81 (.A1(n_0_262), .A2(Res[0]), .ZN(n_0_1_41));
   AND2_X1 i_0_1_82 (.A1(Res[0]), .A2(n_0_1_112), .ZN(n_0_1_42));
   INV_X1 i_0_1_83 (.A(n_0_1_43), .ZN(n_0_198));
   AOI22_X1 i_0_1_84 (.A1(multiplicand[1]), .A2(n_0_1_112), .B1(n_0_1_78), 
      .B2(B[0]), .ZN(n_0_1_43));
   INV_X1 i_0_1_85 (.A(n_0_1_44), .ZN(n_0_199));
   AOI222_X1 i_0_1_86 (.A1(multiplicand[2]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_0), .C1(B[1]), .C2(n_0_1_74), .ZN(n_0_1_44));
   INV_X1 i_0_1_87 (.A(n_0_1_45), .ZN(n_0_200));
   AOI222_X1 i_0_1_88 (.A1(multiplicand[3]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_1), .C1(B[2]), .C2(n_0_1_74), .ZN(n_0_1_45));
   INV_X1 i_0_1_89 (.A(n_0_1_46), .ZN(n_0_201));
   AOI222_X1 i_0_1_90 (.A1(multiplicand[4]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_2), .C1(B[3]), .C2(n_0_1_74), .ZN(n_0_1_46));
   INV_X1 i_0_1_91 (.A(n_0_1_47), .ZN(n_0_202));
   AOI222_X1 i_0_1_92 (.A1(multiplicand[5]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_3), .C1(B[4]), .C2(n_0_1_74), .ZN(n_0_1_47));
   INV_X1 i_0_1_93 (.A(n_0_1_48), .ZN(n_0_203));
   AOI222_X1 i_0_1_94 (.A1(multiplicand[6]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_4), .C1(B[5]), .C2(n_0_1_74), .ZN(n_0_1_48));
   INV_X1 i_0_1_95 (.A(n_0_1_49), .ZN(n_0_204));
   AOI222_X1 i_0_1_96 (.A1(multiplicand[7]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_5), .C1(B[6]), .C2(n_0_1_74), .ZN(n_0_1_49));
   INV_X1 i_0_1_97 (.A(n_0_1_50), .ZN(n_0_205));
   AOI222_X1 i_0_1_98 (.A1(multiplicand[8]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_6), .C1(B[7]), .C2(n_0_1_74), .ZN(n_0_1_50));
   INV_X1 i_0_1_99 (.A(n_0_1_51), .ZN(n_0_206));
   AOI222_X1 i_0_1_100 (.A1(multiplicand[9]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_7), .C1(B[8]), .C2(n_0_1_74), .ZN(n_0_1_51));
   INV_X1 i_0_1_101 (.A(n_0_1_52), .ZN(n_0_207));
   AOI222_X1 i_0_1_102 (.A1(multiplicand[10]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_8), .C1(B[9]), .C2(n_0_1_74), .ZN(n_0_1_52));
   INV_X1 i_0_1_103 (.A(n_0_1_53), .ZN(n_0_208));
   AOI222_X1 i_0_1_104 (.A1(multiplicand[11]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_9), .C1(B[10]), .C2(n_0_1_74), .ZN(n_0_1_53));
   INV_X1 i_0_1_105 (.A(n_0_1_54), .ZN(n_0_209));
   AOI222_X1 i_0_1_106 (.A1(multiplicand[12]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_10), .C1(B[11]), .C2(n_0_1_74), .ZN(n_0_1_54));
   INV_X1 i_0_1_107 (.A(n_0_1_55), .ZN(n_0_210));
   AOI222_X1 i_0_1_108 (.A1(multiplicand[13]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_11), .C1(B[12]), .C2(n_0_1_74), .ZN(n_0_1_55));
   INV_X1 i_0_1_109 (.A(n_0_1_56), .ZN(n_0_211));
   AOI222_X1 i_0_1_110 (.A1(multiplicand[14]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_12), .C1(B[13]), .C2(n_0_1_74), .ZN(n_0_1_56));
   INV_X1 i_0_1_111 (.A(n_0_1_57), .ZN(n_0_212));
   AOI222_X1 i_0_1_112 (.A1(multiplicand[15]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_13), .C1(B[14]), .C2(n_0_1_74), .ZN(n_0_1_57));
   INV_X1 i_0_1_113 (.A(n_0_1_58), .ZN(n_0_213));
   AOI222_X1 i_0_1_114 (.A1(multiplicand[16]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_14), .C1(B[15]), .C2(n_0_1_74), .ZN(n_0_1_58));
   INV_X1 i_0_1_115 (.A(n_0_1_59), .ZN(n_0_214));
   AOI222_X1 i_0_1_116 (.A1(multiplicand[17]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_15), .C1(B[16]), .C2(n_0_1_74), .ZN(n_0_1_59));
   INV_X1 i_0_1_117 (.A(n_0_1_60), .ZN(n_0_215));
   AOI222_X1 i_0_1_118 (.A1(multiplicand[18]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_16), .C1(B[17]), .C2(n_0_1_74), .ZN(n_0_1_60));
   INV_X1 i_0_1_119 (.A(n_0_1_61), .ZN(n_0_216));
   AOI222_X1 i_0_1_120 (.A1(multiplicand[19]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_17), .C1(B[18]), .C2(n_0_1_74), .ZN(n_0_1_61));
   INV_X1 i_0_1_121 (.A(n_0_1_62), .ZN(n_0_217));
   AOI222_X1 i_0_1_122 (.A1(multiplicand[20]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_18), .C1(B[19]), .C2(n_0_1_74), .ZN(n_0_1_62));
   INV_X1 i_0_1_123 (.A(n_0_1_63), .ZN(n_0_218));
   AOI222_X1 i_0_1_124 (.A1(multiplicand[21]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_19), .C1(B[20]), .C2(n_0_1_74), .ZN(n_0_1_63));
   INV_X1 i_0_1_125 (.A(n_0_1_64), .ZN(n_0_219));
   AOI222_X1 i_0_1_126 (.A1(multiplicand[22]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_20), .C1(B[21]), .C2(n_0_1_74), .ZN(n_0_1_64));
   INV_X1 i_0_1_127 (.A(n_0_1_65), .ZN(n_0_220));
   AOI222_X1 i_0_1_128 (.A1(multiplicand[23]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_21), .C1(B[22]), .C2(n_0_1_74), .ZN(n_0_1_65));
   INV_X1 i_0_1_129 (.A(n_0_1_66), .ZN(n_0_221));
   AOI222_X1 i_0_1_130 (.A1(multiplicand[24]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_22), .C1(B[23]), .C2(n_0_1_74), .ZN(n_0_1_66));
   INV_X1 i_0_1_131 (.A(n_0_1_67), .ZN(n_0_222));
   AOI222_X1 i_0_1_132 (.A1(multiplicand[25]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_23), .C1(B[24]), .C2(n_0_1_74), .ZN(n_0_1_67));
   INV_X1 i_0_1_133 (.A(n_0_1_68), .ZN(n_0_223));
   AOI222_X1 i_0_1_134 (.A1(multiplicand[26]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_24), .C1(B[25]), .C2(n_0_1_74), .ZN(n_0_1_68));
   INV_X1 i_0_1_135 (.A(n_0_1_69), .ZN(n_0_224));
   AOI222_X1 i_0_1_136 (.A1(multiplicand[27]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_25), .C1(B[26]), .C2(n_0_1_74), .ZN(n_0_1_69));
   INV_X1 i_0_1_137 (.A(n_0_1_70), .ZN(n_0_225));
   AOI222_X1 i_0_1_138 (.A1(multiplicand[28]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_26), .C1(B[27]), .C2(n_0_1_74), .ZN(n_0_1_70));
   INV_X1 i_0_1_139 (.A(n_0_1_71), .ZN(n_0_226));
   AOI222_X1 i_0_1_140 (.A1(multiplicand[29]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_27), .C1(B[28]), .C2(n_0_1_74), .ZN(n_0_1_71));
   INV_X1 i_0_1_141 (.A(n_0_1_72), .ZN(n_0_227));
   AOI222_X1 i_0_1_142 (.A1(multiplicand[30]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_28), .C1(B[29]), .C2(n_0_1_74), .ZN(n_0_1_72));
   INV_X1 i_0_1_143 (.A(n_0_1_73), .ZN(n_0_228));
   AOI222_X1 i_0_1_144 (.A1(multiplicand[31]), .A2(n_0_1_112), .B1(n_0_1_77), 
      .B2(n_0_29), .C1(B[30]), .C2(n_0_1_74), .ZN(n_0_1_73));
   NOR3_X1 i_0_1_145 (.A1(n_0_1_113), .A2(reset), .A3(B[31]), .ZN(n_0_1_74));
   INV_X1 i_0_1_146 (.A(n_0_1_75), .ZN(n_0_229));
   AOI22_X1 i_0_1_147 (.A1(n_0_1_76), .A2(n_0_1_112), .B1(n_0_30), .B2(n_0_1_77), 
      .ZN(n_0_1_75));
   MUX2_X1 i_0_1_148 (.A(accumulator[0]), .B(n_0_125), .S(Res[0]), .Z(n_0_1_76));
   NOR3_X1 i_0_1_149 (.A1(n_0_1_141), .A2(n_0_1_113), .A3(reset), .ZN(n_0_1_77));
   NOR2_X1 i_0_1_150 (.A1(n_0_1_113), .A2(reset), .ZN(n_0_1_78));
   AND2_X1 i_0_1_151 (.A1(n_0_1_139), .A2(A[0]), .ZN(n_0_230));
   INV_X1 i_0_1_152 (.A(n_0_1_79), .ZN(n_0_231));
   AOI22_X1 i_0_1_153 (.A1(n_0_31), .A2(n_0_266), .B1(n_0_1_109), .B2(A[1]), 
      .ZN(n_0_1_79));
   INV_X1 i_0_1_154 (.A(n_0_1_80), .ZN(n_0_232));
   AOI22_X1 i_0_1_155 (.A1(n_0_32), .A2(n_0_266), .B1(n_0_1_109), .B2(A[2]), 
      .ZN(n_0_1_80));
   INV_X1 i_0_1_156 (.A(n_0_1_81), .ZN(n_0_233));
   AOI22_X1 i_0_1_157 (.A1(n_0_33), .A2(n_0_266), .B1(n_0_1_109), .B2(A[3]), 
      .ZN(n_0_1_81));
   INV_X1 i_0_1_158 (.A(n_0_1_82), .ZN(n_0_234));
   AOI22_X1 i_0_1_159 (.A1(n_0_34), .A2(n_0_266), .B1(n_0_1_109), .B2(A[4]), 
      .ZN(n_0_1_82));
   INV_X1 i_0_1_160 (.A(n_0_1_83), .ZN(n_0_235));
   AOI22_X1 i_0_1_161 (.A1(n_0_35), .A2(n_0_266), .B1(n_0_1_109), .B2(A[5]), 
      .ZN(n_0_1_83));
   INV_X1 i_0_1_162 (.A(n_0_1_84), .ZN(n_0_236));
   AOI22_X1 i_0_1_163 (.A1(n_0_36), .A2(n_0_266), .B1(n_0_1_109), .B2(A[6]), 
      .ZN(n_0_1_84));
   INV_X1 i_0_1_164 (.A(n_0_1_85), .ZN(n_0_237));
   AOI22_X1 i_0_1_165 (.A1(n_0_37), .A2(n_0_266), .B1(n_0_1_109), .B2(A[7]), 
      .ZN(n_0_1_85));
   INV_X1 i_0_1_166 (.A(n_0_1_86), .ZN(n_0_238));
   AOI22_X1 i_0_1_167 (.A1(n_0_38), .A2(n_0_266), .B1(n_0_1_109), .B2(A[8]), 
      .ZN(n_0_1_86));
   INV_X1 i_0_1_168 (.A(n_0_1_87), .ZN(n_0_239));
   AOI22_X1 i_0_1_169 (.A1(n_0_39), .A2(n_0_266), .B1(n_0_1_109), .B2(A[9]), 
      .ZN(n_0_1_87));
   INV_X1 i_0_1_170 (.A(n_0_1_88), .ZN(n_0_240));
   AOI22_X1 i_0_1_171 (.A1(n_0_40), .A2(n_0_266), .B1(n_0_1_109), .B2(A[10]), 
      .ZN(n_0_1_88));
   INV_X1 i_0_1_172 (.A(n_0_1_89), .ZN(n_0_241));
   AOI22_X1 i_0_1_173 (.A1(n_0_41), .A2(n_0_266), .B1(n_0_1_109), .B2(A[11]), 
      .ZN(n_0_1_89));
   INV_X1 i_0_1_174 (.A(n_0_1_90), .ZN(n_0_242));
   AOI22_X1 i_0_1_175 (.A1(n_0_42), .A2(n_0_266), .B1(n_0_1_109), .B2(A[12]), 
      .ZN(n_0_1_90));
   INV_X1 i_0_1_176 (.A(n_0_1_91), .ZN(n_0_243));
   AOI22_X1 i_0_1_177 (.A1(n_0_43), .A2(n_0_266), .B1(n_0_1_109), .B2(A[13]), 
      .ZN(n_0_1_91));
   INV_X1 i_0_1_178 (.A(n_0_1_92), .ZN(n_0_244));
   AOI22_X1 i_0_1_179 (.A1(n_0_44), .A2(n_0_266), .B1(n_0_1_109), .B2(A[14]), 
      .ZN(n_0_1_92));
   INV_X1 i_0_1_180 (.A(n_0_1_93), .ZN(n_0_245));
   AOI22_X1 i_0_1_181 (.A1(n_0_45), .A2(n_0_266), .B1(n_0_1_109), .B2(A[15]), 
      .ZN(n_0_1_93));
   INV_X1 i_0_1_182 (.A(n_0_1_94), .ZN(n_0_246));
   AOI22_X1 i_0_1_183 (.A1(n_0_46), .A2(n_0_266), .B1(n_0_1_109), .B2(A[16]), 
      .ZN(n_0_1_94));
   INV_X1 i_0_1_184 (.A(n_0_1_95), .ZN(n_0_247));
   AOI22_X1 i_0_1_185 (.A1(n_0_47), .A2(n_0_266), .B1(n_0_1_109), .B2(A[17]), 
      .ZN(n_0_1_95));
   INV_X1 i_0_1_186 (.A(n_0_1_96), .ZN(n_0_248));
   AOI22_X1 i_0_1_187 (.A1(n_0_48), .A2(n_0_266), .B1(n_0_1_109), .B2(A[18]), 
      .ZN(n_0_1_96));
   INV_X1 i_0_1_188 (.A(n_0_1_97), .ZN(n_0_249));
   AOI22_X1 i_0_1_189 (.A1(n_0_49), .A2(n_0_266), .B1(n_0_1_109), .B2(A[19]), 
      .ZN(n_0_1_97));
   INV_X1 i_0_1_190 (.A(n_0_1_98), .ZN(n_0_250));
   AOI22_X1 i_0_1_191 (.A1(n_0_50), .A2(n_0_266), .B1(n_0_1_109), .B2(A[20]), 
      .ZN(n_0_1_98));
   INV_X1 i_0_1_192 (.A(n_0_1_99), .ZN(n_0_251));
   AOI22_X1 i_0_1_193 (.A1(n_0_51), .A2(n_0_266), .B1(n_0_1_109), .B2(A[21]), 
      .ZN(n_0_1_99));
   INV_X1 i_0_1_194 (.A(n_0_1_100), .ZN(n_0_252));
   AOI22_X1 i_0_1_195 (.A1(n_0_52), .A2(n_0_266), .B1(n_0_1_109), .B2(A[22]), 
      .ZN(n_0_1_100));
   INV_X1 i_0_1_196 (.A(n_0_1_101), .ZN(n_0_253));
   AOI22_X1 i_0_1_197 (.A1(n_0_53), .A2(n_0_266), .B1(n_0_1_109), .B2(A[23]), 
      .ZN(n_0_1_101));
   INV_X1 i_0_1_198 (.A(n_0_1_102), .ZN(n_0_254));
   AOI22_X1 i_0_1_199 (.A1(n_0_54), .A2(n_0_266), .B1(n_0_1_109), .B2(A[24]), 
      .ZN(n_0_1_102));
   INV_X1 i_0_1_200 (.A(n_0_1_103), .ZN(n_0_255));
   AOI22_X1 i_0_1_201 (.A1(n_0_55), .A2(n_0_266), .B1(n_0_1_109), .B2(A[25]), 
      .ZN(n_0_1_103));
   INV_X1 i_0_1_202 (.A(n_0_1_104), .ZN(n_0_256));
   AOI22_X1 i_0_1_203 (.A1(n_0_56), .A2(n_0_266), .B1(n_0_1_109), .B2(A[26]), 
      .ZN(n_0_1_104));
   INV_X1 i_0_1_204 (.A(n_0_1_105), .ZN(n_0_257));
   AOI22_X1 i_0_1_205 (.A1(n_0_57), .A2(n_0_266), .B1(n_0_1_109), .B2(A[27]), 
      .ZN(n_0_1_105));
   INV_X1 i_0_1_206 (.A(n_0_1_106), .ZN(n_0_258));
   AOI22_X1 i_0_1_207 (.A1(n_0_58), .A2(n_0_266), .B1(n_0_1_109), .B2(A[28]), 
      .ZN(n_0_1_106));
   INV_X1 i_0_1_208 (.A(n_0_1_107), .ZN(n_0_259));
   AOI22_X1 i_0_1_209 (.A1(n_0_59), .A2(n_0_266), .B1(n_0_1_109), .B2(A[29]), 
      .ZN(n_0_1_107));
   INV_X1 i_0_1_210 (.A(n_0_1_108), .ZN(n_0_260));
   AOI22_X1 i_0_1_211 (.A1(n_0_60), .A2(n_0_266), .B1(n_0_1_109), .B2(A[30]), 
      .ZN(n_0_1_108));
   NOR2_X1 i_0_1_212 (.A1(A[31]), .A2(reset), .ZN(n_0_1_109));
   AND2_X1 i_0_1_213 (.A1(n_0_61), .A2(n_0_266), .ZN(n_0_261));
   AND2_X1 i_0_1_214 (.A1(n_0_157), .A2(n_0_1_112), .ZN(n_0_263));
   NAND2_X1 i_0_1_215 (.A1(n_0_1_112), .A2(n_0_1_110), .ZN(n_0_264));
   NAND2_X1 i_0_1_216 (.A1(Res[0]), .A2(n_0_1_111), .ZN(n_0_1_110));
   AOI21_X1 i_0_1_217 (.A(ready), .B1(enable), .B2(clk), .ZN(n_0_1_111));
   INV_X1 i_0_1_218 (.A(n_0_1_112), .ZN(n_0_262));
   AND2_X1 i_0_1_219 (.A1(n_0_1_139), .A2(n_0_1_113), .ZN(n_0_1_112));
   NAND3_X1 i_0_1_220 (.A1(clk), .A2(ready), .A3(enable), .ZN(n_0_1_113));
   NAND2_X1 i_0_1_221 (.A1(clk), .A2(enable), .ZN(n_0_1_114));
   NOR2_X1 i_0_1_222 (.A1(n_0_1_141), .A2(reset), .ZN(n_0_265));
   AND2_X1 i_0_1_223 (.A1(n_0_1_139), .A2(A[31]), .ZN(n_0_266));
   XNOR2_X1 i_0_1_224 (.A(isNeg[0]), .B(n_0_1_115), .ZN(OVF));
   NAND2_X1 i_0_1_225 (.A1(n_0_1_140), .A2(Res[63]), .ZN(n_0_1_115));
   MUX2_X1 i_0_1_226 (.A(n_0_62), .B(multiplicand[1]), .S(n_0_1_116), .Z(Res[1]));
   MUX2_X1 i_0_1_227 (.A(n_0_63), .B(multiplicand[2]), .S(n_0_1_116), .Z(Res[2]));
   MUX2_X1 i_0_1_228 (.A(n_0_64), .B(multiplicand[3]), .S(n_0_1_116), .Z(Res[3]));
   MUX2_X1 i_0_1_229 (.A(n_0_65), .B(multiplicand[4]), .S(n_0_1_116), .Z(Res[4]));
   MUX2_X1 i_0_1_230 (.A(n_0_66), .B(multiplicand[5]), .S(n_0_1_116), .Z(Res[5]));
   MUX2_X1 i_0_1_231 (.A(n_0_67), .B(multiplicand[6]), .S(n_0_1_116), .Z(Res[6]));
   MUX2_X1 i_0_1_232 (.A(n_0_68), .B(multiplicand[7]), .S(n_0_1_116), .Z(Res[7]));
   MUX2_X1 i_0_1_233 (.A(n_0_69), .B(multiplicand[8]), .S(n_0_1_116), .Z(Res[8]));
   MUX2_X1 i_0_1_234 (.A(n_0_70), .B(multiplicand[9]), .S(n_0_1_116), .Z(Res[9]));
   MUX2_X1 i_0_1_235 (.A(n_0_71), .B(multiplicand[10]), .S(n_0_1_116), .Z(
      Res[10]));
   MUX2_X1 i_0_1_236 (.A(n_0_72), .B(multiplicand[11]), .S(n_0_1_116), .Z(
      Res[11]));
   MUX2_X1 i_0_1_237 (.A(n_0_73), .B(multiplicand[12]), .S(n_0_1_116), .Z(
      Res[12]));
   MUX2_X1 i_0_1_238 (.A(n_0_74), .B(multiplicand[13]), .S(n_0_1_116), .Z(
      Res[13]));
   MUX2_X1 i_0_1_239 (.A(n_0_75), .B(multiplicand[14]), .S(n_0_1_116), .Z(
      Res[14]));
   MUX2_X1 i_0_1_240 (.A(n_0_76), .B(multiplicand[15]), .S(n_0_1_116), .Z(
      Res[15]));
   MUX2_X1 i_0_1_241 (.A(n_0_77), .B(multiplicand[16]), .S(n_0_1_116), .Z(
      Res[16]));
   MUX2_X1 i_0_1_242 (.A(n_0_78), .B(multiplicand[17]), .S(n_0_1_116), .Z(
      Res[17]));
   MUX2_X1 i_0_1_243 (.A(n_0_79), .B(multiplicand[18]), .S(n_0_1_116), .Z(
      Res[18]));
   MUX2_X1 i_0_1_244 (.A(n_0_80), .B(multiplicand[19]), .S(n_0_1_116), .Z(
      Res[19]));
   MUX2_X1 i_0_1_245 (.A(n_0_81), .B(multiplicand[20]), .S(n_0_1_116), .Z(
      Res[20]));
   MUX2_X1 i_0_1_246 (.A(n_0_82), .B(multiplicand[21]), .S(n_0_1_116), .Z(
      Res[21]));
   MUX2_X1 i_0_1_247 (.A(n_0_83), .B(multiplicand[22]), .S(n_0_1_116), .Z(
      Res[22]));
   MUX2_X1 i_0_1_248 (.A(n_0_84), .B(multiplicand[23]), .S(n_0_1_116), .Z(
      Res[23]));
   MUX2_X1 i_0_1_249 (.A(n_0_85), .B(multiplicand[24]), .S(n_0_1_116), .Z(
      Res[24]));
   MUX2_X1 i_0_1_250 (.A(n_0_86), .B(multiplicand[25]), .S(n_0_1_116), .Z(
      Res[25]));
   MUX2_X1 i_0_1_251 (.A(n_0_87), .B(multiplicand[26]), .S(n_0_1_116), .Z(
      Res[26]));
   MUX2_X1 i_0_1_252 (.A(n_0_88), .B(multiplicand[27]), .S(n_0_1_116), .Z(
      Res[27]));
   MUX2_X1 i_0_1_253 (.A(n_0_89), .B(multiplicand[28]), .S(n_0_1_116), .Z(
      Res[28]));
   MUX2_X1 i_0_1_254 (.A(n_0_90), .B(multiplicand[29]), .S(n_0_1_116), .Z(
      Res[29]));
   MUX2_X1 i_0_1_255 (.A(n_0_91), .B(multiplicand[30]), .S(n_0_1_116), .Z(
      Res[30]));
   MUX2_X1 i_0_1_256 (.A(n_0_92), .B(multiplicand[31]), .S(n_0_1_116), .Z(
      Res[31]));
   MUX2_X1 i_0_1_257 (.A(n_0_93), .B(accumulator[0]), .S(n_0_1_116), .Z(Res[32]));
   MUX2_X1 i_0_1_258 (.A(n_0_94), .B(accumulator[1]), .S(n_0_1_116), .Z(Res[33]));
   MUX2_X1 i_0_1_259 (.A(n_0_95), .B(accumulator[2]), .S(n_0_1_116), .Z(Res[34]));
   MUX2_X1 i_0_1_260 (.A(n_0_96), .B(accumulator[3]), .S(n_0_1_116), .Z(Res[35]));
   MUX2_X1 i_0_1_261 (.A(n_0_97), .B(accumulator[4]), .S(n_0_1_116), .Z(Res[36]));
   MUX2_X1 i_0_1_262 (.A(n_0_98), .B(accumulator[5]), .S(n_0_1_116), .Z(Res[37]));
   MUX2_X1 i_0_1_263 (.A(n_0_99), .B(accumulator[6]), .S(n_0_1_116), .Z(Res[38]));
   MUX2_X1 i_0_1_264 (.A(n_0_100), .B(accumulator[7]), .S(n_0_1_116), .Z(Res[39]));
   MUX2_X1 i_0_1_265 (.A(n_0_101), .B(accumulator[8]), .S(n_0_1_116), .Z(Res[40]));
   MUX2_X1 i_0_1_266 (.A(n_0_102), .B(accumulator[9]), .S(n_0_1_116), .Z(Res[41]));
   MUX2_X1 i_0_1_267 (.A(n_0_103), .B(accumulator[10]), .S(n_0_1_116), .Z(
      Res[42]));
   MUX2_X1 i_0_1_268 (.A(n_0_104), .B(accumulator[11]), .S(n_0_1_116), .Z(
      Res[43]));
   MUX2_X1 i_0_1_269 (.A(n_0_105), .B(accumulator[12]), .S(n_0_1_116), .Z(
      Res[44]));
   MUX2_X1 i_0_1_270 (.A(n_0_106), .B(accumulator[13]), .S(n_0_1_116), .Z(
      Res[45]));
   MUX2_X1 i_0_1_271 (.A(n_0_107), .B(accumulator[14]), .S(n_0_1_116), .Z(
      Res[46]));
   MUX2_X1 i_0_1_272 (.A(n_0_108), .B(accumulator[15]), .S(n_0_1_116), .Z(
      Res[47]));
   MUX2_X1 i_0_1_273 (.A(n_0_109), .B(accumulator[16]), .S(n_0_1_116), .Z(
      Res[48]));
   MUX2_X1 i_0_1_274 (.A(n_0_110), .B(accumulator[17]), .S(n_0_1_116), .Z(
      Res[49]));
   MUX2_X1 i_0_1_275 (.A(n_0_111), .B(accumulator[18]), .S(n_0_1_116), .Z(
      Res[50]));
   MUX2_X1 i_0_1_276 (.A(n_0_112), .B(accumulator[19]), .S(n_0_1_116), .Z(
      Res[51]));
   MUX2_X1 i_0_1_277 (.A(n_0_113), .B(accumulator[20]), .S(n_0_1_116), .Z(
      Res[52]));
   MUX2_X1 i_0_1_278 (.A(n_0_114), .B(accumulator[21]), .S(n_0_1_116), .Z(
      Res[53]));
   MUX2_X1 i_0_1_279 (.A(n_0_115), .B(accumulator[22]), .S(n_0_1_116), .Z(
      Res[54]));
   MUX2_X1 i_0_1_280 (.A(n_0_116), .B(accumulator[23]), .S(n_0_1_116), .Z(
      Res[55]));
   MUX2_X1 i_0_1_281 (.A(n_0_117), .B(accumulator[24]), .S(n_0_1_116), .Z(
      Res[56]));
   MUX2_X1 i_0_1_282 (.A(n_0_118), .B(accumulator[25]), .S(n_0_1_116), .Z(
      Res[57]));
   MUX2_X1 i_0_1_283 (.A(n_0_119), .B(accumulator[26]), .S(n_0_1_116), .Z(
      Res[58]));
   MUX2_X1 i_0_1_284 (.A(n_0_120), .B(accumulator[27]), .S(n_0_1_116), .Z(
      Res[59]));
   MUX2_X1 i_0_1_285 (.A(n_0_121), .B(accumulator[28]), .S(n_0_1_116), .Z(
      Res[60]));
   MUX2_X1 i_0_1_286 (.A(n_0_122), .B(accumulator[29]), .S(n_0_1_116), .Z(
      Res[61]));
   MUX2_X1 i_0_1_287 (.A(n_0_123), .B(accumulator[30]), .S(n_0_1_116), .Z(
      Res[62]));
   MUX2_X1 i_0_1_288 (.A(n_0_124), .B(accumulator[31]), .S(n_0_1_116), .Z(
      Res[63]));
   OR2_X1 i_0_1_289 (.A1(n_0_1_118), .A2(n_0_1_117), .ZN(n_0_1_116));
   XNOR2_X1 i_0_1_290 (.A(isNeg[1]), .B(isNeg[0]), .ZN(n_0_1_117));
   NOR4_X1 i_0_1_291 (.A1(n_0_1_134), .A2(n_0_1_129), .A3(n_0_1_124), .A4(
      n_0_1_119), .ZN(n_0_1_118));
   NAND4_X1 i_0_1_292 (.A1(n_0_1_123), .A2(n_0_1_122), .A3(n_0_1_121), .A4(
      n_0_1_120), .ZN(n_0_1_119));
   NOR4_X1 i_0_1_293 (.A1(multiplicand[12]), .A2(multiplicand[11]), .A3(
      multiplicand[10]), .A4(multiplicand[9]), .ZN(n_0_1_120));
   NOR4_X1 i_0_1_294 (.A1(multiplicand[14]), .A2(multiplicand[13]), .A3(
      multiplicand[8]), .A4(Res[0]), .ZN(n_0_1_121));
   NOR4_X1 i_0_1_295 (.A1(multiplicand[4]), .A2(multiplicand[3]), .A3(
      multiplicand[2]), .A4(multiplicand[1]), .ZN(n_0_1_122));
   NOR4_X1 i_0_1_296 (.A1(multiplicand[15]), .A2(multiplicand[7]), .A3(
      multiplicand[6]), .A4(multiplicand[5]), .ZN(n_0_1_123));
   NAND4_X1 i_0_1_297 (.A1(n_0_1_128), .A2(n_0_1_127), .A3(n_0_1_126), .A4(
      n_0_1_125), .ZN(n_0_1_124));
   NOR4_X1 i_0_1_298 (.A1(multiplicand[28]), .A2(multiplicand[27]), .A3(
      multiplicand[26]), .A4(multiplicand[25]), .ZN(n_0_1_125));
   NOR4_X1 i_0_1_299 (.A1(multiplicand[31]), .A2(multiplicand[30]), .A3(
      multiplicand[29]), .A4(multiplicand[24]), .ZN(n_0_1_126));
   NOR4_X1 i_0_1_300 (.A1(multiplicand[20]), .A2(multiplicand[19]), .A3(
      multiplicand[18]), .A4(multiplicand[17]), .ZN(n_0_1_127));
   NOR4_X1 i_0_1_301 (.A1(multiplicand[23]), .A2(multiplicand[22]), .A3(
      multiplicand[21]), .A4(multiplicand[16]), .ZN(n_0_1_128));
   NAND4_X1 i_0_1_302 (.A1(n_0_1_133), .A2(n_0_1_132), .A3(n_0_1_131), .A4(
      n_0_1_130), .ZN(n_0_1_129));
   NOR4_X1 i_0_1_303 (.A1(accumulator[12]), .A2(accumulator[11]), .A3(
      accumulator[10]), .A4(accumulator[9]), .ZN(n_0_1_130));
   NOR4_X1 i_0_1_304 (.A1(accumulator[15]), .A2(accumulator[14]), .A3(
      accumulator[13]), .A4(accumulator[8]), .ZN(n_0_1_131));
   NOR4_X1 i_0_1_305 (.A1(accumulator[4]), .A2(accumulator[3]), .A3(
      accumulator[2]), .A4(accumulator[1]), .ZN(n_0_1_132));
   NOR4_X1 i_0_1_306 (.A1(accumulator[16]), .A2(accumulator[7]), .A3(
      accumulator[6]), .A4(accumulator[5]), .ZN(n_0_1_133));
   NAND4_X1 i_0_1_307 (.A1(n_0_1_138), .A2(n_0_1_137), .A3(n_0_1_136), .A4(
      n_0_1_135), .ZN(n_0_1_134));
   NOR4_X1 i_0_1_308 (.A1(accumulator[29]), .A2(accumulator[28]), .A3(
      accumulator[27]), .A4(accumulator[26]), .ZN(n_0_1_135));
   NOR4_X1 i_0_1_309 (.A1(accumulator[31]), .A2(accumulator[30]), .A3(
      accumulator[25]), .A4(accumulator[0]), .ZN(n_0_1_136));
   NOR4_X1 i_0_1_310 (.A1(accumulator[21]), .A2(accumulator[20]), .A3(
      accumulator[19]), .A4(accumulator[18]), .ZN(n_0_1_137));
   NOR4_X1 i_0_1_311 (.A1(accumulator[24]), .A2(accumulator[23]), .A3(
      accumulator[22]), .A4(accumulator[17]), .ZN(n_0_1_138));
   INV_X1 i_0_1_312 (.A(reset), .ZN(n_0_1_139));
   INV_X1 i_0_1_313 (.A(isNeg[1]), .ZN(n_0_1_140));
   INV_X1 i_0_1_314 (.A(B[31]), .ZN(n_0_1_141));
   INV_X1 i_0_1_315 (.A(counter[4]), .ZN(n_0_1_142));
endmodule
