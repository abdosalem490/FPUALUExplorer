* SPICE NETLIST
***************************************

.SUBCKT MGC_via1_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X2
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_3
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2_X1 A2 VSS A1 ZN VDD 6 7
** N=8 EP=7 IP=0 FDC=4
M0 8 A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN A1 8 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A2 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A1 ZN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2_X1 A1 A2 VSS VDD ZN 6 7
** N=9 EP=7 IP=0 FDC=6
M0 8 A1 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 9 A1 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 9 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT via1_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT OAI22_X1 B2 B1 VSS ZN A1 A2 VDD 8 9
** N=12 EP=9 IP=0 FDC=8
M0 VSS B2 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 10 B1 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A1 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 10 A2 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 11 B2 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 ZN B1 11 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 12 A1 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 VDD A2 12 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NAND4_X1 A4 VSS A3 A2 A1 ZN VDD 8 9
** N=12 EP=9 IP=0 FDC=8
M0 10 A4 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 11 A3 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 12 A2 11 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A1 12 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN A4 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 VDD A3 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 ZN A2 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 VDD A1 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FILLCELL_X4
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_12
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT XOR2_X1 VDD A Z B VSS 6 7
** N=11 EP=7 IP=0 FDC=10
M0 8 A VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 11 A Z 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 11 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 10 A 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 10 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 9 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 9 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 9 B Z 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XNOR2_X1 VSS A ZN B VDD 6 7
** N=11 EP=7 IP=0 FDC=10
M0 11 A 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=155 $Y=90 $D=1
M1 VSS B 11 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=345 $Y=90 $D=1
M2 9 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=540 $Y=90 $D=1
M3 ZN A 9 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 9 B ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 8 A VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=155 $Y=995 $D=0
M6 VDD B 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=345 $Y=995 $D=0
M7 ZN 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=540 $Y=680 $D=0
M8 10 A ZN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M9 VDD B 10 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT INV_X1 A VSS VDD ZN 5 6
** N=6 EP=6 IP=0 FDC=2
M0 ZN A VSS 5 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN A VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=2
X1 3 1 2 4 5 6 INV_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT OAI221_X1 B2 B1 VSS A C2 VDD C1 ZN 9 10
** N=14 EP=10 IP=0 FDC=10
M0 VSS B2 11 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 11 B1 VSS 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 12 A 11 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN C2 12 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 12 C1 ZN 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 13 B2 VDD 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 ZN B1 13 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 VDD A ZN 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 14 C2 VDD 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 ZN C1 14 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X8
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_17
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4 5 6 7 8 9 10 11 12 13 14
** N=14 EP=14 IP=18 FDC=16
X0 1 2 3 4 5 6 7 13 14 OAI22_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 8 9 3 10 11 12 7 13 14 OAI22_X1 $T=950 0 0 0 $X=835 $Y=-115
.ENDS
***************************************
.SUBCKT OAI21_X1 B2 B1 ZN A VSS VDD 7 8
** N=10 EP=8 IP=0 FDC=6
M0 ZN B2 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 9 B1 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS A 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=550 $Y=90 $D=1
M3 10 B2 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M4 ZN B1 10 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M5 VDD A ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=550 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=13 FDC=8
X0 1 2 3 4 5 6 7 8 9 OAI22_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_22
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=13 FDC=8
X1 3 4 1 5 6 7 2 8 9 OAI22_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_24
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_25
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_26
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT HA_X1 S B A VSS VDD CO 7 8
** N=14 EP=8 IP=0 FDC=16
M0 13 B VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 S A 13 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS 10 S 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.48e-14 AS=5.81e-14 PD=1.12e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 10 B VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.48e-14 PD=7e-07 PS=1.12e-06 $X=760 $Y=90 $D=1
M4 VSS A 10 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=950 $Y=90 $D=1
M5 14 A 11 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1320 $Y=90 $D=1
M6 VSS B 14 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=1510 $Y=90 $D=1
M7 CO 11 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1700 $Y=90 $D=1
M8 S B 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M9 9 A S 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M10 VDD 10 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.7725e-14 AS=8.82e-14 PD=1.55e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M11 12 B VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.7725e-14 PD=9.1e-07 PS=1.55e-06 $X=760 $Y=870 $D=0
M12 10 A 12 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=950 $Y=870 $D=0
M13 11 A VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1320 $Y=870 $D=0
M14 VDD B 11 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=1510 $Y=870 $D=0
M15 CO 11 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1700 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=2
X1 3 1 2 4 5 6 INV_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_28
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT AOI21_X1 B2 B1 ZN A VSS VDD 7 8
** N=10 EP=8 IP=0 FDC=6
M0 10 B2 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN B1 10 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS A ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B2 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M4 9 B1 ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M5 VDD A 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR2_X1 A2 VDD A1 ZN VSS 6 7
** N=8 EP=7 IP=0 FDC=4
M0 ZN A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A1 ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 8 A2 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 ZN A1 8 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FA_X1 CO CI B A VDD VSS S 8 9
** N=21 EP=9 IP=0 FDC=28
M0 VSS 10 CO 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 19 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06 $X=360 $Y=215 $D=1
M2 10 A 19 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=550 $Y=215 $D=1
M3 11 CI 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07 $X=740 $Y=215 $D=1
M4 VSS A 11 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07 $X=935 $Y=215 $D=1
M5 11 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1125 $Y=215 $D=1
M6 13 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1465 $Y=90 $D=1
M7 VSS CI 13 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1655 $Y=90 $D=1
M8 13 A VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1845 $Y=90 $D=1
M9 15 10 13 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07 $X=2035 $Y=90 $D=1
M10 20 CI 15 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.15e-14 PD=7e-07 PS=7.2e-07 $X=2235 $Y=90 $D=1
M11 21 B 20 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2425 $Y=90 $D=1
M12 VSS A 21 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=2615 $Y=90 $D=1
M13 S 15 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=2805 $Y=90 $D=1
M14 VDD 10 CO 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M15 16 B VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.54e-06 $X=360 $Y=870 $D=0
M16 10 A 16 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=550 $Y=870 $D=0
M17 12 CI 10 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06 PS=9.1e-07 $X=740 $Y=870 $D=0
M18 VDD A 12 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.53e-14 PD=9.1e-07 PS=1.07e-06 $X=935 $Y=945 $D=0
M19 12 B VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1125 $Y=945 $D=0
M20 14 B VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1465 $Y=995 $D=0
M21 VDD CI 14 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1655 $Y=995 $D=0
M22 14 A VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1845 $Y=995 $D=0
M23 15 10 14 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07 $X=2035 $Y=995 $D=0
M24 17 CI 15 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.725e-14 PD=9.1e-07 PS=9.3e-07 $X=2235 $Y=995 $D=0
M25 18 B 17 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=2425 $Y=995 $D=0
M26 VDD A 18 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2615 $Y=995 $D=0
M27 S 15 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2805 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_29
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT AOI22_X1 B2 B1 VDD A1 ZN A2 VSS 8 9
** N=12 EP=9 IP=0 FDC=8
M0 11 B2 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN B1 11 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 12 A1 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 VSS A2 12 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 VDD B2 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 10 B1 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 ZN A1 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 10 A2 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OR4_X1 A1 A2 A3 A4 VSS VDD ZN 8 9
** N=13 EP=9 IP=0 FDC=10
M0 10 A1 VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 10 A3 VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 VSS A4 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=715 $Y=90 $D=1
M4 ZN 10 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 11 A1 10 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 12 A2 11 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 13 A3 12 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M8 VDD A4 13 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=715 $Y=995 $D=0
M9 ZN 10 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_30
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_31
** N=3 EP=0 IP=3 FDC=0
.ENDS
***************************************
.SUBCKT ICV_32
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_33
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_34
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_35 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=4
X0 1 2 3 4 7 8 INV_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 5 2 3 6 7 8 INV_X1 $T=380 0 0 0 $X=265 $Y=-115
.ENDS
***************************************
.SUBCKT FILLCELL_X16
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_36
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_37
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_38 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=2
X1 3 1 2 4 5 6 INV_X1 $T=760 0 0 0 $X=645 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_39 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=15 FDC=10
X0 1 2 3 4 5 6 7 10 11 OAI22_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 8 3 7 9 10 11 INV_X1 $T=950 0 0 0 $X=835 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_40
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_41
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_42
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via1_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2_X2 A1 ZN A2 VSS VDD 6 7
** N=9 EP=7 IP=0 FDC=8
M0 ZN A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A1 ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 ZN A1 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS A2 ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 8 A2 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN A1 8 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 9 A1 ZN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 VDD A2 9 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_43
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_44
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT NAND3_X1 A3 VSS A2 A1 VDD ZN 7 8
** N=10 EP=8 IP=0 FDC=6
M0 9 A3 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 10 A2 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 10 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A3 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 VDD A2 ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI33_X1 B3 B2 B1 VSS A1 A2 A3 ZN VDD 10 11
** N=16 EP=11 IP=0 FDC=12
M0 12 B3 VSS 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS B2 12 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 12 B1 VSS 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 ZN A1 12 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 12 A2 ZN 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 ZN A3 12 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1110 $Y=90 $D=1
M6 13 B3 VDD 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M7 14 B2 13 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M8 ZN B1 14 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M9 15 A1 ZN 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M10 16 A2 15 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
M11 VDD A3 16 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1110 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_45 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=6
X1 3 5 4 6 1 2 7 8 OAI21_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI222_X1 C2 C1 VSS B1 B2 A2 VDD A1 ZN 10 11
** N=16 EP=11 IP=0 FDC=12
M0 12 C2 VSS 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=155 $Y=90 $D=1
M1 VSS C1 12 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=345 $Y=90 $D=1
M2 12 B1 13 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=710 $Y=90 $D=1
M3 13 B2 12 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=900 $Y=90 $D=1
M4 ZN A2 13 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1090 $Y=90 $D=1
M5 13 A1 ZN 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1280 $Y=90 $D=1
M6 14 C2 VDD 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=155 $Y=680 $D=0
M7 ZN C1 14 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=1.9845e-13 AS=8.82e-14 PD=1.89e-06 PS=1.54e-06 $X=345 $Y=680 $D=0
M8 15 B1 ZN 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.9845e-13 PD=1.54e-06 PS=1.89e-06 $X=710 $Y=680 $D=0
M9 VDD B2 15 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=900 $Y=680 $D=0
M10 16 A2 VDD 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1090 $Y=680 $D=0
M11 ZN A1 16 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1280 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI21_X2 A VDD B1 ZN B2 VSS 7 8
** N=11 EP=8 IP=0 FDC=12
M0 ZN A VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 10 B2 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B1 10 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 11 B1 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=945 $Y=90 $D=1
M5 VSS B2 11 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1135 $Y=90 $D=1
M6 VDD A 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M7 9 A VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M8 ZN B2 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M9 9 B1 ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
M10 ZN B1 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=945 $Y=680 $D=0
M11 9 B2 ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1135 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_46
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X32
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT NOR3_X1 A3 VDD A2 A1 VSS ZN 7 8
** N=10 EP=8 IP=0 FDC=6
M0 ZN A3 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A2 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 9 A3 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 10 A2 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 10 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI211_X1 C2 C1 A VDD B ZN VSS 8 9
** N=12 EP=9 IP=0 FDC=8
M0 ZN C2 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 10 C1 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 12 A 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS B 12 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 11 C2 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN C1 11 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 VDD A ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 ZN B VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_47
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT AND2_X1 A1 A2 VSS VDD ZN 6 7
** N=9 EP=7 IP=0 FDC=6
M0 9 A1 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 9 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 8 A1 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OR3_X1 A1 A2 A3 VSS VDD ZN 7 8
** N=11 EP=8 IP=0 FDC=8
M0 VSS A1 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 9 A2 VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 VSS A3 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=525 $Y=90 $D=1
M3 ZN 9 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 10 A1 9 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M5 11 A2 10 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M6 VDD A3 11 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=525 $Y=995 $D=0
M7 ZN 9 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT CLKBUF_X2 A Z VSS VDD 5 6
** N=7 EP=6 IP=0 FDC=6
M0 VSS A 7 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07 $X=145 $Y=90 $D=1
M1 Z 7 VSS 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=335 $Y=90 $D=1
M2 VSS 7 Z 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=525 $Y=90 $D=1
M3 VDD A 7 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 Z 7 VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 VDD 7 Z 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_48 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=16 FDC=18
X0 1 2 3 4 5 6 7 11 12 OAI22_X1 $T=1140 0 0 0 $X=1025 $Y=-115
X1 7 8 9 10 3 11 12 XOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_49
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI221_X1 B2 B1 VDD A C2 VSS C1 ZN 9 10
** N=14 EP=10 IP=0 FDC=10
M0 13 B2 VSS 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN B1 13 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 VSS A ZN 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 14 C2 VSS 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN C1 14 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 VDD B2 11 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 11 B1 VDD 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 12 A 11 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 ZN C2 12 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 12 C1 ZN 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FPU_VA B[31] A[31] B[24] A[25] A[27] A[23] B[28] B[30] A[30] A[20] A[4] B[15] B[26] SUM[19] SUM[15] B[27] SUM[6] A[28] SUM[3] B[16]
+ B[13] B[12] B[10] B[21] B[19] B[8] A[8] A[19] A[11] B[11] A[15] B[0] B[7] B[20] SUM[31] SUM[13] SUM[22] B[29] SUM[4] B[23]
+ SUM[8] B[25] SUM[10] SUM[7] SUM[5] A[29] B[17] B[14] A[16] A[13] A[18] A[14] A[12] B[18] A[22] B[2] B[1] A[9] A[21] A[7]
+ B[6] B[4] A[26] SUM[20] SUM[24] SUM[2] SUM[28] A[24] A[17] B[22] A[10] B[9] A[5] A[6] SUM[21] A[1] SUM[18] SUM[17] SUM[23] SUM[9]
+ SUM[12] SUM[14] SUM[16] A[2] A[0] A[3] B[5] B[3] SUM[26] SUM[27] SUM[11] SUM[25] SUM[29] SUM[30] SUM[0] SUM[1]
** N=1029 EP=96 IP=15994 FDC=6266
M0 299 316 31 998 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.03e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07 $X=14085 $Y=43160 $D=1
M1 316 10 299 998 NMOS_VTL L=5e-08 W=9.5e-08 AD=9.975e-15 AS=2.03e-14 PD=4e-07 PS=6.7e-07 $X=14275 $Y=43160 $D=1
M2 991 158 323 999 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=27555 $Y=6300 $D=1
M3 992 172 991 999 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=27745 $Y=6300 $D=1
M4 993 253 992 999 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=27935 $Y=6300 $D=1
M5 299 154 993 999 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=28125 $Y=6300 $D=1
M6 324 323 299 999 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=28315 $Y=6095 $D=1
M7 994 325 299 1000 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=28735 $Y=9490 $D=1
M8 329 174 994 1000 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=28925 $Y=9490 $D=1
M9 299 176 329 1000 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=29115 $Y=9490 $D=1
M10 329 328 299 1000 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=29305 $Y=9490 $D=1
M11 299 10 337 998 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07 $X=31925 $Y=42700 $D=1
M12 338 337 299 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=32115 $Y=42495 $D=1
M13 995 340 299 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=34585 $Y=40290 $D=1
M14 343 236 995 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=1.2035e-13 AS=5.81e-14 PD=1.41e-06 PS=1.11e-06 $X=34775 $Y=40290 $D=1
M15 996 B[28] 343 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=1.2035e-13 PD=1.11e-06 PS=1.41e-06 $X=35115 $Y=40290 $D=1
M16 299 240 996 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=35305 $Y=40290 $D=1
M17 997 242 299 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=35495 $Y=40290 $D=1
M18 343 B[27] 997 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=35685 $Y=40290 $D=1
M19 299 346 348 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=37245 $Y=43090 $D=1
M20 348 346 299 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37435 $Y=43090 $D=1
M21 299 346 348 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37625 $Y=43090 $D=1
M22 348 346 299 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37815 $Y=43090 $D=1
M23 10 351 348 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38005 $Y=43090 $D=1
M24 348 B[30] 10 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38195 $Y=43090 $D=1
M25 10 B[30] 348 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38385 $Y=43090 $D=1
M26 348 351 10 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38575 $Y=43090 $D=1
M27 10 351 348 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38765 $Y=43090 $D=1
M28 348 B[30] 10 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38955 $Y=43090 $D=1
M29 10 B[30] 348 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=39145 $Y=43090 $D=1
M30 348 351 10 998 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=39335 $Y=43090 $D=1
M31 4 357 299 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=42565 $Y=40290 $D=1
M32 299 357 4 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=42755 $Y=40290 $D=1
M33 4 357 299 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=42945 $Y=40290 $D=1
M34 299 357 4 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43135 $Y=40290 $D=1
M35 4 360 299 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43325 $Y=40290 $D=1
M36 299 360 4 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43515 $Y=40290 $D=1
M37 4 360 299 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43705 $Y=40290 $D=1
M38 299 360 4 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=43895 $Y=40290 $D=1
M39 4 363 299 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=44270 $Y=40290 $D=1
M40 299 363 4 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=44460 $Y=40290 $D=1
M41 4 363 299 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=44650 $Y=40290 $D=1
M42 299 363 4 1001 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=44840 $Y=40290 $D=1
M43 300 316 31 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=14085 $Y=43680 $D=0
M44 316 10 300 1014 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=6.615e-14 PD=8.4e-07 PS=1.54e-06 $X=14275 $Y=43995 $D=0
M45 323 158 300 1015 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=27555 $Y=5290 $D=0
M46 300 172 323 1015 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=27745 $Y=5290 $D=0
M47 323 253 300 1015 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=27935 $Y=5290 $D=0
M48 300 154 323 1015 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=28125 $Y=5290 $D=0
M49 324 323 300 1015 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=28315 $Y=5290 $D=0
M50 329 325 327 1016 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=28735 $Y=10080 $D=0
M51 327 174 329 1016 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=28925 $Y=10080 $D=0
M52 986 176 327 1016 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=29115 $Y=10080 $D=0
M53 300 328 986 1016 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=29305 $Y=10080 $D=0
M54 300 10 337 1017 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=31925 $Y=41690 $D=0
M55 338 337 300 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=32115 $Y=41690 $D=0
M56 341 340 300 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=34585 $Y=40880 $D=0
M57 300 236 341 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=34775 $Y=40880 $D=0
M58 341 B[28] 344 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=35115 $Y=40880 $D=0
M59 344 240 341 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=35305 $Y=40880 $D=0
M60 343 242 344 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=35495 $Y=40880 $D=0
M61 344 B[27] 343 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=35685 $Y=40880 $D=0
M62 10 346 300 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=37245 $Y=43680 $D=0
M63 300 346 10 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37435 $Y=43680 $D=0
M64 10 346 300 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37625 $Y=43680 $D=0
M65 300 346 10 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37815 $Y=43680 $D=0
M66 987 351 300 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38005 $Y=43680 $D=0
M67 10 B[30] 987 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38195 $Y=43680 $D=0
M68 988 B[30] 10 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38385 $Y=43680 $D=0
M69 300 351 988 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38575 $Y=43680 $D=0
M70 989 351 300 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38765 $Y=43680 $D=0
M71 10 B[30] 989 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38955 $Y=43680 $D=0
M72 990 B[30] 10 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=39145 $Y=43680 $D=0
M73 300 351 990 1014 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=39335 $Y=43680 $D=0
M74 4 357 361 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=42565 $Y=40880 $D=0
M75 361 357 4 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=42755 $Y=40880 $D=0
M76 4 357 361 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=42945 $Y=40880 $D=0
M77 361 357 4 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43135 $Y=40880 $D=0
M78 364 360 361 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43325 $Y=40880 $D=0
M79 361 360 364 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43515 $Y=40880 $D=0
M80 364 360 361 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43705 $Y=40880 $D=0
M81 361 360 364 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=43895 $Y=40880 $D=0
M82 364 363 300 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=44270 $Y=40880 $D=0
M83 300 363 364 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=44460 $Y=40880 $D=0
M84 364 363 300 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=44650 $Y=40880 $D=0
M85 300 363 364 1017 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=44840 $Y=40880 $D=0
X5849 881 299 303 882 300 1007 1028 NAND2_X1 $T=2140 15000 1 0 $X=2025 $Y=13485
X5850 654 299 2 656 300 1010 1029 NAND2_X1 $T=2140 20600 0 0 $X=2025 $Y=20485
X5851 828 299 29 674 300 999 1020 NAND2_X1 $T=5180 6600 0 0 $X=5065 $Y=6485
X5852 414 299 44 885 300 1004 1025 NAND2_X1 $T=7650 26200 1 0 $X=7535 $Y=24685
X5853 52 299 405 386 300 1011 1026 NAND2_X1 $T=8030 31800 1 0 $X=7915 $Y=30285
X5854 427 299 58 836 300 1011 1026 NAND2_X1 $T=12780 31800 1 0 $X=12665 $Y=30285
X5855 85 299 71 18 300 1001 1017 NAND2_X1 $T=13730 40200 0 0 $X=13615 $Y=40085
X5856 712 299 65 464 300 1009 1024 NAND2_X1 $T=14110 1000 0 0 $X=13995 $Y=885
X5857 491 299 499 900 300 1000 1020 NAND2_X1 $T=19810 9400 1 0 $X=19695 $Y=7885
X5858 493 299 114 490 300 999 1015 NAND2_X1 $T=20000 6600 1 0 $X=19885 $Y=5085
X5859 321 299 127 902 300 1007 1028 NAND2_X1 $T=21140 15000 1 0 $X=21025 $Y=13485
X5860 154 299 245 530 300 1000 1020 NAND2_X1 $T=26650 9400 1 0 $X=26535 $Y=7885
X5861 253 299 209 162 300 1003 1016 NAND2_X1 $T=26650 12200 1 0 $X=26535 $Y=10685
X5862 172 299 185 163 300 1003 1028 NAND2_X1 $T=27980 12200 0 0 $X=27865 $Y=12085
X5863 233 299 286 191 300 1007 1028 NAND2_X1 $T=29500 15000 1 0 $X=29385 $Y=13485
X5864 559 299 561 262 300 1010 1021 NAND2_X1 $T=31970 20600 1 0 $X=31855 $Y=19085
X5865 220 299 770 219 300 1004 1019 NAND2_X1 $T=32920 26200 0 0 $X=32805 $Y=26085
X5866 207 299 214 564 300 1000 1020 NAND2_X1 $T=33110 9400 1 0 $X=32995 $Y=7885
X5867 261 299 262 224 300 1007 1028 NAND2_X1 $T=34440 15000 1 0 $X=34325 $Y=13485
X5868 218 299 582 263 300 1013 1029 NAND2_X1 $T=35770 23400 1 0 $X=35655 $Y=21885
X5869 784 299 241 352 300 1010 1021 NAND2_X1 $T=36910 20600 1 0 $X=36795 $Y=19085
X5870 872 299 597 SUM[27] 300 1008 1026 NAND2_X1 $T=37100 29000 0 0 $X=36985 $Y=28885
X5871 258 299 597 SUM[26] 300 1011 1018 NAND2_X1 $T=37480 31800 0 0 $X=37365 $Y=31685
X5872 259 299 597 SUM[25] 300 1002 1018 NAND2_X1 $T=37480 34600 1 0 $X=37365 $Y=33085
X5873 260 299 597 SUM[24] 300 1011 1026 NAND2_X1 $T=38810 31800 1 0 $X=38695 $Y=30285
X5874 214 299 251 607 300 1000 1020 NAND2_X1 $T=39950 9400 1 0 $X=39835 $Y=7885
X5875 279 299 597 SUM[23] 300 1004 1019 NAND2_X1 $T=40520 26200 0 0 $X=40405 $Y=26085
X5876 214 299 241 595 300 999 1020 NAND2_X1 $T=40710 6600 0 0 $X=40595 $Y=6485
X5877 214 299 246 627 300 999 1020 NAND2_X1 $T=42420 6600 0 0 $X=42305 $Y=6485
X5878 214 299 228 806 300 1000 1020 NAND2_X1 $T=42420 9400 1 0 $X=42305 $Y=7885
X5879 280 299 597 SUM[29] 300 1011 1026 NAND2_X1 $T=42610 31800 1 0 $X=42495 $Y=30285
X5880 281 299 597 SUM[28] 300 1008 1019 NAND2_X1 $T=42800 29000 1 0 $X=42685 $Y=27485
X5881 597 299 801 SUM[30] 300 1008 1026 NAND2_X1 $T=43370 29000 0 0 $X=43255 $Y=28885
X5882 A[30] 299 B[30] 642 300 998 1014 NAND2_X1 $T=44510 43000 0 0 $X=44395 $Y=42885
X6064 656 9 299 300 660 1010 1021 OR2_X1 $T=2330 20600 1 0 $X=2215 $Y=19085
X6065 882 11 299 300 385 1003 1028 OR2_X1 $T=2520 12200 0 0 $X=2405 $Y=12085
X6066 674 15 299 300 673 999 1015 OR2_X1 $T=4990 6600 1 0 $X=4875 $Y=5085
X6067 660 27 299 300 36 1010 1021 OR2_X1 $T=5750 20600 1 0 $X=5635 $Y=19085
X6068 885 30 299 300 829 1013 1025 OR2_X1 $T=5940 23400 0 0 $X=5825 $Y=23285
X6069 449 60 299 300 447 1002 1022 OR2_X1 $T=12590 34600 0 0 $X=12475 $Y=34485
X6070 715 84 299 300 80 1008 1019 OR2_X1 $T=15250 29000 1 0 $X=15135 $Y=27485
X6071 464 86 299 300 456 1012 1024 OR2_X1 $T=15440 3800 1 0 $X=15325 $Y=2285
X6072 421 87 299 300 473 1000 1016 OR2_X1 $T=15440 9400 0 0 $X=15325 $Y=9285
X6073 503 101 299 300 68 1010 1029 OR2_X1 $T=18100 20600 0 0 $X=17985 $Y=20485
X6074 903 107 299 300 100 1011 1018 OR2_X1 $T=19430 31800 0 0 $X=19315 $Y=31685
X6075 490 113 299 300 500 1012 1024 OR2_X1 $T=20570 3800 1 0 $X=20455 $Y=2285
X6076 732 115 299 300 903 1002 1018 OR2_X1 $T=20760 34600 1 0 $X=20645 $Y=33085
X6077 500 120 299 300 131 1012 1024 OR2_X1 $T=21330 3800 1 0 $X=21215 $Y=2285
X6078 133 135 299 300 116 1010 1021 OR2_X1 $T=24180 20600 1 0 $X=24065 $Y=19085
X6079 515 136 299 300 118 1013 1025 OR2_X1 $T=24180 23400 0 0 $X=24065 $Y=23285
X6080 SUM[31] 137 299 300 525 1007 1028 OR2_X1 $T=24370 15000 1 0 $X=24255 $Y=13485
X6081 165 143 299 300 153 1005 1023 OR2_X1 $T=24940 17800 1 0 $X=24825 $Y=16285
X6082 155 147 299 300 156 1007 1023 OR2_X1 $T=25510 15000 0 0 $X=25395 $Y=14885
X6083 534 160 299 300 515 1004 1019 OR2_X1 $T=27220 26200 0 0 $X=27105 $Y=26085
X6084 753 166 299 300 141 1013 1029 OR2_X1 $T=27790 23400 1 0 $X=27675 $Y=21885
X6085 326 177 299 300 753 1013 1025 OR2_X1 $T=28930 23400 0 0 $X=28815 $Y=23285
X6086 554 198 299 300 951 1010 1029 OR2_X1 $T=31020 20600 0 0 $X=30905 $Y=20485
X6087 262 207 299 300 222 1007 1028 OR2_X1 $T=32730 15000 1 0 $X=32615 $Y=13485
X6088 854 235 299 300 229 1013 1025 OR2_X1 $T=34630 23400 0 0 $X=34515 $Y=23285
X6089 241 257 299 300 592 1010 1021 OR2_X1 $T=37480 20600 1 0 $X=37365 $Y=19085
X6090 241 266 299 300 958 1005 1021 OR2_X1 $T=39000 17800 0 0 $X=38885 $Y=17685
X6091 632 269 299 300 272 1004 1025 OR2_X1 $T=39380 26200 1 0 $X=39265 $Y=24685
X6092 263 272 299 300 349 1004 1025 OR2_X1 $T=40140 26200 1 0 $X=40025 $Y=24685
X6093 B[30] A[30] 299 300 289 1006 1022 OR2_X1 $T=44320 37400 1 0 $X=44205 $Y=35885
X7250 302 421 299 662 B[31] 819 300 1003 1016 OAI22_X1 $T=3090 12200 1 0 $X=2975 $Y=10685
X7251 954 421 299 383 B[31] 301 300 1005 1023 OAI22_X1 $T=3280 17800 1 0 $X=3165 $Y=16285
X7252 653 A[31] 299 664 472 661 300 1005 1021 OAI22_X1 $T=3280 17800 0 0 $X=3165 $Y=17685
X7253 663 421 299 394 B[31] 369 300 999 1020 OAI22_X1 $T=3660 6600 0 0 $X=3545 $Y=6485
X7254 820 A[31] 299 389 472 665 300 1004 1025 OAI22_X1 $T=4040 26200 1 0 $X=3925 $Y=24685
X7255 667 405 299 6 58 883 300 1011 1018 OAI22_X1 $T=4040 31800 0 0 $X=3925 $Y=31685
X7256 373 A[31] 299 670 472 676 300 1010 1029 OAI22_X1 $T=4230 20600 0 0 $X=4115 $Y=20485
X7257 825 A[31] 299 409 472 671 300 1013 1029 OAI22_X1 $T=4800 23400 1 0 $X=4685 $Y=21885
X7258 392 677 299 395 35 45 300 1006 1022 OAI22_X1 $T=4990 37400 1 0 $X=4875 $Y=35885
X7259 824 421 299 407 B[31] 393 300 1012 1015 OAI22_X1 $T=5180 3800 0 0 $X=5065 $Y=3685
X7260 25 421 299 933 B[31] 15 300 999 1015 OAI22_X1 $T=5750 6600 1 0 $X=5635 $Y=5085
X7261 386 399 299 28 405 398 300 1011 1026 OAI22_X1 $T=5940 31800 1 0 $X=5825 $Y=30285
X7262 45 372 299 442 677 23 300 1006 1027 OAI22_X1 $T=5940 37400 0 0 $X=5825 $Y=37285
X7263 682 421 299 698 B[31] 307 300 1009 1024 OAI22_X1 $T=6320 1000 0 0 $X=6205 $Y=885
X7264 402 421 299 686 B[31] 306 300 1005 1023 OAI22_X1 $T=6510 17800 1 0 $X=6395 $Y=16285
X7265 305 A[31] 299 408 472 961 300 1005 1021 OAI22_X1 $T=6700 17800 0 0 $X=6585 $Y=17685
X7266 687 677 299 309 399 45 300 1006 1027 OAI22_X1 $T=6890 37400 0 0 $X=6775 $Y=37285
X7267 403 A[31] 299 690 472 308 300 1013 1025 OAI22_X1 $T=7080 23400 0 0 $X=6965 $Y=23285
X7268 888 696 299 700 17 401 300 1001 1017 OAI22_X1 $T=8980 40200 0 0 $X=8865 $Y=40085
X7269 411 A[31] 299 702 472 891 300 1010 1029 OAI22_X1 $T=9360 20600 0 0 $X=9245 $Y=20485
X7270 416 A[31] 299 51 472 890 300 1013 1025 OAI22_X1 $T=9360 23400 0 0 $X=9245 $Y=23285
X7271 10 310 299 429 834 298 300 1005 1021 OAI22_X1 $T=10500 17800 0 0 $X=10385 $Y=17685
X7272 705 677 299 706 56 45 300 1006 1027 OAI22_X1 $T=10690 37400 0 0 $X=10575 $Y=37285
X7273 64 677 299 463 423 45 300 1001 1017 OAI22_X1 $T=10880 40200 0 0 $X=10765 $Y=40085
X7274 420 A[31] 299 722 472 711 300 1013 1025 OAI22_X1 $T=12590 23400 0 0 $X=12475 $Y=23285
X7275 707 405 299 70 58 311 300 1011 1018 OAI22_X1 $T=12590 31800 0 0 $X=12475 $Y=31685
X7276 452 421 299 459 B[31] 315 300 1003 1016 OAI22_X1 $T=13350 12200 1 0 $X=13235 $Y=10685
X7277 453 421 299 467 B[31] 69 300 1007 1023 OAI22_X1 $T=13540 15000 0 0 $X=13425 $Y=14885
X7278 463 17 299 466 322 894 300 1006 1022 OAI22_X1 $T=14110 37400 1 0 $X=13995 $Y=35885
X7279 77 58 299 89 405 830 300 1002 1022 OAI22_X1 $T=14490 34600 0 0 $X=14375 $Y=34485
X7280 317 405 299 476 58 478 300 1001 1027 OAI22_X1 $T=15820 40200 1 0 $X=15705 $Y=38685
X7281 721 A[31] 299 482 472 963 300 1004 1019 OAI22_X1 $T=17720 26200 0 0 $X=17605 $Y=26085
X7282 10 843 299 101 724 72 300 1002 1022 OAI22_X1 $T=17720 34600 0 0 $X=17605 $Y=34485
X7283 113 SUM[31] 299 245 155 492 300 1012 1015 OAI22_X1 $T=21520 3800 0 0 $X=21405 $Y=3685
X7284 506 421 299 940 B[31] 125 300 1013 1029 OAI22_X1 $T=22090 23400 1 0 $X=21975 $Y=21885
X7285 510 A[31] 299 978 472 848 300 1011 1026 OAI22_X1 $T=22850 31800 1 0 $X=22735 $Y=30285
X7286 511 421 299 943 B[31] 124 300 1013 1029 OAI22_X1 $T=23040 23400 1 0 $X=22925 $Y=21885
X7287 513 SUM[31] 299 288 155 518 300 1007 1028 OAI22_X1 $T=23420 15000 1 0 $X=23305 $Y=13485
X7288 396 SUM[31] 299 193 155 905 300 1000 1020 OAI22_X1 $T=23610 9400 1 0 $X=23495 $Y=7885
X7289 730 SUM[31] 299 183 155 742 300 1000 1016 OAI22_X1 $T=23990 9400 0 0 $X=23875 $Y=9285
X7290 835 SUM[31] 299 209 155 744 300 1009 1024 OAI22_X1 $T=24370 1000 0 0 $X=24255 $Y=885
X7291 157 421 299 947 B[31] 160 300 1008 1019 OAI22_X1 $T=25700 29000 1 0 $X=25585 $Y=27485
X7292 132 SUM[31] 299 158 155 745 300 999 1020 OAI22_X1 $T=26080 6600 0 0 $X=25965 $Y=6485
X7293 135 SUM[31] 299 216 155 746 300 1010 1021 OAI22_X1 $T=26080 20600 1 0 $X=25965 $Y=19085
X7294 726 SUM[31] 299 172 155 520 300 1012 1015 OAI22_X1 $T=26270 3800 0 0 $X=26155 $Y=3685
X7295 145 SUM[31] 299 225 155 749 300 1010 1029 OAI22_X1 $T=26650 20600 0 0 $X=26535 $Y=20485
X7296 130 SUM[31] 299 185 155 956 300 1012 1024 OAI22_X1 $T=27220 3800 1 0 $X=27105 $Y=2285
X7297 856 421 299 528 B[31] 541 300 1008 1026 OAI22_X1 $T=27220 29000 0 0 $X=27105 $Y=28885
X7298 756 751 299 152 203 540 300 1006 1027 OAI22_X1 $T=27410 37400 0 0 $X=27295 $Y=37285
X7299 10 206 299 254 189 298 300 1001 1017 OAI22_X1 $T=27410 40200 0 0 $X=27295 $Y=40085
X7300 10 203 299 239 751 298 300 1006 1022 OAI22_X1 $T=27600 37400 1 0 $X=27485 $Y=35885
X7301 144 SUM[31] 299 787 155 760 300 1010 1029 OAI22_X1 $T=28740 20600 0 0 $X=28625 $Y=20485
X7302 166 SUM[31] 299 331 155 542 300 1013 1029 OAI22_X1 $T=29690 23400 1 0 $X=29575 $Y=21885
X7303 10 339 299 231 211 298 300 1001 1027 OAI22_X1 $T=31780 40200 1 0 $X=31665 $Y=38685
X7304 207 154 299 265 233 564 300 1000 1020 OAI22_X1 $T=32160 9400 1 0 $X=32045 $Y=7885
X7305 222 331 299 570 568 574 300 1007 1028 OAI22_X1 $T=33490 15000 1 0 $X=33375 $Y=13485
X7306 571 568 299 773 787 222 300 1000 1020 OAI22_X1 $T=34060 9400 1 0 $X=33945 $Y=7885
X7307 563 218 299 568 591 262 300 1010 1029 OAI22_X1 $T=34630 20600 0 0 $X=34515 $Y=20485
X7308 207 176 299 615 234 261 300 1000 1020 OAI22_X1 $T=35770 9400 1 0 $X=35655 $Y=7885
X7309 207 328 299 589 772 261 300 1000 1016 OAI22_X1 $T=36530 9400 0 0 $X=36415 $Y=9285
X7310 10 588 299 274 779 298 300 1006 1027 OAI22_X1 $T=36720 37400 0 0 $X=36605 $Y=37285
X7311 592 210 299 599 238 958 300 1013 1029 OAI22_X1 $T=38050 23400 1 0 $X=37935 $Y=21885
X7312 592 331 299 355 247 958 300 1010 1029 OAI22_X1 $T=38240 20600 0 0 $X=38125 $Y=20485
X7313 347 595 299 603 589 607 300 1000 1020 OAI22_X1 $T=39000 9400 1 0 $X=38885 $Y=7885
X7314 791 602 299 SUM[2] 210 349 300 1013 1025 OAI22_X1 $T=39190 23400 0 0 $X=39075 $Y=23285
X7315 793 595 299 953 593 607 300 999 1020 OAI22_X1 $T=39760 6600 0 0 $X=39645 $Y=6485
X7316 257 604 299 624 266 600 300 1005 1021 OAI22_X1 $T=39760 17800 0 0 $X=39645 $Y=17685
X7317 352 787 299 610 241 793 300 1007 1028 OAI22_X1 $T=40140 15000 1 0 $X=40025 $Y=13485
X7318 609 595 299 612 615 607 300 1000 1020 OAI22_X1 $T=40520 9400 1 0 $X=40405 $Y=7885
X7319 352 233 299 798 241 585 300 1000 1016 OAI22_X1 $T=40520 9400 0 0 $X=40405 $Y=9285
X7320 967 602 299 SUM[4] 787 349 300 1010 1029 OAI22_X1 $T=40900 20600 0 0 $X=40785 $Y=20485
X7321 257 619 299 807 266 873 300 1005 1023 OAI22_X1 $T=41850 17800 1 0 $X=41735 $Y=16285
X7322 621 220 299 959 268 624 300 1010 1021 OAI22_X1 $T=42040 20600 1 0 $X=41925 $Y=19085
X7323 800 627 299 293 805 806 300 1003 1016 OAI22_X1 $T=42420 12200 1 0 $X=42305 $Y=10685
X7324 622 627 299 291 246 630 300 999 1015 OAI22_X1 $T=42610 6600 1 0 $X=42495 $Y=5085
X7325 606 246 299 810 228 804 300 1012 1015 OAI22_X1 $T=42990 3800 0 0 $X=42875 $Y=3685
X7326 805 627 299 292 246 804 300 999 1020 OAI22_X1 $T=42990 6600 0 0 $X=42875 $Y=6485
X7327 811 628 299 632 879 816 300 1004 1019 OAI22_X1 $T=42990 26200 0 0 $X=42875 $Y=26085
X7328 636 602 299 SUM[5] 225 349 300 1013 1029 OAI22_X1 $T=44130 23400 1 0 $X=44015 $Y=21885
X7329 926 263 299 640 633 365 300 1011 1026 OAI22_X1 $T=44130 31800 1 0 $X=44015 $Y=30285
X7330 544 299 539 172 185 204 300 1003 1028 NAND4_X1 $T=28930 12200 0 0 $X=28815 $Y=12085
X7331 561 299 562 867 763 559 300 1010 1021 NAND4_X1 $T=32540 20600 1 0 $X=32425 $Y=19085
X7332 B[27] 299 B[28] B[29] B[30] 811 300 1004 1019 NAND4_X1 $T=42040 26200 0 0 $X=41925 $Y=26085
X7333 B[23] 299 B[24] B[25] B[26] 628 300 1004 1025 NAND4_X1 $T=42610 26200 1 0 $X=42495 $Y=24685
X7334 A[27] 299 A[28] A[29] A[30] 816 300 1013 1025 NAND4_X1 $T=44130 23400 0 0 $X=44015 $Y=23285
X7335 A[23] 299 A[24] A[25] A[26] 879 300 1008 1019 NAND4_X1 $T=44130 29000 1 0 $X=44015 $Y=27485
X7426 300 819 302 385 299 1000 1016 XOR2_X1 $T=1000 9400 0 0 $X=885 $Y=9285
X7427 300 11 821 882 299 1003 1028 XOR2_X1 $T=1000 12200 0 0 $X=885 $Y=12085
X7428 300 9 376 656 299 1005 1021 XOR2_X1 $T=1000 17800 0 0 $X=885 $Y=17685
X7429 300 378 388 829 299 1013 1029 XOR2_X1 $T=1000 23400 1 0 $X=885 $Y=21885
X7430 300 393 824 673 299 1012 1015 XOR2_X1 $T=2900 3800 0 0 $X=2785 $Y=3685
X7431 300 15 25 674 299 999 1015 XOR2_X1 $T=3850 6600 1 0 $X=3735 $Y=5085
X7432 300 27 683 660 299 1010 1021 XOR2_X1 $T=4610 20600 1 0 $X=4495 $Y=19085
X7433 300 30 680 885 299 1004 1025 XOR2_X1 $T=4990 26200 1 0 $X=4875 $Y=24685
X7434 300 306 402 708 299 1007 1028 XOR2_X1 $T=5180 15000 1 0 $X=5065 $Y=13485
X7435 300 53 430 54 299 1013 1029 XOR2_X1 $T=9930 23400 1 0 $X=9815 $Y=21885
X7436 300 434 441 439 299 1004 1025 XOR2_X1 $T=11260 26200 1 0 $X=11145 $Y=24685
X7437 300 74 475 80 299 1004 1025 XOR2_X1 $T=15060 26200 1 0 $X=14945 $Y=24685
X7438 300 86 479 464 299 1009 1024 XOR2_X1 $T=15630 1000 0 0 $X=15515 $Y=885
X7439 300 84 719 715 299 1008 1019 XOR2_X1 $T=16010 29000 1 0 $X=15895 $Y=27485
X7440 300 96 489 100 299 1008 1026 XOR2_X1 $T=18480 29000 0 0 $X=18365 $Y=28885
X7441 300 113 492 490 299 1012 1015 XOR2_X1 $T=19050 3800 0 0 $X=18935 $Y=3685
X7442 300 115 497 732 299 1002 1018 XOR2_X1 $T=19620 34600 1 0 $X=19505 $Y=33085
X7443 300 107 734 903 299 1011 1018 XOR2_X1 $T=20190 31800 0 0 $X=20075 $Y=31685
X7444 300 136 517 515 299 1004 1025 XOR2_X1 $T=23040 26200 1 0 $X=22925 $Y=24685
X7445 300 835 744 131 299 1009 1024 XOR2_X1 $T=23230 1000 0 0 $X=23115 $Y=885
X7446 300 124 511 118 299 1010 1029 XOR2_X1 $T=23800 20600 0 0 $X=23685 $Y=20485
X7447 300 112 743 119 299 1002 1022 XOR2_X1 $T=23990 34600 0 0 $X=23875 $Y=34485
X7448 300 135 746 133 299 1010 1021 XOR2_X1 $T=24940 20600 1 0 $X=24825 $Y=19085
X7449 300 160 157 534 299 1004 1019 XOR2_X1 $T=26080 26200 0 0 $X=25965 $Y=26085
X7450 300 144 760 141 299 1010 1029 XOR2_X1 $T=27600 20600 0 0 $X=27485 $Y=20485
X7451 300 166 542 753 299 1013 1029 XOR2_X1 $T=28550 23400 1 0 $X=28435 $Y=21885
X7452 300 177 557 326 299 1013 1025 XOR2_X1 $T=30830 23400 0 0 $X=30715 $Y=23285
X7453 300 188 572 192 299 1004 1025 XOR2_X1 $T=33110 26200 1 0 $X=32995 $Y=24685
X7454 300 642 927 808 299 998 1017 XOR2_X1 $T=43940 43000 1 0 $X=43825 $Y=41485
X7455 299 369 663 1 300 999 1020 XNOR2_X1 $T=1000 6600 0 0 $X=885 $Y=6485
X7456 299 658 931 2 300 1010 1029 XNOR2_X1 $T=1000 20600 0 0 $X=885 $Y=20485
X7457 299 651 384 3 300 1004 1025 XNOR2_X1 $T=1000 26200 1 0 $X=885 $Y=24685
X7458 299 301 954 303 300 1007 1023 XNOR2_X1 $T=2140 15000 0 0 $X=2025 $Y=14885
X7459 299 307 682 21 300 1009 1024 XNOR2_X1 $T=5180 1000 0 0 $X=5065 $Y=885
X7460 299 455 701 29 300 1000 1020 XNOR2_X1 $T=5750 9400 1 0 $X=5635 $Y=7885
X7461 299 693 419 44 300 1004 1025 XNOR2_X1 $T=8220 26200 1 0 $X=8105 $Y=24685
X7462 299 315 452 62 300 1000 1016 XNOR2_X1 $T=12590 9400 0 0 $X=12475 $Y=9285
X7463 299 438 446 65 300 1009 1024 XNOR2_X1 $T=12970 1000 0 0 $X=12855 $Y=885
X7464 299 504 509 114 300 999 1015 XNOR2_X1 $T=20570 6600 1 0 $X=20455 $Y=5085
X7465 299 513 518 127 300 1007 1028 XNOR2_X1 $T=22280 15000 1 0 $X=22165 $Y=13485
X7466 299 396 905 499 300 1000 1020 XNOR2_X1 $T=22470 9400 1 0 $X=22355 $Y=7885
X7467 299 730 742 128 300 1000 1016 XNOR2_X1 $T=22850 9400 0 0 $X=22735 $Y=9285
X7468 299 137 143 741 300 1003 1028 XNOR2_X1 $T=23800 12200 0 0 $X=23685 $Y=12085
X7469 299 SUM[31] 147 150 300 1007 1028 XNOR2_X1 $T=25700 15000 1 0 $X=25585 $Y=13485
X7470 299 130 956 164 300 1009 1024 XNOR2_X1 $T=27410 1000 0 0 $X=27295 $Y=885
X7471 299 608 290 274 300 1002 1022 XNOR2_X1 $T=39950 34600 0 0 $X=39835 $Y=34485
X7472 299 814 926 289 300 1002 1018 XNOR2_X1 $T=43940 34600 1 0 $X=43825 $Y=33085
X7473 299 289 365 290 300 1002 1022 XNOR2_X1 $T=43940 34600 0 0 $X=43825 $Y=34485
X7474 374 299 300 819 1000 1020 INV_X1 $T=1950 9400 1 0 $X=1835 $Y=7885
X7475 375 299 300 301 1005 1023 INV_X1 $T=1950 17800 1 0 $X=1835 $Y=16285
X7476 648 299 300 11 1003 1028 INV_X1 $T=2140 12200 0 0 $X=2025 $Y=12085
X7477 653 299 300 9 1005 1021 INV_X1 $T=2140 17800 0 0 $X=2025 $Y=17685
X7478 373 299 300 658 1013 1029 INV_X1 $T=2140 23400 1 0 $X=2025 $Y=21885
X7479 379 299 300 369 999 1015 INV_X1 $T=2330 6600 1 0 $X=2215 $Y=5085
X7480 817 299 300 393 1012 1024 INV_X1 $T=2520 3800 1 0 $X=2405 $Y=2285
X7481 657 299 300 15 1012 1015 INV_X1 $T=2520 3800 0 0 $X=2405 $Y=3685
X7482 658 299 300 654 1010 1029 INV_X1 $T=2710 20600 0 0 $X=2595 $Y=20485
X7483 825 299 300 378 1013 1025 INV_X1 $T=2710 23400 0 0 $X=2595 $Y=23285
X7484 820 299 300 651 1004 1025 INV_X1 $T=2710 26200 1 0 $X=2595 $Y=24685
X7485 659 299 300 307 1009 1024 INV_X1 $T=2900 1000 0 0 $X=2785 $Y=885
X7486 376 299 300 661 1005 1021 INV_X1 $T=2900 17800 0 0 $X=2785 $Y=17685
X7487 384 299 300 665 1004 1025 INV_X1 $T=3660 26200 1 0 $X=3545 $Y=24685
X7488 662 299 300 672 1003 1016 INV_X1 $T=4610 12200 1 0 $X=4495 $Y=10685
X7489 675 299 300 827 1003 1028 INV_X1 $T=4990 12200 0 0 $X=4875 $Y=12085
X7490 397 299 300 883 1011 1018 INV_X1 $T=4990 31800 0 0 $X=4875 $Y=31685
X7491 669 299 300 306 1005 1023 INV_X1 $T=5180 17800 1 0 $X=5065 $Y=16285
X7492 394 299 300 932 1000 1020 INV_X1 $T=5370 9400 1 0 $X=5255 $Y=7885
X7493 683 299 300 961 1005 1021 INV_X1 $T=6320 17800 0 0 $X=6205 $Y=17685
X7494 886 299 300 377 1002 1018 INV_X1 $T=6510 34600 1 0 $X=6395 $Y=33085
X7495 680 299 300 308 1013 1025 INV_X1 $T=6700 23400 0 0 $X=6585 $Y=23285
X7496 407 299 300 887 999 1015 INV_X1 $T=7080 6600 1 0 $X=6965 $Y=5085
X7497 411 299 300 39 1013 1029 INV_X1 $T=7460 23400 1 0 $X=7345 $Y=21885
X7498 383 299 300 935 1007 1023 INV_X1 $T=7650 15000 0 0 $X=7535 $Y=14885
X7499 686 299 300 695 1005 1023 INV_X1 $T=8410 17800 1 0 $X=8295 $Y=16285
X7500 693 299 300 414 1013 1025 INV_X1 $T=8410 23400 0 0 $X=8295 $Y=23285
X7501 694 299 300 399 1008 1026 INV_X1 $T=8410 29000 0 0 $X=8295 $Y=28885
X7502 52 299 300 33 1011 1018 INV_X1 $T=8600 31800 0 0 $X=8485 $Y=31685
X7503 50 299 300 891 1013 1029 INV_X1 $T=9550 23400 1 0 $X=9435 $Y=21885
X7504 A[21] 299 300 834 1005 1021 INV_X1 $T=10120 17800 0 0 $X=10005 $Y=17685
X7505 405 299 300 58 1002 1018 INV_X1 $T=10500 34600 1 0 $X=10385 $Y=33085
X7506 426 299 300 434 1004 1019 INV_X1 $T=11070 26200 0 0 $X=10955 $Y=26085
X7507 322 299 300 17 1006 1022 INV_X1 $T=11070 37400 1 0 $X=10955 $Y=35885
X7508 420 299 300 53 1013 1025 INV_X1 $T=11260 23400 0 0 $X=11145 $Y=23285
X7509 430 299 300 711 1013 1025 INV_X1 $T=12210 23400 0 0 $X=12095 $Y=23285
X7510 B[15] 299 300 457 1002 1018 INV_X1 $T=12590 34600 1 0 $X=12475 $Y=33085
X7511 979 299 300 315 1003 1016 INV_X1 $T=12970 12200 1 0 $X=12855 $Y=10685
X7512 936 299 300 710 1012 1015 INV_X1 $T=13160 3800 0 0 $X=13045 $Y=3685
X7513 713 299 300 838 999 1020 INV_X1 $T=14490 6600 0 0 $X=14375 $Y=6485
X7514 462 299 300 728 1003 1028 INV_X1 $T=14680 12200 0 0 $X=14565 $Y=12085
X7515 467 299 300 839 1005 1023 INV_X1 $T=14680 17800 1 0 $X=14565 $Y=16285
X7516 47 299 300 7 1008 1026 INV_X1 $T=15440 29000 0 0 $X=15325 $Y=28885
X7517 459 299 300 477 1000 1016 INV_X1 $T=16200 9400 0 0 $X=16085 $Y=9285
X7518 475 299 300 896 1004 1025 INV_X1 $T=17340 26200 1 0 $X=17225 $Y=24685
X7519 719 299 300 963 1004 1019 INV_X1 $T=17340 26200 0 0 $X=17225 $Y=26085
X7520 841 299 300 99 1008 1026 INV_X1 $T=17340 29000 0 0 $X=17225 $Y=28885
X7521 480 299 300 85 998 1017 INV_X1 $T=17340 43000 1 0 $X=17225 $Y=41485
X7522 B[7] 299 300 843 1002 1018 INV_X1 $T=18100 34600 1 0 $X=17985 $Y=33085
X7523 731 299 300 96 1011 1026 INV_X1 $T=18480 31800 1 0 $X=18365 $Y=30285
X7524 A[7] 299 300 724 1002 1022 INV_X1 $T=18670 34600 0 0 $X=18555 $Y=34485
X7525 723 299 300 727 1010 1029 INV_X1 $T=18860 20600 0 0 $X=18745 $Y=20485
X7526 10 299 300 72 998 1017 INV_X1 $T=18860 43000 1 0 $X=18745 $Y=41485
X7527 504 299 300 493 999 1015 INV_X1 $T=19050 6600 1 0 $X=18935 $Y=5085
X7528 396 299 300 491 1000 1020 INV_X1 $T=19430 9400 1 0 $X=19315 $Y=7885
X7529 510 299 300 107 1011 1026 INV_X1 $T=19810 31800 1 0 $X=19695 $Y=30285
X7530 513 299 300 321 1007 1028 INV_X1 $T=20570 15000 1 0 $X=20455 $Y=13485
X7531 940 299 300 942 1013 1029 INV_X1 $T=20950 23400 1 0 $X=20835 $Y=21885
X7532 516 299 300 498 1006 1027 INV_X1 $T=21140 37400 0 0 $X=21025 $Y=37285
X7533 941 299 300 124 1010 1021 INV_X1 $T=21520 20600 1 0 $X=21405 $Y=19085
X7534 734 299 300 848 1011 1026 INV_X1 $T=22470 31800 1 0 $X=22355 $Y=30285
X7535 849 299 300 125 1010 1029 INV_X1 $T=22660 20600 0 0 $X=22545 $Y=20485
X7536 943 299 300 740 1013 1025 INV_X1 $T=22850 23400 0 0 $X=22735 $Y=23285
X7537 507 299 300 850 1002 1022 INV_X1 $T=23040 34600 0 0 $X=22925 $Y=34485
X7538 514 299 300 112 1006 1022 INV_X1 $T=23420 37400 1 0 $X=23305 $Y=35885
X7539 SUM[31] 299 300 155 1010 1021 INV_X1 $T=23800 20600 1 0 $X=23685 $Y=19085
X7540 164 299 300 140 1012 1024 INV_X1 $T=24560 3800 1 0 $X=24445 $Y=2285
X7541 947 299 300 527 1008 1019 INV_X1 $T=26650 29000 1 0 $X=26535 $Y=27485
X7542 948 299 300 159 998 1014 INV_X1 $T=26650 43000 0 0 $X=26535 $Y=42885
X7543 528 299 300 529 1011 1026 INV_X1 $T=26840 31800 1 0 $X=26725 $Y=30285
X7544 A[26] 299 300 189 1001 1017 INV_X1 $T=27030 40200 0 0 $X=26915 $Y=40085
X7545 532 299 300 169 1005 1023 INV_X1 $T=27600 17800 1 0 $X=27485 $Y=16285
X7546 165 299 300 536 1005 1021 INV_X1 $T=27980 17800 0 0 $X=27865 $Y=17685
X7547 949 299 300 160 1004 1019 INV_X1 $T=27980 26200 0 0 $X=27865 $Y=26085
X7548 253 299 300 170 1009 1024 INV_X1 $T=28550 1000 0 0 $X=28435 $Y=885
X7549 759 299 300 545 1005 1023 INV_X1 $T=28740 17800 1 0 $X=28625 $Y=16285
X7550 185 299 300 858 1012 1015 INV_X1 $T=29310 3800 0 0 $X=29195 $Y=3685
X7551 158 299 300 173 999 1015 INV_X1 $T=29310 6600 1 0 $X=29195 $Y=5085
X7552 183 299 300 202 1000 1016 INV_X1 $T=29500 9400 0 0 $X=29385 $Y=9285
X7553 546 299 300 161 1002 1018 INV_X1 $T=29880 34600 1 0 $X=29765 $Y=33085
X7554 549 299 300 198 1010 1021 INV_X1 $T=30260 20600 1 0 $X=30145 $Y=19085
X7555 980 299 300 178 1008 1026 INV_X1 $T=30260 29000 0 0 $X=30145 $Y=28885
X7556 A[23] 299 300 180 1006 1022 INV_X1 $T=30260 37400 1 0 $X=30145 $Y=35885
X7557 861 299 300 541 1008 1019 INV_X1 $T=30450 29000 1 0 $X=30335 $Y=27485
X7558 186 299 300 913 1003 1016 INV_X1 $T=31210 12200 1 0 $X=31095 $Y=10685
X7559 190 299 300 328 1000 1016 INV_X1 $T=31400 9400 0 0 $X=31285 $Y=9285
X7560 A[25] 299 300 211 1001 1027 INV_X1 $T=31400 40200 1 0 $X=31285 $Y=38685
X7561 277 299 300 197 1007 1028 INV_X1 $T=31590 15000 1 0 $X=31475 $Y=13485
X7562 559 299 300 243 1013 1029 INV_X1 $T=32160 23400 1 0 $X=32045 $Y=21885
X7563 A[27] 299 300 242 998 1014 INV_X1 $T=32730 43000 0 0 $X=32615 $Y=42885
X7564 535 299 300 275 998 1014 INV_X1 $T=33110 43000 0 0 $X=32995 $Y=42885
X7565 565 299 300 770 1008 1019 INV_X1 $T=33300 29000 1 0 $X=33185 $Y=27485
X7566 566 299 300 569 998 1017 INV_X1 $T=33300 43000 1 0 $X=33185 $Y=41485
X7567 201 299 300 567 1005 1021 INV_X1 $T=33490 17800 0 0 $X=33375 $Y=17685
X7568 248 299 300 916 999 1020 INV_X1 $T=33680 6600 0 0 $X=33565 $Y=6485
X7569 568 299 300 214 1000 1020 INV_X1 $T=33680 9400 1 0 $X=33565 $Y=7885
X7570 225 299 300 234 1005 1023 INV_X1 $T=34060 17800 1 0 $X=33945 $Y=16285
X7571 238 299 300 576 1005 1021 INV_X1 $T=34820 17800 0 0 $X=34705 $Y=17685
X7572 232 299 300 235 1013 1029 INV_X1 $T=34820 23400 1 0 $X=34705 $Y=21885
X7573 756 299 300 540 1006 1027 INV_X1 $T=34820 37400 0 0 $X=34705 $Y=37285
X7574 579 299 300 775 1005 1023 INV_X1 $T=35200 17800 1 0 $X=35085 $Y=16285
X7575 A[29] 299 300 779 1006 1027 INV_X1 $T=35200 37400 0 0 $X=35085 $Y=37285
X7576 247 299 300 581 1005 1021 INV_X1 $T=36150 17800 0 0 $X=36035 $Y=17685
X7577 583 299 300 784 1004 1025 INV_X1 $T=36150 26200 1 0 $X=36035 $Y=24685
X7578 220 299 300 268 1013 1029 INV_X1 $T=36340 23400 1 0 $X=36225 $Y=21885
X7579 331 299 300 256 1007 1023 INV_X1 $T=36720 15000 0 0 $X=36605 $Y=14885
X7580 261 299 300 207 1003 1028 INV_X1 $T=37290 12200 0 0 $X=37175 $Y=12085
X7581 A[30] 299 300 351 998 1017 INV_X1 $T=38240 43000 0 180 $X=37745 $Y=41485
X7582 603 299 300 606 999 1015 INV_X1 $T=39950 6600 1 0 $X=39835 $Y=5085
X7583 241 299 300 251 1003 1028 INV_X1 $T=40140 12200 0 0 $X=40025 $Y=12085
X7584 612 299 300 630 999 1015 INV_X1 $T=40710 6600 1 0 $X=40595 $Y=5085
X7585 274 299 300 629 1002 1022 INV_X1 $T=41090 34600 0 0 $X=40975 $Y=34485
X7586 605 299 300 285 998 1014 INV_X1 $T=41090 43000 0 0 $X=40975 $Y=42885
X7587 798 299 300 622 1000 1016 INV_X1 $T=41470 9400 0 0 $X=41355 $Y=9285
X7588 613 299 300 356 1003 1028 INV_X1 $T=41850 12200 0 0 $X=41735 $Y=12085
X7589 953 299 300 804 999 1020 INV_X1 $T=42040 6600 0 0 $X=41925 $Y=6485
X7590 213 299 300 602 1013 1025 INV_X1 $T=43180 23400 0 0 $X=43065 $Y=23285
X7591 345 299 300 633 1011 1026 INV_X1 $T=43180 31800 1 0 $X=43065 $Y=30285
X7592 299 300 403 30 1004 1025 ICV_13 $T=6130 26200 1 0 $X=6015 $Y=24685
X7593 299 300 698 934 1009 1024 ICV_13 $T=8980 1000 0 0 $X=8865 $Y=885
X7594 299 300 415 832 1003 1016 ICV_13 $T=9550 12200 1 0 $X=9435 $Y=10685
X7595 299 300 B[21] 310 1010 1021 ICV_13 $T=10120 20600 1 0 $X=10005 $Y=19085
X7596 299 300 714 895 1013 1025 ICV_13 $T=15250 23400 0 0 $X=15135 $Y=23285
X7597 299 300 721 84 1008 1026 ICV_13 $T=16200 29000 0 0 $X=16085 $Y=28885
X7598 299 300 B[31] 421 1007 1023 ICV_13 $T=18860 15000 0 0 $X=18745 $Y=14885
X7599 299 300 497 904 1002 1018 ICV_13 $T=22660 34600 1 0 $X=22545 $Y=33085
X7600 299 300 743 908 1002 1022 ICV_13 $T=25130 34600 0 0 $X=25015 $Y=34485
X7601 299 300 B[25] 339 1006 1027 ICV_13 $T=33680 37400 0 0 $X=33565 $Y=37285
X7602 299 300 A[28] 240 1001 1027 ICV_13 $T=34630 40200 1 0 $X=34515 $Y=38685
X7603 299 300 210 350 1007 1023 ICV_13 $T=38620 15000 0 0 $X=38505 $Y=14885
X7604 299 300 640 801 1008 1026 ICV_13 $T=43940 29000 0 0 $X=43825 $Y=28885
X7605 14 7 299 4 5 300 47 653 1004 1019 OAI221_X1 $T=1000 26200 0 0 $X=885 $Y=26085
X7606 5 7 299 4 6 300 47 373 1008 1019 OAI221_X1 $T=1000 29000 1 0 $X=885 $Y=27485
X7607 380 47 299 4 6 300 7 820 1008 1026 OAI221_X1 $T=1000 29000 0 0 $X=885 $Y=28885
X7608 72 B[6] 299 8 10 300 A[6] 16 1006 1022 OAI221_X1 $T=1950 37400 1 0 $X=1835 $Y=35885
X7609 72 B[5] 299 8 10 300 A[5] 24 1001 1017 OAI221_X1 $T=1950 40200 0 0 $X=1835 $Y=40085
X7610 72 B[4] 299 8 10 300 A[4] 19 998 1017 OAI221_X1 $T=2140 43000 1 0 $X=2025 $Y=41485
X7611 380 7 299 4 13 300 47 825 1008 1026 OAI221_X1 $T=3470 29000 0 0 $X=3355 $Y=28885
X7612 72 B[2] 299 8 10 300 A[2] 20 998 1014 OAI221_X1 $T=3660 43000 0 0 $X=3545 $Y=42885
X7613 390 7 299 4 14 300 47 305 1004 1019 OAI221_X1 $T=4230 26200 0 0 $X=4115 $Y=26085
X7614 392 45 299 16 18 300 35 678 1006 1027 OAI221_X1 $T=4800 37400 0 0 $X=4685 $Y=37285
X7615 18 372 299 19 23 300 45 59 1001 1027 OAI221_X1 $T=4990 40200 1 0 $X=4875 $Y=38685
X7616 685 45 299 20 18 300 668 400 998 1017 OAI221_X1 $T=4990 43000 1 0 $X=4875 $Y=41485
X7617 687 45 299 24 18 300 399 401 1001 1017 OAI221_X1 $T=5180 40200 0 0 $X=5065 $Y=40085
X7618 390 47 299 4 28 300 7 404 1004 1019 OAI221_X1 $T=5370 26200 0 0 $X=5255 $Y=26085
X7619 72 B[1] 299 8 31 300 A[1] 417 998 1014 OAI221_X1 $T=5750 43000 0 0 $X=5635 $Y=42885
X7620 412 47 299 4 13 300 7 403 1008 1019 OAI221_X1 $T=6320 29000 1 0 $X=6205 $Y=27485
X7621 406 7 299 4 28 300 47 411 1004 1019 OAI221_X1 $T=6890 26200 0 0 $X=6775 $Y=26085
X7622 412 7 299 4 40 300 47 416 1008 1019 OAI221_X1 $T=7460 29000 1 0 $X=7345 $Y=27485
X7623 448 47 299 4 40 300 7 426 1008 1019 OAI221_X1 $T=9550 29000 1 0 $X=9435 $Y=27485
X7624 437 435 299 58 59 300 17 88 1001 1027 OAI221_X1 $T=12020 40200 1 0 $X=11905 $Y=38685
X7625 18 423 299 61 64 300 45 450 998 1017 OAI221_X1 $T=12400 43000 1 0 $X=12285 $Y=41485
X7626 448 7 299 4 70 300 47 460 1008 1019 OAI221_X1 $T=13160 29000 1 0 $X=13045 $Y=27485
X7627 314 47 299 4 70 300 7 469 1008 1026 OAI221_X1 $T=14300 29000 0 0 $X=14185 $Y=28885
X7628 314 7 299 4 83 300 47 721 1011 1026 OAI221_X1 $T=14680 31800 1 0 $X=14565 $Y=30285
X7629 72 B[0] 299 8 10 300 A[0] 443 998 1017 OAI221_X1 $T=15060 43000 1 0 $X=14945 $Y=41485
X7630 83 7 299 4 89 300 47 841 1011 1018 OAI221_X1 $T=15440 31800 0 0 $X=15325 $Y=31685
X7631 72 B[3] 299 8 10 300 A[3] 61 998 1014 OAI221_X1 $T=15820 43000 0 0 $X=15705 $Y=42885
X7632 840 47 299 4 89 300 7 731 1011 1018 OAI221_X1 $T=16580 31800 0 0 $X=16465 $Y=31685
X7633 10 724 299 8 72 300 843 471 1006 1022 OAI221_X1 $T=17150 37400 1 0 $X=17035 $Y=35885
X7634 476 47 299 4 104 300 7 487 1006 1022 OAI221_X1 $T=18290 37400 1 0 $X=18175 $Y=35885
X7635 840 7 299 4 104 300 47 510 1002 1018 OAI221_X1 $T=18480 34600 1 0 $X=18365 $Y=33085
X7636 842 47 299 4 105 300 7 514 1001 1027 OAI221_X1 $T=18670 40200 1 0 $X=18555 $Y=38685
X7637 476 7 299 4 105 300 47 516 1006 1027 OAI221_X1 $T=18860 37400 0 0 $X=18745 $Y=37285
X7638 A[24] 203 299 179 A[25] 300 339 184 1001 1027 OAI221_X1 $T=28740 40200 1 0 $X=28625 $Y=38685
X7639 211 B[25] 299 184 189 300 B[26] 194 1001 1017 OAI221_X1 $T=29690 40200 0 0 $X=29575 $Y=40085
X7640 A[26] 206 299 194 A[27] 300 859 863 998 1017 OAI221_X1 $T=30450 43000 1 0 $X=30335 $Y=41485
X7641 751 B[24] 299 208 211 300 B[25] 212 1006 1027 OAI221_X1 $T=32540 37400 0 0 $X=32425 $Y=37285
X7642 A[26] 206 299 212 A[25] 300 339 236 1001 1027 OAI221_X1 $T=32730 40200 1 0 $X=32615 $Y=38685
X7643 771 220 299 213 215 300 268 196 1012 1024 OAI221_X1 $T=32920 3800 1 0 $X=32805 $Y=2285
X7644 916 251 299 217 221 300 228 227 999 1015 OAI221_X1 $T=33300 6600 1 0 $X=33185 $Y=5085
X7645 771 268 299 213 223 300 220 573 1009 1024 OAI221_X1 $T=33490 1000 0 0 $X=33375 $Y=885
X7646 222 225 299 228 230 300 568 774 1000 1016 OAI221_X1 $T=33870 9400 0 0 $X=33755 $Y=9285
X7647 223 268 299 213 249 300 220 333 1009 1024 OAI221_X1 $T=36150 1000 0 0 $X=36035 $Y=885
X7648 783 220 299 213 249 300 268 769 1009 1024 OAI221_X1 $T=37290 1000 0 0 $X=37175 $Y=885
X7649 783 268 299 213 270 300 220 789 1009 1024 OAI221_X1 $T=39190 1000 0 0 $X=39075 $Y=885
X7650 287 220 299 213 270 300 268 611 1009 1024 OAI221_X1 $T=40330 1000 0 0 $X=40215 $Y=885
X7651 810 220 299 213 287 300 268 767 1009 1024 OAI221_X1 $T=42800 1000 0 0 $X=42685 $Y=885
X7652 810 268 299 213 291 300 220 334 1009 1024 OAI221_X1 $T=43940 1000 0 0 $X=43825 $Y=885
X7653 291 268 299 213 292 300 220 552 1012 1015 OAI221_X1 $T=43940 3800 0 0 $X=43825 $Y=3685
X7654 631 220 299 213 292 300 268 548 999 1020 OAI221_X1 $T=43940 6600 0 0 $X=43825 $Y=6485
X7655 631 268 299 213 293 300 220 796 1000 1016 OAI221_X1 $T=43940 9400 0 0 $X=43825 $Y=9285
X7656 293 268 299 213 294 300 220 813 1003 1028 OAI221_X1 $T=43940 12200 0 0 $X=43825 $Y=12085
X7657 294 268 299 213 295 300 220 641 1007 1028 OAI221_X1 $T=43940 15000 1 0 $X=43825 $Y=13485
X7658 807 220 299 213 295 300 268 358 1007 1023 OAI221_X1 $T=43940 15000 0 0 $X=43825 $Y=14885
X7862 367 405 299 5 58 822 300 367 58 380 405 884 1011 1026 ICV_19 $T=1000 31800 1 0 $X=885 $Y=30285
X7863 377 372 299 381 33 56 300 668 33 382 35 377 1002 1018 ICV_19 $T=1950 34600 1 0 $X=1835 $Y=33085
X7864 386 372 299 390 405 822 300 883 405 14 58 398 1011 1026 ICV_19 $T=4040 31800 1 0 $X=3925 $Y=30285
X7865 684 405 299 412 58 884 300 667 58 13 405 692 1011 1018 ICV_19 $T=6320 31800 0 0 $X=6205 $Y=31685
X7866 685 677 299 418 668 45 300 689 677 691 41 45 1001 1017 ICV_19 $T=6320 40200 0 0 $X=6205 $Y=40085
X7867 699 405 299 448 58 684 300 692 58 40 405 311 1011 1018 ICV_19 $T=8980 31800 0 0 $X=8865 $Y=31685
X7868 468 405 299 105 58 319 300 319 405 104 58 830 1006 1027 ICV_19 $T=15820 37400 0 0 $X=15705 $Y=37285
X7869 516 A[31] 299 523 472 850 300 514 A[31] 521 472 908 1002 1018 ICV_19 $T=23800 34600 1 0 $X=23685 $Y=33085
X7870 756 242 299 754 859 540 300 338 859 264 242 298 998 1014 ICV_19 $T=30830 43000 0 0 $X=30715 $Y=42885
X7871 964 228 299 771 246 221 300 868 246 223 228 252 1012 1015 ICV_19 $T=34440 3800 0 0 $X=34325 $Y=3685
X7872 207 197 299 609 581 261 300 207 869 793 576 261 1007 1028 ICV_19 $T=35770 15000 1 0 $X=35655 $Y=13485
X7873 779 B[29] 299 244 B[28] 240 300 756 240 786 785 540 1001 1017 ICV_19 $T=35960 40200 0 0 $X=35845 $Y=40085
X7874 207 913 299 585 256 261 300 207 202 593 590 261 1003 1016 ICV_19 $T=36150 12200 1 0 $X=36035 $Y=10685
X7875 756 779 299 586 588 540 300 10 785 276 240 298 1001 1027 ICV_19 $T=36150 40200 1 0 $X=36035 $Y=38685
X7876 964 246 299 249 228 794 300 252 246 783 228 966 1012 1015 ICV_19 $T=37480 3800 0 0 $X=37365 $Y=3685
X7877 600 257 299 282 210 958 300 257 873 621 331 958 1010 1021 ICV_19 $T=40140 20600 1 0 $X=40025 $Y=19085
X7878 251 331 299 618 233 241 300 604 266 295 806 800 1007 1023 ICV_19 $T=40710 15000 0 0 $X=40595 $Y=14885
X7879 355 220 299 967 268 282 300 282 220 636 268 621 1010 1029 ICV_19 $T=41850 20600 0 0 $X=41735 $Y=20485
X7880 624 220 299 635 268 807 300 635 602 SUM[7] 233 349 1005 1021 ICV_19 $T=43180 17800 0 0 $X=43065 $Y=17685
X7881 18 41 888 417 299 300 998 1017 OAI21_X1 $T=7650 43000 1 0 $X=7535 $Y=41485
X7882 689 45 696 17 299 300 1001 1017 OAI21_X1 $T=8220 40200 0 0 $X=8105 $Y=40085
X7883 422 33 49 47 299 300 1008 1026 OAI21_X1 $T=8790 29000 0 0 $X=8675 $Y=28885
X7884 53 54 57 55 299 300 1013 1029 OAI21_X1 $T=11070 23400 1 0 $X=10955 $Y=21885
X7885 705 45 437 443 299 300 998 1017 OAI21_X1 $T=11640 43000 1 0 $X=11525 $Y=41485
X7886 440 7 893 427 299 300 1011 1026 OAI21_X1 $T=12020 31800 1 0 $X=11905 $Y=30285
X7887 66 68 63 69 299 300 1003 1028 OAI21_X1 $T=13160 12200 0 0 $X=13045 $Y=12085
X7888 73 78 82 75 299 300 1010 1029 OAI21_X1 $T=14300 20600 0 0 $X=14185 $Y=20485
X7889 74 80 79 76 299 300 1004 1019 OAI21_X1 $T=14300 26200 0 0 $X=14185 $Y=26085
X7890 60 85 929 471 299 300 1006 1022 OAI21_X1 $T=15060 37400 1 0 $X=14945 $Y=35885
X7891 96 100 103 99 299 300 1008 1026 OAI21_X1 $T=17720 29000 0 0 $X=17605 $Y=28885
X7892 119 112 122 498 299 300 1006 1022 OAI21_X1 $T=20190 37400 1 0 $X=20075 $Y=35885
X7893 109 116 117 110 299 300 1005 1021 OAI21_X1 $T=20760 17800 0 0 $X=20645 $Y=17685
X7894 124 118 121 125 299 300 1010 1029 OAI21_X1 $T=20950 20600 0 0 $X=20835 $Y=20485
X7895 144 141 151 145 299 300 1013 1029 OAI21_X1 $T=25510 23400 1 0 $X=25395 $Y=21885
X7896 156 143 852 525 299 300 1005 1023 OAI21_X1 $T=25700 17800 1 0 $X=25585 $Y=16285
X7897 153 155 532 525 299 300 1007 1023 OAI21_X1 $T=26270 15000 0 0 $X=26155 $Y=14885
X7898 153 156 550 525 299 300 1005 1023 OAI21_X1 $T=26460 17800 1 0 $X=26345 $Y=16285
X7899 755 163 171 539 299 300 1003 1028 OAI21_X1 $T=27220 12200 0 0 $X=27105 $Y=12085
X7900 910 169 854 538 299 300 1005 1023 OAI21_X1 $T=27980 17800 1 0 $X=27865 $Y=16285
X7901 245 170 855 209 299 300 1012 1024 OAI21_X1 $T=28170 3800 1 0 $X=28055 $Y=2285
X7902 537 173 857 200 299 300 999 1015 OAI21_X1 $T=28550 6600 1 0 $X=28435 $Y=5085
X7903 161 178 168 541 299 300 1008 1019 OAI21_X1 $T=28740 29000 1 0 $X=28625 $Y=27485
X7904 761 176 167 190 299 300 1000 1020 OAI21_X1 $T=28930 9400 1 0 $X=28815 $Y=7885
X7905 950 182 759 544 299 300 1005 1023 OAI21_X1 $T=29120 17800 1 0 $X=29005 $Y=16285
X7906 536 155 582 550 299 300 1005 1021 OAI21_X1 $T=29120 17800 0 0 $X=29005 $Y=17685
X7907 349 183 SUM[12] 548 299 300 1000 1020 OAI21_X1 $T=29690 9400 1 0 $X=29575 $Y=7885
X7908 261 186 766 172 299 300 1003 1028 OAI21_X1 $T=29880 12200 0 0 $X=29765 $Y=12085
X7909 545 187 549 550 299 300 1005 1023 OAI21_X1 $T=29880 17800 1 0 $X=29765 $Y=16285
X7910 261 190 764 200 299 300 999 1020 OAI21_X1 $T=30070 6600 0 0 $X=29955 $Y=6485
X7911 192 188 199 558 299 300 1004 1019 OAI21_X1 $T=30260 26200 0 0 $X=30145 $Y=26085
X7912 349 172 SUM[19] 333 299 300 1009 1024 OAI21_X1 $T=30640 1000 0 0 $X=30525 $Y=885
X7913 349 190 SUM[14] 334 299 300 1012 1024 OAI21_X1 $T=30640 3800 1 0 $X=30525 $Y=2285
X7914 349 158 SUM[21] 196 299 300 1012 1015 OAI21_X1 $T=30640 3800 0 0 $X=30525 $Y=3685
X7915 917 197 553 288 299 300 1007 1028 OAI21_X1 $T=30830 15000 1 0 $X=30715 $Y=13485
X7916 349 200 SUM[22] 556 299 300 999 1015 OAI21_X1 $T=31020 6600 1 0 $X=30905 $Y=5085
X7917 349 154 SUM[15] 767 299 300 1012 1015 OAI21_X1 $T=31400 3800 0 0 $X=31285 $Y=3685
X7918 562 204 583 563 299 300 1010 1029 OAI21_X1 $T=31780 20600 0 0 $X=31665 $Y=20485
X7919 222 216 866 220 299 300 1000 1016 OAI21_X1 $T=33110 9400 0 0 $X=32995 $Y=9285
X7920 220 232 228 229 299 300 1010 1021 OAI21_X1 $T=34250 20600 1 0 $X=34135 $Y=19085
X7921 775 234 918 216 299 300 1005 1023 OAI21_X1 $T=34440 17800 1 0 $X=34325 $Y=16285
X7922 343 244 346 580 299 300 998 1017 OAI21_X1 $T=35200 43000 1 0 $X=35085 $Y=41485
X7923 778 244 782 580 299 300 998 1014 OAI21_X1 $T=35580 43000 0 0 $X=35465 $Y=42885
X7924 351 B[30] 756 782 299 300 998 1014 OAI21_X1 $T=36340 43000 0 0 $X=36225 $Y=42885
X7925 922 256 579 787 299 300 1007 1023 OAI21_X1 $T=37100 15000 0 0 $X=36985 $Y=14885
X7926 349 253 SUM[17] 789 299 300 1009 1024 OAI21_X1 $T=38430 1000 0 0 $X=38315 $Y=885
X7927 599 268 791 594 299 300 1013 1029 OAI21_X1 $T=39000 23400 1 0 $X=38885 $Y=21885
X7928 349 186 SUM[11] 796 299 300 1000 1016 OAI21_X1 $T=39760 9400 0 0 $X=39645 $Y=9285
X7929 349 245 SUM[16] 611 299 300 1012 1024 OAI21_X1 $T=40330 3800 1 0 $X=40215 $Y=2285
X7930 349 277 SUM[9] 641 299 300 1007 1028 OAI21_X1 $T=41090 15000 1 0 $X=40975 $Y=13485
X7931 349 286 SUM[8] 358 299 300 1005 1023 OAI21_X1 $T=42800 17800 1 0 $X=42685 $Y=16285
X7932 349 288 SUM[10] 813 299 300 1003 1028 OAI21_X1 $T=43180 12200 0 0 $X=43065 $Y=12085
X7942 821 421 299 675 B[31] 11 300 1003 1028 ICV_21 $T=3280 12200 0 0 $X=3165 $Y=12085
X7943 699 58 299 314 405 77 300 1002 1018 ICV_21 $T=10880 34600 1 0 $X=10765 $Y=33085
X7944 504 SUM[31] 299 154 155 509 300 999 1015 ICV_21 $T=21710 6600 1 0 $X=21595 $Y=5085
X7945 517 421 299 945 B[31] 136 300 1004 1025 ICV_21 $T=24180 26200 1 0 $X=24065 $Y=24685
X7946 756 180 299 126 560 540 300 1006 1027 ICV_21 $T=29500 37400 0 0 $X=29385 $Y=37285
X7947 352 216 299 353 241 347 300 1003 1016 ICV_21 $T=39760 12200 1 0 $X=39645 $Y=10685
X7948 966 246 299 287 228 630 300 1012 1015 ICV_21 $T=40330 3800 0 0 $X=40215 $Y=3685
X7949 619 266 299 294 806 356 300 1007 1028 ICV_21 $T=41850 15000 1 0 $X=41735 $Y=13485
X7950 959 602 299 SUM[6] 216 349 300 1010 1021 ICV_21 $T=42990 20600 1 0 $X=42875 $Y=19085
X7961 299 300 41 33 397 399 377 1002 1018 ICV_23 $T=4990 34600 1 0 $X=4875 $Y=33085
X7962 299 300 10 834 694 310 298 1010 1021 ICV_23 $T=8980 20600 1 0 $X=8865 $Y=19085
X7963 299 300 474 472 318 A[31] 75 1010 1021 ICV_23 $T=15820 20600 1 0 $X=15705 $Y=19085
X7964 299 300 469 A[31] 718 472 896 1013 1025 ICV_23 $T=16770 23400 0 0 $X=16655 $Y=23285
X7965 299 300 487 A[31] 750 472 904 1011 1018 ICV_23 $T=22470 31800 0 0 $X=22355 $Y=31685
X7966 299 300 756 211 758 339 540 1001 1017 ICV_23 $T=28550 40200 0 0 $X=28435 $Y=40085
X7967 299 300 599 220 617 268 355 1013 1029 ICV_23 $T=40710 23400 1 0 $X=40595 $Y=21885
X7968 299 300 617 602 SUM[3] 331 349 1013 1025 ICV_23 $T=42040 23400 0 0 $X=41925 $Y=23285
X7969 299 300 356 627 631 622 806 1000 1016 ICV_23 $T=42800 9400 0 0 $X=42685 $Y=9285
X8011 777 575 231 299 300 781 1006 1022 HA_X1 $T=33490 37400 1 0 $X=33375 $Y=35885
X8012 776 565 239 299 300 575 1002 1022 HA_X1 $T=34250 34600 0 0 $X=34135 $Y=34485
X8013 780 781 254 299 300 788 1002 1022 HA_X1 $T=36150 34600 0 0 $X=36035 $Y=34485
X8014 596 264 262 299 300 973 1004 1019 HA_X1 $T=37670 26200 0 0 $X=37555 $Y=26085
X8015 598 788 264 299 300 797 1002 1022 HA_X1 $T=38050 34600 0 0 $X=37935 $Y=34485
X8016 802 797 276 299 300 620 1006 1027 HA_X1 $T=40140 37400 0 0 $X=40025 $Y=37285
X8017 803 620 274 299 300 814 1006 1022 HA_X1 $T=42420 37400 1 0 $X=42305 $Y=35885
X8018 299 300 388 671 1013 1029 ICV_27 $T=4230 23400 1 0 $X=4115 $Y=21885
X8019 299 300 305 27 1005 1021 ICV_27 $T=5180 17800 0 0 $X=5065 $Y=17685
X8020 299 300 455 828 999 1020 ICV_27 $T=6130 6600 0 0 $X=6015 $Y=6485
X8021 299 300 404 38 1013 1029 ICV_27 $T=6130 23400 1 0 $X=6015 $Y=21885
X8022 299 300 933 410 999 1020 ICV_27 $T=7080 6600 0 0 $X=6965 $Y=6485
X8023 299 300 8 677 1001 1027 ICV_27 $T=7650 40200 1 0 $X=7535 $Y=38685
X8024 299 300 433 66 1007 1028 ICV_27 $T=11070 15000 1 0 $X=10955 $Y=13485
X8025 299 300 312 438 1012 1024 ICV_27 $T=11640 3800 1 0 $X=11525 $Y=2285
X8026 299 300 929 894 1006 1027 ICV_27 $T=15250 37400 0 0 $X=15135 $Y=37285
X8027 299 300 487 115 1002 1022 ICV_27 $T=20760 34600 0 0 $X=20645 $Y=34485
X8028 299 300 945 946 1004 1019 ICV_27 $T=23990 26200 0 0 $X=23875 $Y=26085
X8029 299 300 526 136 1004 1025 ICV_27 $T=26270 26200 1 0 $X=26155 $Y=24685
X8030 299 300 193 176 1000 1020 ICV_27 $T=28360 9400 1 0 $X=28245 $Y=7885
X8031 299 300 547 757 1011 1018 ICV_27 $T=28550 31800 0 0 $X=28435 $Y=31685
X8032 299 300 B[27] 859 998 1014 ICV_27 $T=30260 43000 0 0 $X=30145 $Y=42885
X8033 299 300 766 574 1003 1028 ICV_27 $T=31020 12200 0 0 $X=30905 $Y=12085
X8034 299 300 276 273 1006 1022 ICV_27 $T=39570 37400 1 0 $X=39455 $Y=35885
X8035 299 300 353 805 1003 1016 ICV_27 $T=41850 12200 1 0 $X=41735 $Y=10685
X8036 299 300 228 246 1012 1015 ICV_27 $T=42420 3800 0 0 $X=42305 $Y=3685
X8045 395 17 884 391 299 300 1002 1022 AOI21_X1 $T=4990 34600 0 0 $X=4875 $Y=34485
X8046 442 17 684 688 299 300 1006 1022 AOI21_X1 $T=6890 37400 1 0 $X=6775 $Y=35885
X8047 309 17 692 889 299 300 1002 1022 AOI21_X1 $T=8410 34600 0 0 $X=8295 $Y=34485
X8048 422 7 55 893 299 300 1008 1026 AOI21_X1 $T=11260 29000 0 0 $X=11145 $Y=28885
X8049 35 7 73 836 299 300 1008 1019 AOI21_X1 $T=12400 29000 1 0 $X=12285 $Y=27485
X8050 758 142 906 748 299 300 1001 1017 AOI21_X1 $T=24560 40200 0 0 $X=24445 $Y=40085
X8051 524 149 939 948 299 300 998 1017 AOI21_X1 $T=25320 43000 1 0 $X=25205 $Y=41485
X8052 126 152 944 853 299 300 1001 1027 AOI21_X1 $T=25890 40200 1 0 $X=25775 $Y=38685
X8053 754 159 909 535 299 300 998 1014 AOI21_X1 $T=27030 43000 0 0 $X=26915 $Y=42885
X8054 324 167 910 857 299 300 999 1020 AOI21_X1 $T=27790 6600 0 0 $X=27675 $Y=6485
X8055 852 171 232 554 299 300 1005 1021 AOI21_X1 $T=28360 17800 0 0 $X=28245 $Y=17685
X8056 855 172 537 858 299 300 1012 1015 AOI21_X1 $T=28550 3800 0 0 $X=28435 $Y=3685
X8057 553 186 761 202 299 300 1003 1016 AOI21_X1 $T=29500 12200 1 0 $X=29385 $Y=10685
X8058 207 176 230 173 299 300 999 1020 AOI21_X1 $T=30830 6600 0 0 $X=30715 $Y=6485
X8059 768 201 950 335 299 300 1005 1023 AOI21_X1 $T=31210 17800 1 0 $X=31095 $Y=16285
X8060 207 202 571 858 299 300 1000 1020 AOI21_X1 $T=31400 9400 1 0 $X=31285 $Y=7885
X8061 A[26] 206 340 566 299 300 1001 1017 AOI21_X1 $T=32350 40200 0 0 $X=32235 $Y=40085
X8062 247 210 914 567 299 300 1005 1021 AOI21_X1 $T=32730 17800 0 0 $X=32615 $Y=17685
X8063 764 214 217 866 299 300 999 1020 AOI21_X1 $T=32920 6600 0 0 $X=32805 $Y=6485
X8064 918 233 917 869 299 300 1007 1023 AOI21_X1 $T=34440 15000 0 0 $X=34325 $Y=14885
X8065 255 241 221 773 299 300 999 1020 AOI21_X1 $T=35010 6600 0 0 $X=34895 $Y=6485
X8066 952 241 972 774 299 300 1000 1020 AOI21_X1 $T=35010 9400 1 0 $X=34895 $Y=7885
X8067 868 246 215 972 299 300 999 1015 AOI21_X1 $T=35770 6600 1 0 $X=35655 $Y=5085
X8068 248 251 964 919 299 300 999 1015 AOI21_X1 $T=36530 6600 1 0 $X=36415 $Y=5085
X8069 952 251 252 920 299 300 1000 1020 AOI21_X1 $T=36720 9400 1 0 $X=36605 $Y=7885
X8070 255 251 794 921 299 300 999 1015 AOI21_X1 $T=37290 6600 1 0 $X=37175 $Y=5085
X8071 576 247 922 350 299 300 1007 1023 AOI21_X1 $T=37860 15000 0 0 $X=37745 $Y=14885
X8072 265 251 966 601 299 300 999 1015 AOI21_X1 $T=39190 6600 1 0 $X=39075 $Y=5085
X8073 243 273 614 795 299 300 1011 1026 AOI21_X1 $T=39950 31800 1 0 $X=39835 $Y=30285
X8074 786 275 924 605 299 300 998 1014 AOI21_X1 $T=40330 43000 0 0 $X=40215 $Y=42885
X8075 586 285 925 808 299 300 998 1014 AOI21_X1 $T=42230 43000 0 0 $X=42115 $Y=42885
X8076 819 300 385 1 299 1000 1016 NOR2_X1 $T=2140 9400 0 0 $X=2025 $Y=9285
X8077 378 300 829 3 299 1004 1025 NOR2_X1 $T=2140 26200 1 0 $X=2025 $Y=24685
X8078 668 300 377 391 299 1002 1022 NOR2_X1 $T=4420 34600 0 0 $X=4305 $Y=34485
X8079 393 300 673 21 299 1009 1024 NOR2_X1 $T=4610 1000 0 0 $X=4495 $Y=885
X8080 306 300 708 303 299 1007 1023 NOR2_X1 $T=5180 15000 0 0 $X=5065 $Y=14885
X8081 677 300 17 886 299 1002 1022 NOR2_X1 $T=5750 34600 0 0 $X=5635 $Y=34485
X8082 886 300 833 398 299 1002 1018 NOR2_X1 $T=6890 34600 1 0 $X=6775 $Y=33085
X8083 56 300 377 688 299 1002 1022 NOR2_X1 $T=7080 34600 0 0 $X=6965 $Y=34485
X8084 41 300 377 889 299 1002 1018 NOR2_X1 $T=7460 34600 1 0 $X=7345 $Y=33085
X8085 677 300 322 52 299 1002 1022 NOR2_X1 $T=9170 34600 0 0 $X=9055 $Y=34485
X8086 694 300 405 422 299 1008 1026 NOR2_X1 $T=9550 29000 0 0 $X=9435 $Y=28885
X8087 423 300 677 833 299 1006 1027 NOR2_X1 $T=10120 37400 0 0 $X=10005 $Y=37285
X8088 35 300 405 440 299 1011 1026 NOR2_X1 $T=11450 31800 1 0 $X=11335 $Y=30285
X8089 434 300 439 44 299 1013 1025 NOR2_X1 $T=11640 23400 0 0 $X=11525 $Y=23285
X8090 429 300 456 62 299 1000 1020 NOR2_X1 $T=13160 9400 1 0 $X=13045 $Y=7885
X8091 85 300 71 449 299 1006 1022 NOR2_X1 $T=13540 37400 1 0 $X=13425 $Y=35885
X8092 836 300 47 75 299 1008 1019 NOR2_X1 $T=14300 29000 1 0 $X=14185 $Y=27485
X8093 480 300 71 8 299 998 1017 NOR2_X1 $T=17720 43000 1 0 $X=17605 $Y=41485
X8094 738 300 900 114 299 999 1020 NOR2_X1 $T=20000 6600 0 0 $X=19885 $Y=6485
X8095 729 300 501 127 299 1007 1023 NOR2_X1 $T=20000 15000 0 0 $X=19885 $Y=14885
X8096 733 300 902 128 299 1000 1016 NOR2_X1 $T=21140 9400 0 0 $X=21025 $Y=9285
X8097 495 300 519 741 299 1003 1016 NOR2_X1 $T=23990 12200 1 0 $X=23875 $Y=10685
X8098 150 300 SUM[31] 165 299 1007 1028 NOR2_X1 $T=25130 15000 1 0 $X=25015 $Y=13485
X8099 758 300 142 748 299 1001 1017 NOR2_X1 $T=25320 40200 0 0 $X=25205 $Y=40085
X8100 524 300 149 948 299 998 1017 NOR2_X1 $T=26080 43000 1 0 $X=25965 $Y=41485
X8101 126 300 152 853 299 1001 1027 NOR2_X1 $T=26650 40200 1 0 $X=26535 $Y=38685
X8102 329 300 530 533 299 1000 1016 NOR2_X1 $T=26840 9400 0 0 $X=26725 $Y=9285
X8103 530 300 162 544 299 1003 1016 NOR2_X1 $T=27220 12200 1 0 $X=27105 $Y=10685
X8104 533 300 162 755 299 1003 1016 NOR2_X1 $T=27790 12200 1 0 $X=27675 $Y=10685
X8105 754 300 159 535 299 998 1014 NOR2_X1 $T=27790 43000 0 0 $X=27675 $Y=42885
X8106 335 300 182 562 299 1005 1023 NOR2_X1 $T=30640 17800 1 0 $X=30525 $Y=16285
X8107 913 300 202 174 299 1000 1016 NOR2_X1 $T=30830 9400 0 0 $X=30715 $Y=9285
X8108 204 300 582 561 299 1005 1021 NOR2_X1 $T=31400 17800 0 0 $X=31285 $Y=17685
X8109 197 300 578 765 299 1007 1028 NOR2_X1 $T=32160 15000 1 0 $X=32045 $Y=13485
X8110 243 300 582 563 299 1010 1029 NOR2_X1 $T=32540 20600 0 0 $X=32425 $Y=20485
X8111 234 300 772 768 299 1007 1023 NOR2_X1 $T=32730 15000 0 0 $X=32615 $Y=14885
X8112 242 300 B[27] 566 299 998 1017 NOR2_X1 $T=32730 43000 1 0 $X=32615 $Y=41485
X8113 198 300 229 218 299 1010 1029 NOR2_X1 $T=34060 20600 0 0 $X=33945 $Y=20485
X8114 256 300 590 201 299 1005 1023 NOR2_X1 $T=36720 17800 1 0 $X=36605 $Y=16285
X8115 784 300 218 591 299 1010 1029 NOR2_X1 $T=37480 20600 1 180 $X=36795 $Y=20485
X8116 589 300 595 919 299 999 1020 NOR2_X1 $T=37100 6600 0 0 $X=36985 $Y=6485
X8117 615 300 595 920 299 1000 1020 NOR2_X1 $T=37480 9400 1 0 $X=37365 $Y=7885
X8118 593 300 595 921 299 999 1015 NOR2_X1 $T=38050 6600 1 0 $X=37935 $Y=5085
X8119 585 300 595 601 299 999 1015 NOR2_X1 $T=38620 6600 1 0 $X=38505 $Y=5085
X8120 809 300 875 269 299 1008 1026 NOR2_X1 $T=39190 29000 0 0 $X=39075 $Y=28885
X8121 354 300 243 345 299 1011 1026 NOR2_X1 $T=39380 31800 1 0 $X=39265 $Y=30285
X8122 786 300 275 605 299 998 1014 NOR2_X1 $T=39760 43000 0 0 $X=39645 $Y=42885
X8123 243 300 273 795 299 1011 1018 NOR2_X1 $T=39950 31800 0 0 $X=39835 $Y=31685
X8124 586 300 285 808 299 998 1017 NOR2_X1 $T=42230 43000 1 0 $X=42115 $Y=41485
X8125 37 12 389 932 300 299 396 1000 1016 FA_X1 $T=2710 9400 0 0 $X=2595 $Y=9285
X8126 12 22 409 672 300 299 730 1003 1016 FA_X1 $T=4990 12200 1 0 $X=4875 $Y=10685
X8127 22 26 690 827 300 299 733 1003 1028 FA_X1 $T=5370 12200 0 0 $X=5255 $Y=12085
X8128 679 32 832 934 300 299 120 1012 1024 FA_X1 $T=5940 3800 1 0 $X=5825 $Y=2285
X8129 32 34 408 887 300 299 113 1012 1015 FA_X1 $T=6130 3800 0 0 $X=6015 $Y=3685
X8130 42 37 670 892 300 299 738 1000 1020 FA_X1 $T=6890 9400 1 0 $X=6775 $Y=7885
X8131 34 42 664 410 300 299 504 999 1020 FA_X1 $T=7650 6600 0 0 $X=7535 $Y=6485
X8132 26 43 51 935 300 299 513 1007 1023 FA_X1 $T=8030 15000 0 0 $X=7915 $Y=14885
X8133 43 48 436 695 300 299 729 1005 1023 FA_X1 $T=8790 17800 1 0 $X=8675 $Y=16285
X8134 90 679 702 710 300 299 835 1012 1015 FA_X1 $T=9170 3800 0 0 $X=9055 $Y=3685
X8135 48 897 969 839 300 299 110 1005 1023 FA_X1 $T=15060 17800 1 0 $X=14945 $Y=16285
X8136 94 90 722 717 300 299 726 1012 1015 FA_X1 $T=16010 3800 0 0 $X=15895 $Y=3685
X8137 97 92 486 477 300 299 132 1000 1020 FA_X1 $T=16390 9400 1 0 $X=16275 $Y=7885
X8138 981 93 844 B[31] 300 299 320 1007 1028 FA_X1 $T=16770 15000 1 0 $X=16655 $Y=13485
X8139 92 94 728 838 300 299 130 999 1020 FA_X1 $T=16960 6600 0 0 $X=16845 $Y=6485
X8140 134 95 254 939 300 299 480 998 1014 FA_X1 $T=16960 43000 0 0 $X=16845 $Y=42885
X8141 98 97 898 473 300 299 495 1000 1016 FA_X1 $T=17340 9400 0 0 $X=17225 $Y=9285
X8142 93 98 844 B[31] 300 299 137 1003 1028 FA_X1 $T=17340 12200 0 0 $X=17225 $Y=12085
X8143 897 102 718 970 300 299 109 1005 1021 FA_X1 $T=17720 17800 0 0 $X=17605 $Y=17685
X8144 102 899 482 727 300 299 135 1010 1021 FA_X1 $T=18480 20600 1 0 $X=18365 $Y=19085
X8145 95 108 231 906 300 299 322 1001 1017 FA_X1 $T=19430 40200 0 0 $X=19315 $Y=40085
X8146 899 901 488 942 300 299 145 1013 1025 FA_X1 $T=19810 23400 0 0 $X=19695 $Y=23285
X8147 901 111 508 740 300 299 144 1004 1025 FA_X1 $T=20000 26200 1 0 $X=19885 $Y=24685
X8148 108 123 239 944 300 299 405 1001 1027 FA_X1 $T=20950 40200 1 0 $X=20835 $Y=38685
X8149 123 126 565 299 300 299 47 1006 1027 FA_X1 $T=21520 37400 0 0 $X=21405 $Y=37285
X8150 111 129 978 946 300 299 166 1008 1019 FA_X1 $T=22660 29000 1 0 $X=22545 $Y=27485
X8151 271 134 264 909 300 299 71 998 1014 FA_X1 $T=23610 43000 0 0 $X=23495 $Y=42885
X8152 139 907 523 529 300 299 558 1011 1026 FA_X1 $T=23800 31800 1 0 $X=23685 $Y=30285
X8153 129 139 750 527 300 299 177 1008 1026 FA_X1 $T=24180 29000 0 0 $X=24065 $Y=28885
X8154 907 148 521 757 300 299 188 1011 1018 FA_X1 $T=25130 31800 0 0 $X=25015 $Y=31685
X8155 148 161 119 299 300 299 192 1002 1022 FA_X1 $T=26840 34600 0 0 $X=26725 $Y=34485
X8156 226 971 231 951 300 299 577 1011 1018 FA_X1 $T=32160 31800 0 0 $X=32045 $Y=31685
X8157 971 219 239 235 300 299 870 1008 1026 FA_X1 $T=33110 29000 0 0 $X=32995 $Y=28885
X8158 915 226 784 254 300 299 871 1002 1018 FA_X1 $T=33490 34600 1 0 $X=33375 $Y=33085
X8159 267 915 596 583 300 299 587 1008 1019 FA_X1 $T=35580 29000 1 0 $X=35465 $Y=27485
X8160 278 267 614 973 300 299 799 1008 1019 FA_X1 $T=38620 29000 1 0 $X=38505 $Y=27485
X8161 284 271 276 924 300 299 363 998 1017 FA_X1 $T=39190 43000 1 0 $X=39075 $Y=41485
X8162 608 278 629 795 300 299 878 1002 1018 FA_X1 $T=40900 34600 1 0 $X=40785 $Y=33085
X8163 982 283 289 927 300 299 357 1006 1027 FA_X1 $T=42040 37400 0 0 $X=41925 $Y=37285
X8164 283 284 274 925 300 299 360 1001 1027 FA_X1 $T=42040 40200 1 0 $X=41925 $Y=38685
X8177 298 B[17] 300 A[17] 817 10 299 1009 1024 AOI22_X1 $T=1000 1000 0 0 $X=885 $Y=885
X8178 298 B[16] 300 A[16] 657 10 299 1012 1015 AOI22_X1 $T=1000 3800 0 0 $X=885 $Y=3685
X8179 298 B[14] 300 A[14] 379 10 299 999 1015 AOI22_X1 $T=1000 6600 1 0 $X=885 $Y=5085
X8180 298 B[13] 300 A[13] 374 10 299 1000 1020 AOI22_X1 $T=1000 9400 1 0 $X=885 $Y=7885
X8181 298 B[12] 300 A[12] 648 10 299 1003 1016 AOI22_X1 $T=1000 12200 1 0 $X=885 $Y=10685
X8182 298 B[11] 300 A[11] 375 10 299 1005 1023 AOI22_X1 $T=1000 17800 1 0 $X=885 $Y=16285
X8183 72 A[20] 300 B[20] 372 10 299 1002 1022 AOI22_X1 $T=1000 34600 0 0 $X=885 $Y=34485
X8184 72 A[14] 300 B[14] 392 10 299 1006 1022 AOI22_X1 $T=1000 37400 1 0 $X=885 $Y=35885
X8185 72 A[16] 300 B[16] 56 10 299 1006 1027 AOI22_X1 $T=1000 37400 0 0 $X=885 $Y=37285
X8186 72 A[13] 300 B[13] 687 10 299 1001 1027 AOI22_X1 $T=1000 40200 1 0 $X=885 $Y=38685
X8187 72 A[18] 300 B[18] 668 10 299 1001 1017 AOI22_X1 $T=1000 40200 0 0 $X=885 $Y=40085
X8188 72 A[10] 300 B[10] 685 10 299 998 1014 AOI22_X1 $T=1000 43000 0 0 $X=885 $Y=42885
X8189 298 B[18] 300 A[18] 659 10 299 1009 1024 AOI22_X1 $T=1950 1000 0 0 $X=1835 $Y=885
X8190 72 A[22] 300 B[22] 35 10 299 1002 1022 AOI22_X1 $T=1950 34600 0 0 $X=1835 $Y=34485
X8191 72 A[12] 300 B[12] 23 10 299 1001 1027 AOI22_X1 $T=1950 40200 1 0 $X=1835 $Y=38685
X8192 298 B[10] 300 A[10] 669 10 299 1005 1023 AOI22_X1 $T=4230 17800 1 0 $X=4115 $Y=16285
X8193 72 A[17] 300 B[17] 41 10 299 998 1014 AOI22_X1 $T=4800 43000 0 0 $X=4685 $Y=42885
X8194 395 322 300 17 699 418 299 1006 1022 AOI22_X1 $T=7650 37400 1 0 $X=7535 $Y=35885
X8195 418 322 300 17 830 678 299 1006 1027 AOI22_X1 $T=7840 37400 0 0 $X=7725 $Y=37285
X8196 678 322 300 17 468 400 299 1001 1027 AOI22_X1 $T=8220 40200 1 0 $X=8105 $Y=38685
X8197 72 A[9] 300 B[9] 689 31 299 998 1014 AOI22_X1 $T=8600 43000 0 0 $X=8485 $Y=42885
X8198 691 17 300 322 707 309 299 1006 1022 AOI22_X1 $T=9550 37400 1 0 $X=9435 $Y=35885
X8199 72 A[19] 300 B[19] 423 31 299 998 1014 AOI22_X1 $T=9550 43000 0 0 $X=9435 $Y=42885
X8200 833 322 300 17 667 447 299 1002 1022 AOI22_X1 $T=9740 34600 0 0 $X=9625 $Y=34485
X8201 401 17 300 322 478 691 299 1001 1017 AOI22_X1 $T=9930 40200 0 0 $X=9815 $Y=40085
X8202 298 B[19] 300 A[19] 312 10 299 1009 1024 AOI22_X1 $T=10500 1000 0 0 $X=10385 $Y=885
X8203 298 B[8] 300 A[8] 433 10 299 1003 1028 AOI22_X1 $T=10500 12200 0 0 $X=10385 $Y=12085
X8204 72 A[8] 300 B[8] 705 31 299 998 1017 AOI22_X1 $T=10690 43000 1 0 $X=10575 $Y=41485
X8205 298 B[22] 300 A[22] 979 10 299 1003 1016 AOI22_X1 $T=11070 12200 1 0 $X=10955 $Y=10685
X8206 298 B[9] 300 A[9] 928 10 299 1003 1028 AOI22_X1 $T=11450 12200 0 0 $X=11335 $Y=12085
X8207 706 17 300 322 77 442 299 1006 1022 AOI22_X1 $T=11450 37400 1 0 $X=11335 $Y=35885
X8208 447 322 300 17 311 463 299 1002 1022 AOI22_X1 $T=11640 34600 0 0 $X=11525 $Y=34485
X8209 72 A[11] 300 B[11] 64 31 299 998 1014 AOI22_X1 $T=12970 43000 0 0 $X=12855 $Y=42885
X8210 59 17 300 322 319 706 299 1006 1027 AOI22_X1 $T=13160 37400 0 0 $X=13045 $Y=37285
X8211 55 472 300 A[31] 462 465 299 1013 1029 AOI22_X1 $T=13730 23400 1 0 $X=13615 $Y=21885
X8212 894 322 300 17 317 450 299 1001 1017 AOI22_X1 $T=14300 40200 0 0 $X=14185 $Y=40085
X8213 707 405 300 58 83 466 299 1011 1018 AOI22_X1 $T=14490 31800 0 0 $X=14375 $Y=31685
X8214 478 58 300 405 840 466 299 1002 1018 AOI22_X1 $T=15440 34600 1 0 $X=15325 $Y=33085
X8215 317 405 300 58 842 700 299 1001 1017 AOI22_X1 $T=16580 40200 0 0 $X=16465 $Y=40085
X8216 298 B[20] 300 A[20] 484 10 299 1009 1024 AOI22_X1 $T=18290 1000 0 0 $X=18175 $Y=885
X8217 298 B[5] 300 A[5] 941 10 299 1010 1021 AOI22_X1 $T=21900 20600 1 0 $X=21785 $Y=19085
X8218 847 SUM[31] 300 155 286 110 299 1007 1023 AOI22_X1 $T=22660 15000 0 0 $X=22545 $Y=14885
X8219 298 B[6] 300 A[6] 849 10 299 1010 1021 AOI22_X1 $T=22850 20600 1 0 $X=22735 $Y=19085
X8220 298 B[4] 300 A[4] 526 10 299 1013 1025 AOI22_X1 $T=26080 23400 0 0 $X=25965 $Y=23285
X8221 A[31] 421 300 B[31] 531 472 299 1004 1025 AOI22_X1 $T=26840 26200 1 0 $X=26725 $Y=24685
X8222 298 B[3] 300 A[3] 949 10 299 1004 1025 AOI22_X1 $T=27790 26200 1 0 $X=27675 $Y=24685
X8223 298 B[0] 300 A[0] 546 10 299 1002 1018 AOI22_X1 $T=30260 34600 1 0 $X=30145 $Y=33085
X8224 298 B[1] 300 A[1] 980 10 299 1008 1026 AOI22_X1 $T=30640 29000 0 0 $X=30525 $Y=28885
X8225 298 B[2] 300 A[2] 861 10 299 1008 1019 AOI22_X1 $T=30830 29000 1 0 $X=30715 $Y=27485
X8226 864 SUM[31] 300 155 247 558 299 1004 1025 AOI22_X1 $T=31020 26200 1 0 $X=30905 $Y=24685
X8227 557 SUM[31] 300 155 210 177 299 1013 1025 AOI22_X1 $T=31970 23400 0 0 $X=31855 $Y=23285
X8228 854 565 300 770 279 220 299 1004 1019 AOI22_X1 $T=33490 26200 0 0 $X=33375 $Y=26085
X8229 863 569 300 B[28] 778 240 299 998 1014 AOI22_X1 $T=33490 43000 0 0 $X=33375 $Y=42885
X8230 265 241 300 251 868 570 299 999 1020 AOI22_X1 $T=34060 6600 0 0 $X=33945 $Y=6485
X8231 572 SUM[31] 300 155 238 188 299 1004 1025 AOI22_X1 $T=34250 26200 1 0 $X=34135 $Y=24685
X8232 354 776 300 870 260 345 299 1011 1026 AOI22_X1 $T=35200 31800 1 0 $X=35085 $Y=30285
X8233 354 777 300 577 259 345 299 1011 1018 AOI22_X1 $T=35200 31800 0 0 $X=35085 $Y=31685
X8234 232 581 300 576 957 268 299 1010 1021 AOI22_X1 $T=35960 20600 1 0 $X=35845 $Y=19085
X8235 354 598 300 587 872 345 299 1008 1026 AOI22_X1 $T=36150 29000 0 0 $X=36035 $Y=28885
X8236 354 780 300 871 258 345 299 1002 1018 AOI22_X1 $T=36530 34600 1 0 $X=36415 $Y=33085
X8237 779 B[29] 300 B[30] 580 351 299 998 1017 AOI22_X1 $T=36910 43000 1 0 $X=36795 $Y=41485
X8238 241 581 300 234 873 251 299 1005 1023 AOI22_X1 $T=37290 17800 1 0 $X=37175 $Y=16285
X8239 241 576 300 590 600 251 299 1005 1023 AOI22_X1 $T=38240 17800 1 0 $X=38125 $Y=16285
X8240 606 246 300 228 270 794 299 1012 1015 AOI22_X1 $T=39380 3800 0 0 $X=39265 $Y=3685
X8241 241 350 300 772 604 251 299 1007 1023 AOI22_X1 $T=39760 15000 0 0 $X=39645 $Y=14885
X8242 354 802 300 799 281 345 299 1011 1026 AOI22_X1 $T=41660 31800 1 0 $X=41545 $Y=30285
X8243 354 803 300 878 280 345 299 1011 1018 AOI22_X1 $T=41660 31800 0 0 $X=41545 $Y=31685
X8244 872 258 259 260 299 300 875 1011 1026 OR4_X1 $T=37670 31800 1 0 $X=37555 $Y=30285
X8245 801 279 280 281 299 300 809 1008 1019 OR4_X1 $T=41660 29000 1 0 $X=41545 $Y=27485
X8294 381 299 300 367 382 822 1011 1018 ICV_35 $T=1760 31800 0 0 $X=1645 $Y=31685
X8295 419 299 300 890 416 693 1004 1025 ICV_35 $T=9360 26200 1 0 $X=9245 $Y=24685
X8296 928 299 300 69 454 486 1003 1028 ICV_35 $T=13920 12200 0 0 $X=13805 $Y=12085
X8297 460 299 300 76 469 74 1004 1019 ICV_35 $T=15060 26200 0 0 $X=14945 $Y=26085
X8298 481 299 300 970 318 898 1005 1023 ICV_35 $T=18100 17800 1 0 $X=17985 $Y=16285
X8299 853 299 300 142 748 149 1001 1017 ICV_35 $T=25890 40200 0 0 $X=25775 $Y=40085
X8300 A[24] 299 300 751 B[24] 203 1006 1022 ICV_35 $T=26840 37400 1 0 $X=26725 $Y=35885
X8301 288 299 300 578 286 869 1007 1028 ICV_35 $T=35010 15000 1 0 $X=34895 $Y=13485
X8302 632 299 300 597 263 354 1004 1019 ICV_35 $T=41090 26200 0 0 $X=40975 $Y=26085
X8345 299 300 301 881 1007 1023 ICV_38 $T=1000 15000 0 0 $X=885 $Y=14885
X8346 299 300 931 676 1010 1029 ICV_38 $T=3090 20600 0 0 $X=2975 $Y=20485
X8347 299 300 449 45 1006 1022 ICV_38 $T=12400 37400 1 0 $X=12285 $Y=35885
X8348 299 300 720 717 1012 1024 ICV_38 $T=16200 3800 1 0 $X=16085 $Y=2285
X8349 299 300 845 119 1001 1027 ICV_38 $T=19810 40200 1 0 $X=19695 $Y=38685
X8350 299 300 216 772 1007 1023 ICV_38 $T=33300 15000 0 0 $X=33185 $Y=14885
X8351 299 300 B[29] 588 1006 1027 ICV_38 $T=35580 37400 0 0 $X=35465 $Y=37285
X8352 299 300 B[28] 785 1001 1027 ICV_38 $T=38050 40200 1 0 $X=37935 $Y=38685
X8353 299 300 618 619 1005 1023 ICV_38 $T=40710 17800 1 0 $X=40595 $Y=16285
X8354 701 421 299 704 B[31] 455 300 704 892 1000 1016 ICV_39 $T=9550 9400 0 0 $X=9435 $Y=9285
X8355 426 A[31] 299 436 472 444 300 441 444 1004 1019 ICV_39 $T=11450 26200 0 0 $X=11335 $Y=26085
X8356 446 421 299 936 B[31] 438 300 438 712 1012 1024 ICV_39 $T=12970 3800 1 0 $X=12855 $Y=2285
X8357 10 457 299 455 837 72 300 A[15] 837 1002 1018 ICV_39 $T=12970 34600 1 0 $X=12855 $Y=33085
X8358 460 A[31] 299 969 472 895 300 A[31] 472 1013 1029 ICV_39 $T=14680 23400 1 0 $X=14565 $Y=21885
X8359 479 421 299 720 B[31] 86 300 484 86 1012 1024 ICV_39 $T=17340 3800 1 0 $X=17225 $Y=2285
X8360 841 A[31] 299 488 472 955 300 494 955 1008 1019 ICV_39 $T=19050 29000 1 0 $X=18935 $Y=27485
X8361 731 A[31] 299 508 472 737 300 489 737 1008 1026 ICV_39 $T=20760 29000 0 0 $X=20645 $Y=28885
X8362 756 189 299 524 206 540 300 B[26] 206 998 1017 ICV_39 $T=28360 43000 1 0 $X=28245 $Y=41485
X8363 10 560 299 565 180 298 300 B[23] 560 1002 1022 ICV_39 $T=29880 34600 0 0 $X=29765 $Y=34485
X8364 207 578 299 347 350 261 300 787 590 1007 1028 ICV_39 $T=37670 15000 1 0 $X=37555 $Y=13485
X8365 352 225 299 613 241 609 300 610 800 1003 1028 ICV_39 $T=40520 12200 0 0 $X=40405 $Y=12085
X8470 243 220 854 299 300 1004 1025 NOR2_X2 $T=35200 26200 1 0 $X=35085 $Y=24685
X8471 354 213 272 299 300 1004 1019 NOR2_X2 $T=39570 26200 0 0 $X=39455 $Y=26085
X8491 174 299 193 190 300 182 1003 1016 NAND3_X1 $T=28740 12200 1 0 $X=28625 $Y=10685
X8492 539 299 172 185 300 187 1007 1028 NAND3_X1 $T=28740 15000 1 0 $X=28625 $Y=13485
X8493 765 299 233 286 300 335 1007 1023 NAND3_X1 $T=30830 15000 0 0 $X=30715 $Y=14885
X8494 246 299 261 262 300 266 1003 1028 NAND3_X1 $T=38240 12200 0 0 $X=38125 $Y=12085
X8495 228 299 261 262 300 257 1005 1021 NAND3_X1 $T=38240 17800 0 0 $X=38125 $Y=17685
X8496 602 957 592 299 263 272 247 SUM[1] 300 1013 1025 OAI33_X1 $T=37860 23400 0 0 $X=37745 $Y=23285
X8497 269 531 597 299 263 272 238 SUM[0] 300 1004 1025 OAI33_X1 $T=38050 26200 1 0 $X=37935 $Y=24685
X8508 299 300 38 46 36 39 1010 1029 ICV_45 $T=6700 20600 0 0 $X=6585 $Y=20485
X8509 299 300 18 435 56 17 1001 1027 ICV_45 $T=11070 40200 1 0 $X=10955 $Y=38685
X8510 299 300 835 138 131 726 1012 1015 ICV_45 $T=23610 3800 0 0 $X=23495 $Y=3685
X8511 299 300 130 146 140 132 999 1020 ICV_45 $T=24370 6600 0 0 $X=24255 $Y=6485
X8512 299 300 147 538 165 SUM[31] 1007 1023 ICV_45 $T=27410 15000 0 0 $X=27295 $Y=14885
X8513 299 300 536 554 155 559 1010 1021 ICV_45 $T=29310 20600 1 0 $X=29195 $Y=19085
X8514 299 300 349 SUM[20] 185 573 1009 1024 ICV_45 $T=29690 1000 0 0 $X=29575 $Y=885
X8515 299 300 763 325 191 765 1007 1023 ICV_45 $T=29880 15000 0 0 $X=29765 $Y=14885
X8516 299 300 349 SUM[13] 193 552 999 1015 ICV_45 $T=30070 6600 1 0 $X=29955 $Y=5085
X8517 299 300 349 SUM[18] 209 769 1009 1024 ICV_45 $T=32540 1000 0 0 $X=32425 $Y=885
X8518 299 300 592 594 247 268 1013 1029 ICV_45 $T=37100 23400 1 0 $X=36985 $Y=21885
X8532 564 288 299 210 222 224 300 209 248 1003 1016 OAI222_X1 $T=33110 12200 1 0 $X=32995 $Y=10685
X8533 564 286 299 238 222 224 300 245 255 1003 1016 OAI222_X1 $T=34630 12200 1 0 $X=34515 $Y=10685
X8534 564 277 299 247 222 224 300 253 952 1003 1028 OAI222_X1 $T=35770 12200 0 0 $X=35655 $Y=12085
X8535 218 300 229 241 951 299 1013 1029 AOI21_X2 $T=33490 23400 1 0 $X=33375 $Y=21885
X8536 591 300 218 261 784 299 1010 1029 AOI21_X2 $T=35580 20600 0 0 $X=35465 $Y=20485
X8550 651 300 378 829 299 2 1013 1025 NOR3_X1 $T=1950 23400 0 0 $X=1835 $Y=23285
X8551 369 300 819 385 299 29 1000 1020 NOR3_X1 $T=3470 9400 1 0 $X=3355 $Y=7885
X8552 307 300 393 673 299 65 1012 1024 NOR3_X1 $T=5180 3800 1 0 $X=5065 $Y=2285
X8553 315 300 429 456 299 87 1000 1020 NOR3_X1 $T=13730 9400 1 0 $X=13615 $Y=7885
X8554 730 300 733 902 299 499 1000 1016 NOR3_X1 $T=20380 9400 0 0 $X=20265 $Y=9285
X8555 726 300 835 131 299 164 1012 1024 NOR3_X1 $T=23800 3800 1 0 $X=23685 $Y=2285
X8556 137 300 495 519 299 150 1003 1016 NOR3_X1 $T=24560 12200 1 0 $X=24445 $Y=10685
X8557 914 300 234 772 299 763 1005 1023 NOR3_X1 $T=33300 17800 1 0 $X=33185 $Y=16285
X8558 567 300 576 192 299 867 1010 1021 NOR3_X1 $T=33490 20600 1 0 $X=33375 $Y=19085
X8559 406 47 4 300 49 420 299 1008 1019 OAI211_X1 $T=8600 29000 1 0 $X=8485 $Y=27485
X8560 468 58 7 300 88 106 299 1001 1027 OAI211_X1 $T=14870 40200 1 0 $X=14755 $Y=38685
X8561 842 7 4 300 106 845 299 1001 1017 OAI211_X1 $T=18480 40200 0 0 $X=18365 $Y=40085
X8562 751 B[24] B[23] 300 180 179 299 1006 1022 OAI211_X1 $T=28550 37400 1 0 $X=28435 $Y=35885
X8563 A[24] 203 560 300 A[23] 208 299 1006 1027 OAI211_X1 $T=31590 37400 0 0 $X=31475 $Y=37285
X8564 215 220 213 300 227 556 299 1012 1015 OAI211_X1 $T=33490 3800 0 0 $X=33375 $Y=3685
X8576 54 46 299 300 50 1010 1029 AND2_X1 $T=8600 20600 0 0 $X=8485 $Y=20485
X8577 4 52 299 300 427 1011 1026 AND2_X1 $T=9930 31800 1 0 $X=9815 $Y=30285
X8578 78 57 299 300 465 1010 1029 AND2_X1 $T=12210 20600 0 0 $X=12095 $Y=20485
X8579 708 63 299 300 453 1007 1023 AND2_X1 $T=12780 15000 0 0 $X=12665 $Y=14885
X8580 439 79 299 300 714 1013 1025 AND2_X1 $T=14490 23400 0 0 $X=14375 $Y=23285
X8581 81 82 299 300 474 1010 1029 AND2_X1 $T=15060 20600 0 0 $X=14945 $Y=20485
X8582 A[31] 81 299 300 844 1007 1023 AND2_X1 $T=18100 15000 0 0 $X=17985 $Y=14885
X8583 715 103 299 300 494 1008 1019 AND2_X1 $T=18290 29000 1 0 $X=18175 $Y=27485
X8584 501 117 299 300 847 1005 1023 AND2_X1 $T=21140 17800 1 0 $X=21025 $Y=16285
X8585 503 121 299 300 506 1013 1029 AND2_X1 $T=21330 23400 1 0 $X=21215 $Y=21885
X8586 732 122 299 300 507 1002 1022 AND2_X1 $T=21330 34600 0 0 $X=21215 $Y=34485
X8587 140 138 299 300 520 1012 1015 AND2_X1 $T=24560 3800 0 0 $X=24445 $Y=3685
X8588 519 146 299 300 745 999 1020 AND2_X1 $T=25320 6600 0 0 $X=25205 $Y=6485
X8589 133 151 299 300 749 1010 1029 AND2_X1 $T=25890 20600 0 0 $X=25775 $Y=20485
X8590 200 158 299 300 539 999 1020 AND2_X1 $T=27030 6600 0 0 $X=26915 $Y=6485
X8591 534 168 299 300 856 1008 1019 AND2_X1 $T=27980 29000 1 0 $X=27865 $Y=27485
X8592 326 199 299 300 864 1004 1019 AND2_X1 $T=31020 26200 0 0 $X=30905 $Y=26085
X8593 36 38 39 299 300 54 1010 1029 OR3_X1 $T=7650 20600 0 0 $X=7535 $Y=20485
X8594 54 53 55 299 300 78 1010 1029 OR3_X1 $T=11260 20600 0 0 $X=11145 $Y=20485
X8595 68 66 69 299 300 708 1007 1028 OR3_X1 $T=13160 15000 1 0 $X=13045 $Y=13485
X8596 78 73 75 299 300 81 1010 1021 OR3_X1 $T=13920 20600 1 0 $X=13805 $Y=19085
X8597 80 74 76 299 300 439 1004 1025 OR3_X1 $T=14110 26200 1 0 $X=13995 $Y=24685
X8598 100 96 99 299 300 715 1011 1026 OR3_X1 $T=17530 31800 1 0 $X=17415 $Y=30285
X8599 116 109 110 299 300 501 1005 1023 OR3_X1 $T=20190 17800 1 0 $X=20075 $Y=16285
X8600 498 112 119 299 300 732 1006 1022 OR3_X1 $T=20950 37400 1 0 $X=20835 $Y=35885
X8601 118 124 125 299 300 503 1010 1029 OR3_X1 $T=21710 20600 0 0 $X=21595 $Y=20485
X8602 140 130 132 299 300 519 999 1015 OR3_X1 $T=23800 6600 1 0 $X=23685 $Y=5085
X8603 141 144 145 299 300 133 1010 1029 OR3_X1 $T=24940 20600 0 0 $X=24825 $Y=20485
X8604 541 178 161 299 300 534 1008 1019 OR3_X1 $T=29500 29000 1 0 $X=29385 $Y=27485
X8605 558 188 192 299 300 326 1004 1025 OR3_X1 $T=30070 26200 1 0 $X=29955 $Y=24685
X8606 320 SUM[31] 299 300 1007 1028 CLKBUF_X2 $T=19810 15000 1 0 $X=19695 $Y=13485
X8607 72 298 299 300 1006 1022 CLKBUF_X2 $T=29500 37400 1 0 $X=29385 $Y=35885
X8608 413 472 299 415 A[31] 38 300 38 413 36 1010 1021 ICV_48 $T=6510 20600 1 0 $X=6395 $Y=19085
X8609 445 472 299 454 A[31] 73 300 73 445 78 1010 1021 ICV_48 $T=11830 20600 1 0 $X=11715 $Y=19085
X8610 709 421 299 713 B[31] 429 300 429 709 456 999 1020 ICV_48 $T=12020 6600 0 0 $X=11905 $Y=6485
X8611 716 421 299 481 B[31] 66 300 66 716 68 1007 1023 ICV_48 $T=16010 15000 0 0 $X=15895 $Y=14885
X8612 880 421 299 723 B[31] 101 300 101 880 503 1013 1029 ICV_48 $T=16770 23400 1 0 $X=16655 $Y=21885
X8613 733 SUM[31] 299 186 155 502 300 733 502 902 1003 1028 ICV_48 $T=20380 12200 0 0 $X=20265 $Y=12085
X8614 738 SUM[31] 299 190 155 735 300 738 735 900 999 1020 ICV_48 $T=20570 6600 0 0 $X=20455 $Y=6485
X8615 729 SUM[31] 299 277 155 736 300 729 736 501 1007 1023 ICV_48 $T=20570 15000 0 0 $X=20455 $Y=14885
X8616 120 SUM[31] 299 253 155 505 300 120 505 500 1009 1024 ICV_48 $T=21140 1000 0 0 $X=21025 $Y=885
X8617 109 SUM[31] 299 233 155 512 300 109 512 116 1005 1021 ICV_48 $T=22470 17800 0 0 $X=22355 $Y=17685
X8618 495 SUM[31] 299 200 155 522 300 495 522 519 1000 1020 ICV_48 $T=24560 9400 1 0 $X=24445 $Y=7885
X8619 543 421 299 547 B[31] 178 300 178 543 161 1011 1026 ICV_48 $T=28550 31800 1 0 $X=28435 $Y=30285
X8630 372 58 300 33 35 299 405 406 1008 1026 AOI221_X1 $T=6130 29000 0 0 $X=6015 $Y=28885
X8631 10 457 300 71 72 299 837 60 1002 1022 AOI221_X1 $T=13350 34600 0 0 $X=13235 $Y=34485
.ENDS
***************************************
