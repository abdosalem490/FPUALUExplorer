/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 16 23:17:26 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2842027065 */

module datapath(B, p_0);
   input [31:0]B;
   output [31:0]p_0;

   XOR2_X1 i_0 (.A(B[1]), .B(B[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(B[2]), .B1(B[1]), .B2(B[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(B[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(B[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(B[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(B[6]), .B1(n_27), .B2(B[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(B[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(B[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(B[9]), .B1(n_25), .B2(B[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(B[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(B[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(B[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(B[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(B[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(B[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(B[16]), .B1(n_19), .B2(B[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(B[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(B[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(B[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(B[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(B[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(B[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(B[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(B[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(B[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(B[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(B[27]), .B1(n_9), .B2(B[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(B[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(B[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(B[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(B[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(B[28]), .A3(B[29]), .A4(B[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(B[28]), .A3(B[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(B[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(B[26]), .A3(B[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(B[23]), .A3(B[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(B[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(B[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(B[18]), .A3(B[19]), .A4(B[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(B[18]), .A3(B[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(B[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(B[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(B[15]), .A3(B[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(B[12]), .A3(B[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(B[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(B[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(B[8]), .A3(B[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(B[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(B[5]), .A3(B[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(B[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(B[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(B[2]), .A2(B[1]), .A3(B[0]), .ZN(n_29));
   INV_X1 i_61 (.A(B[11]), .ZN(n_30));
   INV_X1 i_62 (.A(B[14]), .ZN(n_31));
   INV_X1 i_63 (.A(B[21]), .ZN(n_32));
   INV_X1 i_64 (.A(B[25]), .ZN(n_33));
endmodule

module datapath__0_0(A, p_0);
   input [31:0]A;
   output [31:0]p_0;

   XOR2_X1 i_0 (.A(A[1]), .B(A[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(A[2]), .B1(A[1]), .B2(A[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(A[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(A[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(A[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(A[6]), .B1(n_27), .B2(A[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(A[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(A[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(A[9]), .B1(n_25), .B2(A[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(A[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(A[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(A[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(A[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(A[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(A[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(A[16]), .B1(n_19), .B2(A[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(A[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(A[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(A[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(A[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(A[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(A[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(A[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(A[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(A[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(A[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(A[27]), .B1(n_9), .B2(A[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(A[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(A[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(A[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(A[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(A[28]), .A3(A[29]), .A4(A[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(A[28]), .A3(A[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(A[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(A[26]), .A3(A[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(A[23]), .A3(A[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(A[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(A[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(A[18]), .A3(A[19]), .A4(A[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(A[18]), .A3(A[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(A[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(A[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(A[15]), .A3(A[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(A[12]), .A3(A[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(A[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(A[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(A[8]), .A3(A[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(A[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(A[5]), .A3(A[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(A[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(A[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(A[2]), .A2(A[1]), .A3(A[0]), .ZN(n_29));
   INV_X1 i_61 (.A(A[11]), .ZN(n_30));
   INV_X1 i_62 (.A(A[14]), .ZN(n_31));
   INV_X1 i_63 (.A(A[21]), .ZN(n_32));
   INV_X1 i_64 (.A(A[25]), .ZN(n_33));
endmodule

module datapath__0_17(p_0, p_1);
   input [63:0]p_0;
   output [63:0]p_1;

   XOR2_X1 i_0 (.A(p_0[1]), .B(p_0[0]), .Z(p_1[1]));
   AND2_X1 i_1 (.A1(n_60), .A2(n_0), .ZN(p_1[2]));
   OAI21_X1 i_2 (.A(p_0[2]), .B1(p_0[1]), .B2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_0[3]), .B(n_60), .Z(p_1[3]));
   XOR2_X1 i_4 (.A(p_0[4]), .B(n_59), .Z(p_1[4]));
   XOR2_X1 i_5 (.A(p_0[5]), .B(n_58), .Z(p_1[5]));
   AND2_X1 i_6 (.A1(n_57), .A2(n_1), .ZN(p_1[6]));
   OAI21_X1 i_7 (.A(p_0[6]), .B1(n_58), .B2(p_0[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_0[7]), .B(n_57), .Z(p_1[7]));
   XOR2_X1 i_9 (.A(p_0[8]), .B(n_56), .Z(p_1[8]));
   AND2_X1 i_10 (.A1(n_55), .A2(n_2), .ZN(p_1[9]));
   OAI21_X1 i_11 (.A(p_0[9]), .B1(n_56), .B2(p_0[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_0[10]), .B(n_55), .Z(p_1[10]));
   XNOR2_X1 i_13 (.A(p_0[11]), .B(n_54), .ZN(p_1[11]));
   XOR2_X1 i_14 (.A(p_0[12]), .B(n_53), .Z(p_1[12]));
   XNOR2_X1 i_15 (.A(p_0[13]), .B(n_52), .ZN(p_1[13]));
   XOR2_X1 i_16 (.A(p_0[14]), .B(n_51), .Z(p_1[14]));
   AND2_X1 i_17 (.A1(n_50), .A2(n_3), .ZN(p_1[15]));
   OAI21_X1 i_18 (.A(p_0[15]), .B1(n_51), .B2(p_0[14]), .ZN(n_3));
   XOR2_X1 i_19 (.A(p_0[16]), .B(n_50), .Z(p_1[16]));
   XOR2_X1 i_20 (.A(p_0[17]), .B(n_49), .Z(p_1[17]));
   XOR2_X1 i_21 (.A(p_0[18]), .B(n_48), .Z(p_1[18]));
   XNOR2_X1 i_22 (.A(p_0[19]), .B(n_47), .ZN(p_1[19]));
   XNOR2_X1 i_23 (.A(p_0[20]), .B(n_46), .ZN(p_1[20]));
   XNOR2_X1 i_24 (.A(p_0[21]), .B(n_45), .ZN(p_1[21]));
   XOR2_X1 i_25 (.A(p_0[22]), .B(n_44), .Z(p_1[22]));
   XOR2_X1 i_26 (.A(p_0[23]), .B(n_43), .Z(p_1[23]));
   XNOR2_X1 i_27 (.A(p_0[24]), .B(n_42), .ZN(p_1[24]));
   XNOR2_X1 i_28 (.A(p_0[25]), .B(n_41), .ZN(p_1[25]));
   XNOR2_X1 i_29 (.A(p_0[26]), .B(n_40), .ZN(p_1[26]));
   XOR2_X1 i_30 (.A(p_0[27]), .B(n_39), .Z(p_1[27]));
   XOR2_X1 i_31 (.A(p_0[28]), .B(n_38), .Z(p_1[28]));
   XNOR2_X1 i_32 (.A(p_0[29]), .B(n_37), .ZN(p_1[29]));
   XNOR2_X1 i_33 (.A(p_0[30]), .B(n_36), .ZN(p_1[30]));
   XNOR2_X1 i_34 (.A(p_0[31]), .B(n_35), .ZN(p_1[31]));
   XOR2_X1 i_35 (.A(p_0[32]), .B(n_34), .Z(p_1[32]));
   XOR2_X1 i_36 (.A(p_0[33]), .B(n_33), .Z(p_1[33]));
   XNOR2_X1 i_37 (.A(p_0[34]), .B(n_32), .ZN(p_1[34]));
   XNOR2_X1 i_38 (.A(p_0[35]), .B(n_31), .ZN(p_1[35]));
   XNOR2_X1 i_39 (.A(p_0[36]), .B(n_30), .ZN(p_1[36]));
   XOR2_X1 i_40 (.A(p_0[37]), .B(n_29), .Z(p_1[37]));
   XOR2_X1 i_41 (.A(p_0[38]), .B(n_28), .Z(p_1[38]));
   XNOR2_X1 i_42 (.A(p_0[39]), .B(n_27), .ZN(p_1[39]));
   XNOR2_X1 i_43 (.A(p_0[40]), .B(n_26), .ZN(p_1[40]));
   XOR2_X1 i_44 (.A(p_0[41]), .B(n_25), .Z(p_1[41]));
   XNOR2_X1 i_45 (.A(p_0[42]), .B(n_24), .ZN(p_1[42]));
   XOR2_X1 i_46 (.A(p_0[43]), .B(n_23), .Z(p_1[43]));
   AND2_X1 i_47 (.A1(n_22), .A2(n_4), .ZN(p_1[44]));
   OAI21_X1 i_48 (.A(p_0[44]), .B1(n_23), .B2(p_0[43]), .ZN(n_4));
   XOR2_X1 i_49 (.A(p_0[45]), .B(n_22), .Z(p_1[45]));
   XOR2_X1 i_50 (.A(p_0[46]), .B(n_21), .Z(p_1[46]));
   XOR2_X1 i_51 (.A(p_0[47]), .B(n_20), .Z(p_1[47]));
   XOR2_X1 i_52 (.A(p_0[48]), .B(n_19), .Z(p_1[48]));
   XNOR2_X1 i_53 (.A(p_0[49]), .B(n_18), .ZN(p_1[49]));
   XNOR2_X1 i_54 (.A(p_0[50]), .B(n_17), .ZN(p_1[50]));
   XNOR2_X1 i_55 (.A(p_0[51]), .B(n_16), .ZN(p_1[51]));
   XOR2_X1 i_56 (.A(p_0[52]), .B(n_15), .Z(p_1[52]));
   XNOR2_X1 i_57 (.A(p_0[53]), .B(n_14), .ZN(p_1[53]));
   XNOR2_X1 i_58 (.A(p_0[54]), .B(n_13), .ZN(p_1[54]));
   XNOR2_X1 i_59 (.A(p_0[55]), .B(n_12), .ZN(p_1[55]));
   XOR2_X1 i_60 (.A(p_0[56]), .B(n_11), .Z(p_1[56]));
   AND2_X1 i_61 (.A1(n_10), .A2(n_5), .ZN(p_1[57]));
   OAI21_X1 i_62 (.A(p_0[57]), .B1(n_11), .B2(p_0[56]), .ZN(n_5));
   XOR2_X1 i_63 (.A(p_0[58]), .B(n_10), .Z(p_1[58]));
   XNOR2_X1 i_64 (.A(p_0[59]), .B(n_9), .ZN(p_1[59]));
   XNOR2_X1 i_65 (.A(p_0[60]), .B(n_8), .ZN(p_1[60]));
   XOR2_X1 i_66 (.A(p_0[61]), .B(n_7), .Z(p_1[61]));
   XNOR2_X1 i_67 (.A(p_0[63]), .B(n_6), .ZN(p_1[62]));
   NOR2_X1 i_68 (.A1(p_0[63]), .A2(n_6), .ZN(p_1[63]));
   NOR2_X1 i_69 (.A1(n_7), .A2(p_0[61]), .ZN(n_6));
   NAND2_X1 i_70 (.A1(n_8), .A2(n_71), .ZN(n_7));
   NOR3_X1 i_71 (.A1(n_10), .A2(p_0[58]), .A3(p_0[59]), .ZN(n_8));
   NOR2_X1 i_72 (.A1(n_10), .A2(p_0[58]), .ZN(n_9));
   OR3_X1 i_73 (.A1(n_11), .A2(p_0[56]), .A3(p_0[57]), .ZN(n_10));
   NAND2_X1 i_74 (.A1(n_12), .A2(n_70), .ZN(n_11));
   NOR4_X1 i_75 (.A1(n_15), .A2(p_0[52]), .A3(p_0[53]), .A4(p_0[54]), .ZN(n_12));
   NOR3_X1 i_76 (.A1(n_15), .A2(p_0[52]), .A3(p_0[53]), .ZN(n_13));
   NOR2_X1 i_77 (.A1(n_15), .A2(p_0[52]), .ZN(n_14));
   NAND2_X1 i_78 (.A1(n_16), .A2(n_69), .ZN(n_15));
   NOR4_X1 i_79 (.A1(n_19), .A2(p_0[48]), .A3(p_0[49]), .A4(p_0[50]), .ZN(n_16));
   NOR3_X1 i_80 (.A1(n_19), .A2(p_0[48]), .A3(p_0[49]), .ZN(n_17));
   NOR2_X1 i_81 (.A1(n_19), .A2(p_0[48]), .ZN(n_18));
   OR2_X1 i_82 (.A1(n_20), .A2(p_0[47]), .ZN(n_19));
   OR2_X1 i_83 (.A1(n_21), .A2(p_0[46]), .ZN(n_20));
   OR2_X1 i_84 (.A1(n_22), .A2(p_0[45]), .ZN(n_21));
   OR3_X1 i_85 (.A1(n_23), .A2(p_0[43]), .A3(p_0[44]), .ZN(n_22));
   NAND2_X1 i_86 (.A1(n_24), .A2(n_68), .ZN(n_23));
   NOR2_X1 i_87 (.A1(n_25), .A2(p_0[41]), .ZN(n_24));
   NAND2_X1 i_88 (.A1(n_26), .A2(n_67), .ZN(n_25));
   NOR3_X1 i_89 (.A1(n_28), .A2(p_0[38]), .A3(p_0[39]), .ZN(n_26));
   NOR2_X1 i_90 (.A1(n_28), .A2(p_0[38]), .ZN(n_27));
   OR2_X1 i_91 (.A1(n_29), .A2(p_0[37]), .ZN(n_28));
   NAND2_X1 i_92 (.A1(n_30), .A2(n_66), .ZN(n_29));
   NOR4_X1 i_93 (.A1(n_33), .A2(p_0[33]), .A3(p_0[34]), .A4(p_0[35]), .ZN(n_30));
   NOR3_X1 i_94 (.A1(n_33), .A2(p_0[33]), .A3(p_0[34]), .ZN(n_31));
   NOR2_X1 i_95 (.A1(n_33), .A2(p_0[33]), .ZN(n_32));
   OR2_X1 i_96 (.A1(n_34), .A2(p_0[32]), .ZN(n_33));
   NAND2_X1 i_97 (.A1(n_35), .A2(n_65), .ZN(n_34));
   NOR4_X1 i_98 (.A1(n_38), .A2(p_0[28]), .A3(p_0[29]), .A4(p_0[30]), .ZN(n_35));
   NOR3_X1 i_99 (.A1(n_38), .A2(p_0[28]), .A3(p_0[29]), .ZN(n_36));
   NOR2_X1 i_100 (.A1(n_38), .A2(p_0[28]), .ZN(n_37));
   OR2_X1 i_101 (.A1(n_39), .A2(p_0[27]), .ZN(n_38));
   NAND2_X1 i_102 (.A1(n_40), .A2(n_64), .ZN(n_39));
   NOR4_X1 i_103 (.A1(n_43), .A2(p_0[23]), .A3(p_0[24]), .A4(p_0[25]), .ZN(n_40));
   NOR3_X1 i_104 (.A1(n_43), .A2(p_0[23]), .A3(p_0[24]), .ZN(n_41));
   NOR2_X1 i_105 (.A1(n_43), .A2(p_0[23]), .ZN(n_42));
   OR2_X1 i_106 (.A1(n_44), .A2(p_0[22]), .ZN(n_43));
   NAND2_X1 i_107 (.A1(n_45), .A2(n_63), .ZN(n_44));
   NOR4_X1 i_108 (.A1(n_48), .A2(p_0[18]), .A3(p_0[19]), .A4(p_0[20]), .ZN(n_45));
   NOR3_X1 i_109 (.A1(n_48), .A2(p_0[18]), .A3(p_0[19]), .ZN(n_46));
   NOR2_X1 i_110 (.A1(n_48), .A2(p_0[18]), .ZN(n_47));
   OR2_X1 i_111 (.A1(n_49), .A2(p_0[17]), .ZN(n_48));
   OR2_X1 i_112 (.A1(n_50), .A2(p_0[16]), .ZN(n_49));
   OR3_X1 i_113 (.A1(n_51), .A2(p_0[14]), .A3(p_0[15]), .ZN(n_50));
   NAND2_X1 i_114 (.A1(n_52), .A2(n_62), .ZN(n_51));
   NOR2_X1 i_115 (.A1(n_53), .A2(p_0[12]), .ZN(n_52));
   NAND2_X1 i_116 (.A1(n_54), .A2(n_61), .ZN(n_53));
   NOR2_X1 i_117 (.A1(n_55), .A2(p_0[10]), .ZN(n_54));
   OR3_X1 i_118 (.A1(n_56), .A2(p_0[8]), .A3(p_0[9]), .ZN(n_55));
   OR2_X1 i_119 (.A1(n_57), .A2(p_0[7]), .ZN(n_56));
   OR3_X1 i_120 (.A1(n_58), .A2(p_0[5]), .A3(p_0[6]), .ZN(n_57));
   OR2_X1 i_121 (.A1(n_59), .A2(p_0[4]), .ZN(n_58));
   OR2_X1 i_122 (.A1(n_60), .A2(p_0[3]), .ZN(n_59));
   OR3_X1 i_123 (.A1(p_0[2]), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_60));
   INV_X1 i_124 (.A(p_0[11]), .ZN(n_61));
   INV_X1 i_125 (.A(p_0[13]), .ZN(n_62));
   INV_X1 i_126 (.A(p_0[21]), .ZN(n_63));
   INV_X1 i_127 (.A(p_0[26]), .ZN(n_64));
   INV_X1 i_128 (.A(p_0[31]), .ZN(n_65));
   INV_X1 i_129 (.A(p_0[36]), .ZN(n_66));
   INV_X1 i_130 (.A(p_0[40]), .ZN(n_67));
   INV_X1 i_131 (.A(p_0[42]), .ZN(n_68));
   INV_X1 i_132 (.A(p_0[51]), .ZN(n_69));
   INV_X1 i_133 (.A(p_0[55]), .ZN(n_70));
   INV_X1 i_134 (.A(p_0[60]), .ZN(n_71));
endmodule

module datapath__0_4(multiplier_M, accumulator_A, p_0);
   input [31:0]multiplier_M;
   input [31:0]accumulator_A;
   output [31:0]p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0[0]));
   OAI21_X1 i_1 (.A(n_154), .B1(multiplier_M[0]), .B2(accumulator_A[0]), 
      .ZN(n_0));
   XOR2_X1 i_2 (.A(n_154), .B(n_1), .Z(p_0[1]));
   OAI21_X1 i_3 (.A(n_153), .B1(multiplier_M[1]), .B2(accumulator_A[1]), 
      .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_152), .B(n_2), .ZN(p_0[2]));
   OAI21_X1 i_5 (.A(n_157), .B1(multiplier_M[2]), .B2(accumulator_A[2]), 
      .ZN(n_2));
   XOR2_X1 i_6 (.A(n_151), .B(n_3), .Z(p_0[3]));
   OAI21_X1 i_7 (.A(n_158), .B1(n_164), .B2(n_161), .ZN(n_3));
   XOR2_X1 i_8 (.A(n_149), .B(n_10), .Z(p_0[4]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_0[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_0[6]));
   NOR2_X1 i_11 (.A1(n_146), .A2(n_137), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_0[7]));
   OAI22_X1 i_13 (.A1(multiplier_M[6]), .A2(accumulator_A[6]), .B1(n_137), 
      .B2(n_7), .ZN(n_5));
   AOI21_X1 i_14 (.A(n_147), .B1(multiplier_M[5]), .B2(accumulator_A[5]), 
      .ZN(n_6));
   AOI21_X1 i_15 (.A(n_147), .B1(n_141), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_144), .B1(n_149), .B2(n_142), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_142), .B1(multiplier_M[4]), .B2(accumulator_A[4]), 
      .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_148), .A2(n_139), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_135), .B(n_18), .ZN(p_0[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_0[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_0[10]));
   NOR2_X1 i_23 (.A1(n_132), .A2(n_123), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_0[11]));
   OAI22_X1 i_25 (.A1(multiplier_M[10]), .A2(accumulator_A[10]), .B1(n_123), 
      .B2(n_15), .ZN(n_13));
   AOI21_X1 i_26 (.A(n_133), .B1(multiplier_M[9]), .B2(accumulator_A[9]), 
      .ZN(n_14));
   AOI21_X1 i_27 (.A(n_133), .B1(n_127), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_130), .B1(n_135), .B2(n_128), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_130), .B1(multiplier_M[8]), .B2(accumulator_A[8]), 
      .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_134), .A2(n_125), .ZN(n_19));
   XOR2_X1 i_32 (.A(n_121), .B(n_26), .Z(p_0[12]));
   XOR2_X1 i_33 (.A(n_25), .B(n_22), .Z(p_0[13]));
   XOR2_X1 i_34 (.A(n_23), .B(n_20), .Z(p_0[14]));
   NOR2_X1 i_35 (.A1(n_118), .A2(n_109), .ZN(n_20));
   XNOR2_X1 i_36 (.A(n_27), .B(n_21), .ZN(p_0[15]));
   OAI22_X1 i_37 (.A1(multiplier_M[14]), .A2(accumulator_A[14]), .B1(n_109), 
      .B2(n_23), .ZN(n_21));
   AOI21_X1 i_38 (.A(n_119), .B1(multiplier_M[13]), .B2(accumulator_A[13]), 
      .ZN(n_22));
   AOI21_X1 i_39 (.A(n_119), .B1(n_113), .B2(n_24), .ZN(n_23));
   INV_X1 i_40 (.A(n_25), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_116), .B1(n_121), .B2(n_114), .ZN(n_25));
   OAI21_X1 i_42 (.A(n_114), .B1(multiplier_M[12]), .B2(accumulator_A[12]), 
      .ZN(n_26));
   NOR2_X1 i_43 (.A1(n_120), .A2(n_111), .ZN(n_27));
   XOR2_X1 i_44 (.A(n_107), .B(n_34), .Z(p_0[16]));
   XOR2_X1 i_45 (.A(n_33), .B(n_30), .Z(p_0[17]));
   XOR2_X1 i_46 (.A(n_31), .B(n_28), .Z(p_0[18]));
   NOR2_X1 i_47 (.A1(n_104), .A2(n_95), .ZN(n_28));
   XNOR2_X1 i_48 (.A(n_35), .B(n_29), .ZN(p_0[19]));
   OAI22_X1 i_49 (.A1(multiplier_M[18]), .A2(accumulator_A[18]), .B1(n_95), 
      .B2(n_31), .ZN(n_29));
   AOI21_X1 i_50 (.A(n_105), .B1(multiplier_M[17]), .B2(accumulator_A[17]), 
      .ZN(n_30));
   AOI21_X1 i_51 (.A(n_105), .B1(n_99), .B2(n_32), .ZN(n_31));
   INV_X1 i_52 (.A(n_33), .ZN(n_32));
   AOI21_X1 i_53 (.A(n_102), .B1(n_107), .B2(n_100), .ZN(n_33));
   OAI21_X1 i_54 (.A(n_100), .B1(multiplier_M[16]), .B2(accumulator_A[16]), 
      .ZN(n_34));
   NOR2_X1 i_55 (.A1(n_106), .A2(n_97), .ZN(n_35));
   XOR2_X1 i_56 (.A(n_93), .B(n_42), .Z(p_0[20]));
   XOR2_X1 i_57 (.A(n_41), .B(n_38), .Z(p_0[21]));
   XOR2_X1 i_58 (.A(n_39), .B(n_36), .Z(p_0[22]));
   NOR2_X1 i_59 (.A1(n_82), .A2(n_72), .ZN(n_36));
   XNOR2_X1 i_60 (.A(n_43), .B(n_37), .ZN(p_0[23]));
   OAI21_X1 i_61 (.A(n_81), .B1(n_72), .B2(n_39), .ZN(n_37));
   NOR2_X1 i_62 (.A1(n_84), .A2(n_74), .ZN(n_38));
   INV_X1 i_63 (.A(n_40), .ZN(n_39));
   OAI21_X1 i_64 (.A(n_83), .B1(n_74), .B2(n_41), .ZN(n_40));
   AOI21_X1 i_65 (.A(n_79), .B1(n_93), .B2(n_76), .ZN(n_41));
   OAI21_X1 i_66 (.A(n_76), .B1(multiplier_M[20]), .B2(accumulator_A[20]), 
      .ZN(n_42));
   AOI21_X1 i_67 (.A(n_86), .B1(multiplier_M[23]), .B2(accumulator_A[23]), 
      .ZN(n_43));
   XOR2_X1 i_68 (.A(n_51), .B(n_50), .Z(p_0[24]));
   XOR2_X1 i_69 (.A(n_49), .B(n_47), .Z(p_0[25]));
   XNOR2_X1 i_70 (.A(n_45), .B(n_44), .ZN(p_0[26]));
   NOR2_X1 i_71 (.A1(n_91), .A2(n_48), .ZN(n_44));
   OAI21_X1 i_72 (.A(n_66), .B1(multiplier_M[26]), .B2(accumulator_A[26]), 
      .ZN(n_45));
   XNOR2_X1 i_73 (.A(n_53), .B(n_46), .ZN(p_0[27]));
   OAI21_X1 i_74 (.A(n_66), .B1(n_90), .B2(n_48), .ZN(n_46));
   AOI21_X1 i_75 (.A(n_91), .B1(multiplier_M[25]), .B2(accumulator_A[25]), 
      .ZN(n_47));
   AOI21_X1 i_76 (.A(n_49), .B1(multiplier_M[25]), .B2(accumulator_A[25]), 
      .ZN(n_48));
   AOI21_X1 i_77 (.A(n_88), .B1(n_69), .B2(n_51), .ZN(n_49));
   OAI21_X1 i_78 (.A(n_69), .B1(multiplier_M[24]), .B2(accumulator_A[24]), 
      .ZN(n_50));
   INV_X1 i_79 (.A(n_52), .ZN(n_51));
   OAI21_X1 i_80 (.A(n_71), .B1(n_93), .B2(n_78), .ZN(n_52));
   OAI22_X1 i_81 (.A1(multiplier_M[27]), .A2(accumulator_A[27]), .B1(n_165), 
      .B2(n_162), .ZN(n_53));
   XNOR2_X1 i_82 (.A(n_64), .B(n_63), .ZN(p_0[28]));
   XOR2_X1 i_83 (.A(n_62), .B(n_58), .Z(p_0[29]));
   XNOR2_X1 i_84 (.A(n_55), .B(n_54), .ZN(p_0[30]));
   OAI21_X1 i_85 (.A(n_160), .B1(n_166), .B2(n_163), .ZN(n_54));
   NOR2_X1 i_86 (.A1(n_61), .A2(n_60), .ZN(n_55));
   XOR2_X1 i_87 (.A(n_57), .B(n_56), .Z(p_0[31]));
   XNOR2_X1 i_88 (.A(multiplier_M[31]), .B(multiplier_M[30]), .ZN(n_56));
   OAI21_X1 i_89 (.A(n_160), .B1(n_61), .B2(n_59), .ZN(n_57));
   AOI21_X1 i_90 (.A(n_60), .B1(multiplier_M[29]), .B2(accumulator_A[29]), 
      .ZN(n_58));
   OAI22_X1 i_91 (.A1(n_166), .A2(n_163), .B1(multiplier_M[29]), .B2(
      accumulator_A[29]), .ZN(n_59));
   NOR2_X1 i_92 (.A1(multiplier_M[29]), .A2(accumulator_A[29]), .ZN(n_60));
   AOI21_X1 i_93 (.A(n_62), .B1(multiplier_M[29]), .B2(accumulator_A[29]), 
      .ZN(n_61));
   AOI21_X1 i_94 (.A(n_159), .B1(n_64), .B2(n_63), .ZN(n_62));
   AOI21_X1 i_95 (.A(n_159), .B1(multiplier_M[28]), .B2(accumulator_A[28]), 
      .ZN(n_63));
   NOR4_X1 i_96 (.A1(n_67), .A2(n_65), .A3(n_70), .A4(n_77), .ZN(n_64));
   OAI22_X1 i_97 (.A1(n_165), .A2(n_162), .B1(n_92), .B2(n_66), .ZN(n_65));
   NAND2_X1 i_98 (.A1(multiplier_M[26]), .A2(accumulator_A[26]), .ZN(n_66));
   AOI21_X1 i_99 (.A(n_89), .B1(n_69), .B2(n_68), .ZN(n_67));
   NAND2_X1 i_100 (.A1(multiplier_M[25]), .A2(accumulator_A[25]), .ZN(n_68));
   NAND2_X1 i_101 (.A1(multiplier_M[24]), .A2(accumulator_A[24]), .ZN(n_69));
   NOR2_X1 i_102 (.A1(n_87), .A2(n_71), .ZN(n_70));
   AOI221_X1 i_103 (.A(n_73), .B1(multiplier_M[23]), .B2(accumulator_A[23]), 
      .C1(n_85), .C2(n_72), .ZN(n_71));
   AND2_X1 i_104 (.A1(multiplier_M[22]), .A2(accumulator_A[22]), .ZN(n_72));
   AOI21_X1 i_105 (.A(n_80), .B1(n_76), .B2(n_75), .ZN(n_73));
   INV_X1 i_106 (.A(n_75), .ZN(n_74));
   NAND2_X1 i_107 (.A1(multiplier_M[21]), .A2(accumulator_A[21]), .ZN(n_75));
   NAND2_X1 i_108 (.A1(multiplier_M[20]), .A2(accumulator_A[20]), .ZN(n_76));
   NOR3_X1 i_109 (.A1(n_87), .A2(n_78), .A3(n_93), .ZN(n_77));
   OR2_X1 i_110 (.A1(n_80), .A2(n_79), .ZN(n_78));
   NOR2_X1 i_111 (.A1(multiplier_M[20]), .A2(accumulator_A[20]), .ZN(n_79));
   NAND3_X1 i_112 (.A1(n_85), .A2(n_81), .A3(n_83), .ZN(n_80));
   INV_X1 i_113 (.A(n_82), .ZN(n_81));
   NOR2_X1 i_114 (.A1(multiplier_M[22]), .A2(accumulator_A[22]), .ZN(n_82));
   INV_X1 i_115 (.A(n_84), .ZN(n_83));
   NOR2_X1 i_116 (.A1(multiplier_M[21]), .A2(accumulator_A[21]), .ZN(n_84));
   INV_X1 i_117 (.A(n_86), .ZN(n_85));
   NOR2_X1 i_118 (.A1(multiplier_M[23]), .A2(accumulator_A[23]), .ZN(n_86));
   OR2_X1 i_119 (.A1(n_89), .A2(n_88), .ZN(n_87));
   NOR2_X1 i_120 (.A1(multiplier_M[24]), .A2(accumulator_A[24]), .ZN(n_88));
   OR2_X1 i_121 (.A1(n_92), .A2(n_90), .ZN(n_89));
   OAI22_X1 i_122 (.A1(multiplier_M[25]), .A2(accumulator_A[25]), .B1(
      multiplier_M[26]), .B2(accumulator_A[26]), .ZN(n_90));
   NOR2_X1 i_123 (.A1(multiplier_M[25]), .A2(accumulator_A[25]), .ZN(n_91));
   NOR2_X1 i_124 (.A1(multiplier_M[27]), .A2(accumulator_A[27]), .ZN(n_92));
   NOR4_X1 i_125 (.A1(n_97), .A2(n_94), .A3(n_98), .A4(n_101), .ZN(n_93));
   NOR2_X1 i_126 (.A1(n_106), .A2(n_96), .ZN(n_94));
   INV_X1 i_127 (.A(n_96), .ZN(n_95));
   NAND2_X1 i_128 (.A1(multiplier_M[18]), .A2(accumulator_A[18]), .ZN(n_96));
   AND2_X1 i_129 (.A1(multiplier_M[19]), .A2(accumulator_A[19]), .ZN(n_97));
   AOI21_X1 i_130 (.A(n_103), .B1(n_100), .B2(n_99), .ZN(n_98));
   NAND2_X1 i_131 (.A1(multiplier_M[17]), .A2(accumulator_A[17]), .ZN(n_99));
   NAND2_X1 i_132 (.A1(multiplier_M[16]), .A2(accumulator_A[16]), .ZN(n_100));
   NOR3_X1 i_133 (.A1(n_103), .A2(n_102), .A3(n_107), .ZN(n_101));
   NOR2_X1 i_134 (.A1(multiplier_M[16]), .A2(accumulator_A[16]), .ZN(n_102));
   OR3_X1 i_135 (.A1(n_106), .A2(n_104), .A3(n_105), .ZN(n_103));
   NOR2_X1 i_136 (.A1(multiplier_M[18]), .A2(accumulator_A[18]), .ZN(n_104));
   NOR2_X1 i_137 (.A1(multiplier_M[17]), .A2(accumulator_A[17]), .ZN(n_105));
   NOR2_X1 i_138 (.A1(multiplier_M[19]), .A2(accumulator_A[19]), .ZN(n_106));
   NOR4_X1 i_139 (.A1(n_111), .A2(n_108), .A3(n_112), .A4(n_115), .ZN(n_107));
   NOR2_X1 i_140 (.A1(n_120), .A2(n_110), .ZN(n_108));
   INV_X1 i_141 (.A(n_110), .ZN(n_109));
   NAND2_X1 i_142 (.A1(multiplier_M[14]), .A2(accumulator_A[14]), .ZN(n_110));
   AND2_X1 i_143 (.A1(multiplier_M[15]), .A2(accumulator_A[15]), .ZN(n_111));
   AOI21_X1 i_144 (.A(n_117), .B1(n_114), .B2(n_113), .ZN(n_112));
   NAND2_X1 i_145 (.A1(multiplier_M[13]), .A2(accumulator_A[13]), .ZN(n_113));
   NAND2_X1 i_146 (.A1(multiplier_M[12]), .A2(accumulator_A[12]), .ZN(n_114));
   NOR3_X1 i_147 (.A1(n_117), .A2(n_116), .A3(n_121), .ZN(n_115));
   NOR2_X1 i_148 (.A1(multiplier_M[12]), .A2(accumulator_A[12]), .ZN(n_116));
   OR3_X1 i_149 (.A1(n_120), .A2(n_118), .A3(n_119), .ZN(n_117));
   NOR2_X1 i_150 (.A1(multiplier_M[14]), .A2(accumulator_A[14]), .ZN(n_118));
   NOR2_X1 i_151 (.A1(multiplier_M[13]), .A2(accumulator_A[13]), .ZN(n_119));
   NOR2_X1 i_152 (.A1(multiplier_M[15]), .A2(accumulator_A[15]), .ZN(n_120));
   NOR4_X1 i_153 (.A1(n_125), .A2(n_122), .A3(n_126), .A4(n_129), .ZN(n_121));
   NOR2_X1 i_154 (.A1(n_134), .A2(n_124), .ZN(n_122));
   INV_X1 i_155 (.A(n_124), .ZN(n_123));
   NAND2_X1 i_156 (.A1(multiplier_M[10]), .A2(accumulator_A[10]), .ZN(n_124));
   AND2_X1 i_157 (.A1(multiplier_M[11]), .A2(accumulator_A[11]), .ZN(n_125));
   AOI21_X1 i_158 (.A(n_131), .B1(n_128), .B2(n_127), .ZN(n_126));
   NAND2_X1 i_159 (.A1(multiplier_M[9]), .A2(accumulator_A[9]), .ZN(n_127));
   NAND2_X1 i_160 (.A1(multiplier_M[8]), .A2(accumulator_A[8]), .ZN(n_128));
   NOR3_X1 i_161 (.A1(n_131), .A2(n_130), .A3(n_135), .ZN(n_129));
   NOR2_X1 i_162 (.A1(multiplier_M[8]), .A2(accumulator_A[8]), .ZN(n_130));
   OR3_X1 i_163 (.A1(n_134), .A2(n_132), .A3(n_133), .ZN(n_131));
   NOR2_X1 i_164 (.A1(multiplier_M[10]), .A2(accumulator_A[10]), .ZN(n_132));
   NOR2_X1 i_165 (.A1(multiplier_M[9]), .A2(accumulator_A[9]), .ZN(n_133));
   NOR2_X1 i_166 (.A1(multiplier_M[11]), .A2(accumulator_A[11]), .ZN(n_134));
   NOR4_X1 i_167 (.A1(n_139), .A2(n_136), .A3(n_140), .A4(n_143), .ZN(n_135));
   NOR2_X1 i_168 (.A1(n_148), .A2(n_138), .ZN(n_136));
   INV_X1 i_169 (.A(n_138), .ZN(n_137));
   NAND2_X1 i_170 (.A1(multiplier_M[6]), .A2(accumulator_A[6]), .ZN(n_138));
   AND2_X1 i_171 (.A1(multiplier_M[7]), .A2(accumulator_A[7]), .ZN(n_139));
   AOI21_X1 i_172 (.A(n_145), .B1(n_142), .B2(n_141), .ZN(n_140));
   NAND2_X1 i_173 (.A1(multiplier_M[5]), .A2(accumulator_A[5]), .ZN(n_141));
   NAND2_X1 i_174 (.A1(multiplier_M[4]), .A2(accumulator_A[4]), .ZN(n_142));
   NOR3_X1 i_175 (.A1(n_145), .A2(n_144), .A3(n_149), .ZN(n_143));
   NOR2_X1 i_176 (.A1(multiplier_M[4]), .A2(accumulator_A[4]), .ZN(n_144));
   OR3_X1 i_177 (.A1(n_148), .A2(n_146), .A3(n_147), .ZN(n_145));
   NOR2_X1 i_178 (.A1(multiplier_M[6]), .A2(accumulator_A[6]), .ZN(n_146));
   NOR2_X1 i_179 (.A1(multiplier_M[5]), .A2(accumulator_A[5]), .ZN(n_147));
   NOR2_X1 i_180 (.A1(multiplier_M[7]), .A2(accumulator_A[7]), .ZN(n_148));
   NAND2_X1 i_181 (.A1(n_158), .A2(n_150), .ZN(n_149));
   OAI21_X1 i_182 (.A(n_151), .B1(n_164), .B2(n_161), .ZN(n_150));
   OAI22_X1 i_183 (.A1(multiplier_M[2]), .A2(accumulator_A[2]), .B1(n_156), 
      .B2(n_152), .ZN(n_151));
   AOI21_X1 i_184 (.A(n_155), .B1(n_154), .B2(n_153), .ZN(n_152));
   NAND2_X1 i_185 (.A1(multiplier_M[1]), .A2(accumulator_A[1]), .ZN(n_153));
   NAND2_X1 i_186 (.A1(multiplier_M[0]), .A2(accumulator_A[0]), .ZN(n_154));
   NOR2_X1 i_187 (.A1(multiplier_M[1]), .A2(accumulator_A[1]), .ZN(n_155));
   INV_X1 i_188 (.A(n_157), .ZN(n_156));
   NAND2_X1 i_189 (.A1(multiplier_M[2]), .A2(accumulator_A[2]), .ZN(n_157));
   NAND2_X1 i_190 (.A1(n_164), .A2(n_161), .ZN(n_158));
   NOR2_X1 i_191 (.A1(multiplier_M[28]), .A2(accumulator_A[28]), .ZN(n_159));
   NAND2_X1 i_192 (.A1(n_166), .A2(n_163), .ZN(n_160));
   INV_X1 i_193 (.A(accumulator_A[3]), .ZN(n_161));
   INV_X1 i_194 (.A(accumulator_A[27]), .ZN(n_162));
   INV_X1 i_195 (.A(accumulator_A[30]), .ZN(n_163));
   INV_X1 i_196 (.A(multiplier_M[3]), .ZN(n_164));
   INV_X1 i_197 (.A(multiplier_M[27]), .ZN(n_165));
   INV_X1 i_198 (.A(multiplier_M[30]), .ZN(n_166));
endmodule

module datapath__0_5(accumulator_A, p_0, multiplier_M);
   input [31:0]accumulator_A;
   output [31:0]p_0;
   input [31:0]multiplier_M;

   OAI21_X1 i_0 (.A(n_25), .B1(n_38), .B2(multiplier_M[0]), .ZN(p_0[0]));
   XNOR2_X1 i_1 (.A(n_145), .B(n_0), .ZN(p_0[1]));
   NOR2_X1 i_2 (.A1(n_37), .A2(n_28), .ZN(n_0));
   XOR2_X1 i_3 (.A(n_3), .B(n_1), .Z(p_0[2]));
   NOR2_X1 i_4 (.A1(n_29), .A2(n_27), .ZN(n_1));
   XOR2_X1 i_5 (.A(n_4), .B(n_2), .Z(p_0[3]));
   OAI21_X1 i_6 (.A(n_34), .B1(n_27), .B2(n_3), .ZN(n_2));
   OAI22_X1 i_7 (.A1(n_43), .A2(multiplier_M[1]), .B1(n_37), .B2(n_145), 
      .ZN(n_3));
   OAI21_X1 i_8 (.A(n_36), .B1(n_45), .B2(multiplier_M[3]), .ZN(n_4));
   XNOR2_X1 i_9 (.A(n_11), .B(n_6), .ZN(p_0[5]));
   OAI21_X1 i_10 (.A(n_66), .B1(n_78), .B2(multiplier_M[5]), .ZN(n_6));
   XNOR2_X1 i_11 (.A(n_9), .B(n_7), .ZN(p_0[6]));
   OAI21_X1 i_12 (.A(n_68), .B1(n_79), .B2(multiplier_M[6]), .ZN(n_7));
   XOR2_X1 i_13 (.A(n_12), .B(n_8), .Z(p_0[7]));
   OAI21_X1 i_14 (.A(n_68), .B1(n_63), .B2(n_9), .ZN(n_8));
   INV_X1 i_15 (.A(n_10), .ZN(n_9));
   OAI21_X1 i_16 (.A(n_66), .B1(n_62), .B2(n_11), .ZN(n_10));
   OAI22_X1 i_17 (.A1(n_17), .A2(n_18), .B1(n_46), .B2(multiplier_M[4]), 
      .ZN(n_11));
   OAI21_X1 i_18 (.A(n_67), .B1(n_80), .B2(multiplier_M[7]), .ZN(n_12));
   XNOR2_X1 i_19 (.A(n_55), .B(n_13), .ZN(p_0[8]));
   NOR2_X1 i_20 (.A1(n_69), .A2(n_95), .ZN(n_13));
   XOR2_X1 i_21 (.A(n_54), .B(n_14), .Z(p_0[9]));
   NOR2_X1 i_22 (.A1(n_104), .A2(n_71), .ZN(n_14));
   XNOR2_X1 i_23 (.A(n_53), .B(n_15), .ZN(p_0[10]));
   NOR2_X1 i_24 (.A1(n_73), .A2(n_74), .ZN(n_15));
   XNOR2_X1 i_25 (.A(n_89), .B(n_20), .ZN(p_0[12]));
   OAI21_X1 i_26 (.A(n_97), .B1(n_107), .B2(multiplier_M[12]), .ZN(n_20));
   XNOR2_X1 i_27 (.A(n_88), .B(n_21), .ZN(p_0[13]));
   NOR2_X1 i_28 (.A1(n_132), .A2(n_98), .ZN(n_21));
   XNOR2_X1 i_29 (.A(n_86), .B(n_22), .ZN(p_0[14]));
   NOR2_X1 i_30 (.A1(n_100), .A2(n_101), .ZN(n_22));
   XNOR2_X1 i_31 (.A(n_117), .B(n_30), .ZN(p_0[16]));
   NOR2_X1 i_32 (.A1(n_116), .A2(n_151), .ZN(n_30));
   INV_X1 i_33 (.A(n_31), .ZN(p_0[17]));
   AOI21_X1 i_34 (.A(n_112), .B1(n_115), .B2(n_113), .ZN(n_31));
   XNOR2_X1 i_35 (.A(n_33), .B(n_32), .ZN(p_0[18]));
   OAI21_X1 i_36 (.A(n_126), .B1(n_114), .B2(n_115), .ZN(n_32));
   NOR2_X1 i_37 (.A1(n_125), .A2(n_127), .ZN(n_33));
   XOR2_X1 i_38 (.A(n_146), .B(n_39), .Z(p_0[20]));
   OAI22_X1 i_39 (.A1(accumulator_A[20]), .A2(n_159), .B1(n_161), .B2(
      multiplier_M[20]), .ZN(n_39));
   INV_X1 i_40 (.A(n_40), .ZN(p_0[21]));
   AOI21_X1 i_41 (.A(n_140), .B1(n_143), .B2(n_141), .ZN(n_40));
   XNOR2_X1 i_42 (.A(n_42), .B(n_41), .ZN(p_0[22]));
   OAI21_X1 i_43 (.A(n_154), .B1(n_142), .B2(n_143), .ZN(n_41));
   NOR2_X1 i_44 (.A1(n_153), .A2(n_155), .ZN(n_42));
   XOR2_X1 i_45 (.A(n_170), .B(n_48), .Z(p_0[24]));
   OAI22_X1 i_46 (.A1(accumulator_A[24]), .A2(n_181), .B1(n_183), .B2(
      multiplier_M[24]), .ZN(n_48));
   INV_X1 i_47 (.A(n_49), .ZN(p_0[25]));
   AOI21_X1 i_48 (.A(n_165), .B1(n_168), .B2(n_166), .ZN(n_49));
   XNOR2_X1 i_49 (.A(n_51), .B(n_50), .ZN(p_0[26]));
   OAI21_X1 i_50 (.A(n_178), .B1(n_167), .B2(n_168), .ZN(n_50));
   NOR2_X1 i_51 (.A1(n_177), .A2(n_179), .ZN(n_51));
   XOR2_X1 i_52 (.A(n_56), .B(n_164), .Z(p_0[27]));
   NOR2_X1 i_53 (.A1(n_196), .A2(n_197), .ZN(n_56));
   XOR2_X1 i_54 (.A(multiplier_M[28]), .B(n_57), .Z(p_0[28]));
   OAI21_X1 i_55 (.A(n_191), .B1(accumulator_A[28]), .B2(n_192), .ZN(n_57));
   XOR2_X1 i_56 (.A(n_189), .B(n_206), .Z(p_0[29]));
   XOR2_X1 i_57 (.A(n_204), .B(n_60), .Z(p_0[31]));
   XOR2_X1 i_58 (.A(accumulator_A[30]), .B(multiplier_M[31]), .Z(n_60));
   INV_X1 i_59 (.A(n_25), .ZN(n_145));
   XNOR2_X1 i_60 (.A(n_19), .B(n_5), .ZN(p_0[4]));
   OR2_X1 i_61 (.A1(n_17), .A2(n_16), .ZN(n_5));
   NOR2_X1 i_62 (.A1(n_46), .A2(multiplier_M[4]), .ZN(n_16));
   AND2_X1 i_63 (.A1(n_46), .A2(multiplier_M[4]), .ZN(n_17));
   INV_X1 i_64 (.A(n_19), .ZN(n_18));
   OAI221_X1 i_65 (.A(n_23), .B1(n_45), .B2(multiplier_M[3]), .C1(n_35), 
      .C2(n_26), .ZN(n_19));
   OAI21_X1 i_66 (.A(n_24), .B1(n_28), .B2(n_25), .ZN(n_23));
   NOR3_X1 i_67 (.A1(n_35), .A2(n_29), .A3(n_37), .ZN(n_24));
   NAND2_X1 i_68 (.A1(n_38), .A2(multiplier_M[0]), .ZN(n_25));
   INV_X1 i_69 (.A(n_27), .ZN(n_26));
   NOR2_X1 i_70 (.A1(n_44), .A2(multiplier_M[2]), .ZN(n_27));
   NOR2_X1 i_71 (.A1(n_43), .A2(multiplier_M[1]), .ZN(n_28));
   INV_X1 i_72 (.A(n_34), .ZN(n_29));
   NAND2_X1 i_73 (.A1(n_44), .A2(multiplier_M[2]), .ZN(n_34));
   INV_X1 i_74 (.A(n_36), .ZN(n_35));
   NAND2_X1 i_75 (.A1(n_45), .A2(multiplier_M[3]), .ZN(n_36));
   AND2_X1 i_76 (.A1(n_43), .A2(multiplier_M[1]), .ZN(n_37));
   INV_X1 i_77 (.A(accumulator_A[0]), .ZN(n_38));
   INV_X1 i_78 (.A(accumulator_A[1]), .ZN(n_43));
   INV_X1 i_79 (.A(accumulator_A[2]), .ZN(n_44));
   INV_X1 i_80 (.A(accumulator_A[3]), .ZN(n_45));
   INV_X1 i_81 (.A(accumulator_A[4]), .ZN(n_46));
   XNOR2_X1 i_82 (.A(n_52), .B(n_47), .ZN(p_0[11]));
   OAI21_X1 i_83 (.A(n_75), .B1(n_73), .B2(n_53), .ZN(n_47));
   OAI21_X1 i_84 (.A(n_76), .B1(n_83), .B2(multiplier_M[11]), .ZN(n_52));
   OAI21_X1 i_85 (.A(n_72), .B1(n_71), .B2(n_54), .ZN(n_53));
   OAI22_X1 i_86 (.A1(n_81), .A2(multiplier_M[8]), .B1(n_69), .B2(n_55), 
      .ZN(n_54));
   NOR2_X1 i_87 (.A1(n_64), .A2(n_58), .ZN(n_55));
   OAI221_X1 i_88 (.A(n_59), .B1(n_65), .B2(n_61), .C1(n_80), .C2(
      multiplier_M[7]), .ZN(n_58));
   NAND2_X1 i_89 (.A1(n_67), .A2(n_63), .ZN(n_59));
   NOR2_X1 i_90 (.A1(n_16), .A2(n_62), .ZN(n_61));
   NOR2_X1 i_91 (.A1(n_78), .A2(multiplier_M[5]), .ZN(n_62));
   NOR2_X1 i_92 (.A1(n_79), .A2(multiplier_M[6]), .ZN(n_63));
   NOR3_X1 i_93 (.A1(n_17), .A2(n_65), .A3(n_18), .ZN(n_64));
   NAND3_X1 i_94 (.A1(n_68), .A2(n_66), .A3(n_67), .ZN(n_65));
   NAND2_X1 i_95 (.A1(n_78), .A2(multiplier_M[5]), .ZN(n_66));
   NAND2_X1 i_96 (.A1(n_80), .A2(multiplier_M[7]), .ZN(n_67));
   NAND2_X1 i_97 (.A1(n_79), .A2(multiplier_M[6]), .ZN(n_68));
   INV_X1 i_98 (.A(n_70), .ZN(n_69));
   NAND2_X1 i_99 (.A1(n_81), .A2(multiplier_M[8]), .ZN(n_70));
   NOR2_X1 i_100 (.A1(n_82), .A2(multiplier_M[9]), .ZN(n_71));
   NAND2_X1 i_101 (.A1(n_82), .A2(multiplier_M[9]), .ZN(n_72));
   NOR2_X1 i_102 (.A1(accumulator_A[10]), .A2(n_77), .ZN(n_73));
   INV_X1 i_103 (.A(n_75), .ZN(n_74));
   NAND2_X1 i_104 (.A1(accumulator_A[10]), .A2(n_77), .ZN(n_75));
   NAND2_X1 i_105 (.A1(n_83), .A2(multiplier_M[11]), .ZN(n_76));
   INV_X1 i_106 (.A(multiplier_M[10]), .ZN(n_77));
   INV_X1 i_107 (.A(accumulator_A[5]), .ZN(n_78));
   INV_X1 i_108 (.A(accumulator_A[6]), .ZN(n_79));
   INV_X1 i_109 (.A(accumulator_A[7]), .ZN(n_80));
   INV_X1 i_110 (.A(accumulator_A[8]), .ZN(n_81));
   INV_X1 i_111 (.A(accumulator_A[9]), .ZN(n_82));
   INV_X1 i_112 (.A(accumulator_A[11]), .ZN(n_83));
   XNOR2_X1 i_113 (.A(n_85), .B(n_84), .ZN(p_0[15]));
   OAI21_X1 i_114 (.A(n_102), .B1(n_100), .B2(n_86), .ZN(n_84));
   OAI21_X1 i_115 (.A(n_103), .B1(n_109), .B2(multiplier_M[15]), .ZN(n_85));
   OAI21_X1 i_116 (.A(n_99), .B1(n_98), .B2(n_87), .ZN(n_86));
   INV_X1 i_117 (.A(n_88), .ZN(n_87));
   OAI21_X1 i_118 (.A(n_97), .B1(n_96), .B2(n_89), .ZN(n_88));
   OAI21_X1 i_119 (.A(n_91), .B1(n_55), .B2(n_90), .ZN(n_89));
   NAND2_X1 i_120 (.A1(n_70), .A2(n_94), .ZN(n_90));
   INV_X1 i_121 (.A(n_92), .ZN(n_91));
   OAI221_X1 i_122 (.A(n_93), .B1(multiplier_M[11]), .B2(n_83), .C1(n_105), 
      .C2(n_75), .ZN(n_92));
   OAI21_X1 i_123 (.A(n_94), .B1(n_71), .B2(n_95), .ZN(n_93));
   NOR3_X1 i_124 (.A1(n_105), .A2(n_73), .A3(n_104), .ZN(n_94));
   NOR2_X1 i_125 (.A1(multiplier_M[8]), .A2(n_81), .ZN(n_95));
   NOR2_X1 i_126 (.A1(n_107), .A2(multiplier_M[12]), .ZN(n_96));
   NAND2_X1 i_127 (.A1(n_107), .A2(multiplier_M[12]), .ZN(n_97));
   NOR2_X1 i_128 (.A1(n_108), .A2(multiplier_M[13]), .ZN(n_98));
   NAND2_X1 i_129 (.A1(n_108), .A2(multiplier_M[13]), .ZN(n_99));
   NOR2_X1 i_130 (.A1(accumulator_A[14]), .A2(n_106), .ZN(n_100));
   INV_X1 i_131 (.A(n_102), .ZN(n_101));
   NAND2_X1 i_132 (.A1(accumulator_A[14]), .A2(n_106), .ZN(n_102));
   NAND2_X1 i_133 (.A1(n_109), .A2(multiplier_M[15]), .ZN(n_103));
   INV_X1 i_134 (.A(n_72), .ZN(n_104));
   INV_X1 i_135 (.A(n_76), .ZN(n_105));
   INV_X1 i_136 (.A(multiplier_M[14]), .ZN(n_106));
   INV_X1 i_137 (.A(accumulator_A[12]), .ZN(n_107));
   INV_X1 i_138 (.A(accumulator_A[13]), .ZN(n_108));
   INV_X1 i_139 (.A(accumulator_A[15]), .ZN(n_109));
   XNOR2_X1 i_140 (.A(n_111), .B(n_110), .ZN(p_0[19]));
   OAI21_X1 i_141 (.A(n_128), .B1(n_124), .B2(n_112), .ZN(n_110));
   OR2_X1 i_142 (.A1(n_130), .A2(n_129), .ZN(n_111));
   NOR2_X1 i_143 (.A1(n_115), .A2(n_113), .ZN(n_112));
   OAI21_X1 i_144 (.A(n_126), .B1(n_136), .B2(multiplier_M[17]), .ZN(n_113));
   NOR2_X1 i_145 (.A1(n_136), .A2(multiplier_M[17]), .ZN(n_114));
   OAI22_X1 i_146 (.A1(n_135), .A2(multiplier_M[16]), .B1(n_117), .B2(n_116), 
      .ZN(n_115));
   AND2_X1 i_147 (.A1(n_135), .A2(multiplier_M[16]), .ZN(n_116));
   AOI221_X1 i_148 (.A(n_118), .B1(n_131), .B2(n_122), .C1(n_122), .C2(n_120), 
      .ZN(n_117));
   OAI221_X1 i_149 (.A(n_119), .B1(n_133), .B2(n_102), .C1(multiplier_M[15]), 
      .C2(n_109), .ZN(n_118));
   OAI21_X1 i_150 (.A(n_123), .B1(n_96), .B2(n_98), .ZN(n_119));
   NOR2_X1 i_151 (.A1(n_90), .A2(n_121), .ZN(n_120));
   NOR2_X1 i_152 (.A1(n_58), .A2(n_64), .ZN(n_121));
   AND2_X1 i_153 (.A1(n_97), .A2(n_123), .ZN(n_122));
   NOR3_X1 i_154 (.A1(n_133), .A2(n_100), .A3(n_132), .ZN(n_123));
   OAI21_X1 i_155 (.A(n_126), .B1(accumulator_A[18]), .B2(n_134), .ZN(n_124));
   NOR2_X1 i_156 (.A1(accumulator_A[18]), .A2(n_134), .ZN(n_125));
   NAND2_X1 i_157 (.A1(n_136), .A2(multiplier_M[17]), .ZN(n_126));
   INV_X1 i_158 (.A(n_128), .ZN(n_127));
   NAND2_X1 i_159 (.A1(accumulator_A[18]), .A2(n_134), .ZN(n_128));
   NOR2_X1 i_160 (.A1(n_137), .A2(multiplier_M[19]), .ZN(n_129));
   AND2_X1 i_161 (.A1(n_137), .A2(multiplier_M[19]), .ZN(n_130));
   INV_X1 i_162 (.A(n_91), .ZN(n_131));
   INV_X1 i_163 (.A(n_99), .ZN(n_132));
   INV_X1 i_164 (.A(n_103), .ZN(n_133));
   INV_X1 i_165 (.A(multiplier_M[18]), .ZN(n_134));
   INV_X1 i_166 (.A(accumulator_A[16]), .ZN(n_135));
   INV_X1 i_167 (.A(accumulator_A[17]), .ZN(n_136));
   INV_X1 i_168 (.A(accumulator_A[19]), .ZN(n_137));
   XNOR2_X1 i_169 (.A(n_139), .B(n_138), .ZN(p_0[23]));
   OAI21_X1 i_170 (.A(n_156), .B1(n_152), .B2(n_140), .ZN(n_138));
   OR2_X1 i_171 (.A1(n_158), .A2(n_157), .ZN(n_139));
   NOR2_X1 i_172 (.A1(n_143), .A2(n_141), .ZN(n_140));
   OAI21_X1 i_173 (.A(n_154), .B1(n_162), .B2(multiplier_M[21]), .ZN(n_141));
   NOR2_X1 i_174 (.A1(n_162), .A2(multiplier_M[21]), .ZN(n_142));
   OAI22_X1 i_175 (.A1(n_161), .A2(multiplier_M[20]), .B1(n_146), .B2(n_144), 
      .ZN(n_143));
   NOR2_X1 i_176 (.A1(accumulator_A[20]), .A2(n_159), .ZN(n_144));
   NOR4_X1 i_177 (.A1(n_129), .A2(n_147), .A3(n_149), .A4(n_148), .ZN(n_146));
   NOR2_X1 i_178 (.A1(n_130), .A2(n_128), .ZN(n_147));
   NOR4_X1 i_179 (.A1(n_130), .A2(n_124), .A3(n_116), .A4(n_117), .ZN(n_148));
   NOR3_X1 i_180 (.A1(n_130), .A2(n_124), .A3(n_150), .ZN(n_149));
   NOR2_X1 i_181 (.A1(n_114), .A2(n_151), .ZN(n_150));
   NOR2_X1 i_182 (.A1(multiplier_M[16]), .A2(n_135), .ZN(n_151));
   OAI21_X1 i_183 (.A(n_154), .B1(accumulator_A[22]), .B2(n_160), .ZN(n_152));
   NOR2_X1 i_184 (.A1(accumulator_A[22]), .A2(n_160), .ZN(n_153));
   NAND2_X1 i_185 (.A1(n_162), .A2(multiplier_M[21]), .ZN(n_154));
   INV_X1 i_186 (.A(n_156), .ZN(n_155));
   NAND2_X1 i_187 (.A1(accumulator_A[22]), .A2(n_160), .ZN(n_156));
   NOR2_X1 i_188 (.A1(n_163), .A2(multiplier_M[23]), .ZN(n_157));
   AND2_X1 i_189 (.A1(n_163), .A2(multiplier_M[23]), .ZN(n_158));
   INV_X1 i_190 (.A(multiplier_M[20]), .ZN(n_159));
   INV_X1 i_191 (.A(multiplier_M[22]), .ZN(n_160));
   INV_X1 i_192 (.A(accumulator_A[20]), .ZN(n_161));
   INV_X1 i_193 (.A(accumulator_A[21]), .ZN(n_162));
   INV_X1 i_194 (.A(accumulator_A[23]), .ZN(n_163));
   OAI21_X1 i_195 (.A(n_180), .B1(n_176), .B2(n_165), .ZN(n_164));
   NOR2_X1 i_196 (.A1(n_168), .A2(n_166), .ZN(n_165));
   OAI21_X1 i_197 (.A(n_178), .B1(n_184), .B2(multiplier_M[25]), .ZN(n_166));
   NOR2_X1 i_198 (.A1(n_184), .A2(multiplier_M[25]), .ZN(n_167));
   OAI22_X1 i_199 (.A1(n_183), .A2(multiplier_M[24]), .B1(n_170), .B2(n_169), 
      .ZN(n_168));
   NOR2_X1 i_200 (.A1(accumulator_A[24]), .A2(n_181), .ZN(n_169));
   NOR4_X1 i_201 (.A1(n_157), .A2(n_171), .A3(n_173), .A4(n_172), .ZN(n_170));
   NOR2_X1 i_202 (.A1(n_158), .A2(n_156), .ZN(n_171));
   NOR3_X1 i_203 (.A1(n_144), .A2(n_175), .A3(n_146), .ZN(n_172));
   NOR2_X1 i_204 (.A1(n_175), .A2(n_174), .ZN(n_173));
   AOI21_X1 i_205 (.A(n_142), .B1(accumulator_A[20]), .B2(n_159), .ZN(n_174));
   OR2_X1 i_206 (.A1(n_158), .A2(n_152), .ZN(n_175));
   OAI21_X1 i_207 (.A(n_178), .B1(accumulator_A[26]), .B2(n_182), .ZN(n_176));
   NOR2_X1 i_208 (.A1(accumulator_A[26]), .A2(n_182), .ZN(n_177));
   NAND2_X1 i_209 (.A1(n_184), .A2(multiplier_M[25]), .ZN(n_178));
   INV_X1 i_210 (.A(n_180), .ZN(n_179));
   NAND2_X1 i_211 (.A1(accumulator_A[26]), .A2(n_182), .ZN(n_180));
   INV_X1 i_212 (.A(multiplier_M[24]), .ZN(n_181));
   INV_X1 i_213 (.A(multiplier_M[26]), .ZN(n_182));
   INV_X1 i_214 (.A(accumulator_A[24]), .ZN(n_183));
   INV_X1 i_215 (.A(accumulator_A[25]), .ZN(n_184));
   XNOR2_X1 i_216 (.A(n_186), .B(n_185), .ZN(p_0[30]));
   OAI22_X1 i_217 (.A1(multiplier_M[29]), .A2(n_200), .B1(n_189), .B2(n_187), 
      .ZN(n_185));
   OAI21_X1 i_218 (.A(n_199), .B1(n_203), .B2(accumulator_A[30]), .ZN(n_186));
   INV_X1 i_219 (.A(n_188), .ZN(n_187));
   NAND2_X1 i_220 (.A1(multiplier_M[29]), .A2(n_200), .ZN(n_188));
   OAI22_X1 i_221 (.A1(accumulator_A[28]), .A2(n_192), .B1(n_202), .B2(n_190), 
      .ZN(n_189));
   INV_X1 i_222 (.A(n_191), .ZN(n_190));
   NAND2_X1 i_223 (.A1(accumulator_A[28]), .A2(n_192), .ZN(n_191));
   OAI221_X1 i_224 (.A(n_198), .B1(n_180), .B2(n_196), .C1(n_195), .C2(n_193), 
      .ZN(n_192));
   AOI211_X1 i_225 (.A(n_167), .B(n_194), .C1(accumulator_A[24]), .C2(n_181), 
      .ZN(n_193));
   NOR2_X1 i_226 (.A1(n_169), .A2(n_170), .ZN(n_194));
   OR2_X1 i_227 (.A1(n_176), .A2(n_196), .ZN(n_195));
   NOR2_X1 i_228 (.A1(n_201), .A2(accumulator_A[27]), .ZN(n_196));
   INV_X1 i_229 (.A(n_198), .ZN(n_197));
   NAND2_X1 i_230 (.A1(n_201), .A2(accumulator_A[27]), .ZN(n_198));
   NAND2_X1 i_231 (.A1(n_203), .A2(accumulator_A[30]), .ZN(n_199));
   INV_X1 i_232 (.A(accumulator_A[29]), .ZN(n_200));
   INV_X1 i_233 (.A(multiplier_M[27]), .ZN(n_201));
   INV_X1 i_234 (.A(multiplier_M[28]), .ZN(n_202));
   INV_X1 i_235 (.A(multiplier_M[30]), .ZN(n_203));
   OAI222_X1 i_236 (.A1(accumulator_A[30]), .A2(n_203), .B1(n_188), .B2(n_207), 
      .C1(n_206), .C2(n_205), .ZN(n_204));
   NAND2_X1 i_237 (.A1(n_199), .A2(n_189), .ZN(n_205));
   OAI21_X1 i_238 (.A(n_188), .B1(n_200), .B2(multiplier_M[29]), .ZN(n_206));
   INV_X1 i_239 (.A(n_199), .ZN(n_207));
endmodule

module boothAlgo(Res, OVF, A, B, clk, reset, enable);
   output [63:0]Res;
   output OVF;
   input [31:0]A;
   input [31:0]B;
   input clk;
   input reset;
   input enable;

   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire [1:0]isNeg;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire [31:0]accumulator_A;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_0;
   wire [31:0]multiplier_M;
   wire ready;
   wire [4:0]counter;
   wire n_0_221;
   wire n_0_222;
   wire n_0_2_0;
   wire n_0_223;
   wire n_0_224;
   wire n_0_2_1;
   wire n_0_225;
   wire n_0_2_2;
   wire n_0_226;
   wire n_0_2_3;
   wire n_0_227;
   wire n_0_2_4;
   wire n_0_2_5;
   wire n_0_2_6;
   wire n_0_2_7;
   wire n_0_228;
   wire n_0_2_8;
   wire n_0_229;
   wire n_0_2_9;
   wire n_0_230;
   wire n_0_2_10;
   wire n_0_231;
   wire n_0_2_11;
   wire n_0_232;
   wire n_0_2_12;
   wire n_0_233;
   wire n_0_2_13;
   wire n_0_234;
   wire n_0_2_14;
   wire n_0_235;
   wire n_0_2_15;
   wire n_0_236;
   wire n_0_2_16;
   wire n_0_237;
   wire n_0_2_17;
   wire n_0_238;
   wire n_0_2_18;
   wire n_0_239;
   wire n_0_2_19;
   wire n_0_240;
   wire n_0_2_20;
   wire n_0_241;
   wire n_0_2_21;
   wire n_0_242;
   wire n_0_2_22;
   wire n_0_243;
   wire n_0_2_23;
   wire n_0_244;
   wire n_0_2_24;
   wire n_0_245;
   wire n_0_2_25;
   wire n_0_246;
   wire n_0_2_26;
   wire n_0_247;
   wire n_0_2_27;
   wire n_0_248;
   wire n_0_2_28;
   wire n_0_249;
   wire n_0_2_29;
   wire n_0_250;
   wire n_0_2_30;
   wire n_0_251;
   wire n_0_2_31;
   wire n_0_252;
   wire n_0_2_32;
   wire n_0_253;
   wire n_0_2_33;
   wire n_0_254;
   wire n_0_2_34;
   wire n_0_255;
   wire n_0_2_35;
   wire n_0_256;
   wire n_0_2_36;
   wire n_0_257;
   wire n_0_2_37;
   wire n_0_258;
   wire n_0_2_38;
   wire n_0_259;
   wire n_0_2_39;
   wire n_0_261;
   wire n_0_2_40;
   wire n_0_262;
   wire n_0_2_41;
   wire n_0_263;
   wire n_0_2_42;
   wire n_0_264;
   wire n_0_2_43;
   wire n_0_265;
   wire n_0_2_44;
   wire n_0_266;
   wire n_0_2_45;
   wire n_0_267;
   wire n_0_2_46;
   wire n_0_268;
   wire n_0_2_47;
   wire n_0_269;
   wire n_0_2_48;
   wire n_0_270;
   wire n_0_2_49;
   wire n_0_271;
   wire n_0_2_50;
   wire n_0_272;
   wire n_0_2_51;
   wire n_0_273;
   wire n_0_2_52;
   wire n_0_274;
   wire n_0_2_53;
   wire n_0_275;
   wire n_0_2_54;
   wire n_0_276;
   wire n_0_2_55;
   wire n_0_277;
   wire n_0_2_56;
   wire n_0_278;
   wire n_0_2_57;
   wire n_0_279;
   wire n_0_2_58;
   wire n_0_280;
   wire n_0_2_59;
   wire n_0_281;
   wire n_0_2_60;
   wire n_0_282;
   wire n_0_2_61;
   wire n_0_283;
   wire n_0_2_62;
   wire n_0_284;
   wire n_0_2_63;
   wire n_0_285;
   wire n_0_2_64;
   wire n_0_286;
   wire n_0_2_65;
   wire n_0_287;
   wire n_0_2_66;
   wire n_0_288;
   wire n_0_2_67;
   wire n_0_289;
   wire n_0_2_68;
   wire n_0_290;
   wire n_0_2_69;
   wire n_0_291;
   wire n_0_2_70;
   wire n_0_2_71;
   wire n_0_292;
   wire n_0_2_72;
   wire n_0_2_73;
   wire n_0_2_74;
   wire n_0_2_75;
   wire n_0_260;
   wire n_0_2_76;
   wire n_0_2_77;
   wire n_0_2_78;
   wire n_0_293;
   wire n_0_294;
   wire n_0_2_79;
   wire n_0_295;
   wire n_0_2_80;
   wire n_0_296;
   wire n_0_2_81;
   wire n_0_297;
   wire n_0_2_82;
   wire n_0_298;
   wire n_0_2_83;
   wire n_0_299;
   wire n_0_2_84;
   wire n_0_300;
   wire n_0_2_85;
   wire n_0_301;
   wire n_0_2_86;
   wire n_0_302;
   wire n_0_2_87;
   wire n_0_303;
   wire n_0_2_88;
   wire n_0_304;
   wire n_0_2_89;
   wire n_0_305;
   wire n_0_2_90;
   wire n_0_306;
   wire n_0_2_91;
   wire n_0_307;
   wire n_0_2_92;
   wire n_0_308;
   wire n_0_2_93;
   wire n_0_309;
   wire n_0_2_94;
   wire n_0_310;
   wire n_0_2_95;
   wire n_0_311;
   wire n_0_2_96;
   wire n_0_312;
   wire n_0_2_97;
   wire n_0_313;
   wire n_0_2_98;
   wire n_0_314;
   wire n_0_2_99;
   wire n_0_315;
   wire n_0_2_100;
   wire n_0_316;
   wire n_0_2_101;
   wire n_0_317;
   wire n_0_2_102;
   wire n_0_318;
   wire n_0_2_103;
   wire n_0_319;
   wire n_0_2_104;
   wire n_0_320;
   wire n_0_2_105;
   wire n_0_321;
   wire n_0_2_106;
   wire n_0_322;
   wire n_0_2_107;
   wire n_0_323;
   wire n_0_2_108;
   wire n_0_2_109;
   wire n_0_324;
   wire n_0_325;
   wire n_0_2_110;
   wire n_0_2_111;
   wire n_0_326;
   wire n_0_327;
   wire n_0_2_112;
   wire n_0_2_113;
   wire n_0_2_114;
   wire n_0_2_115;
   wire n_0_2_116;
   wire n_0_2_117;
   wire n_0_2_118;
   wire n_0_2_119;
   wire n_0_2_120;
   wire n_0_2_121;
   wire n_0_2_122;
   wire n_0_2_123;
   wire n_0_2_124;
   wire n_0_2_125;
   wire n_0_2_126;
   wire n_0_2_127;
   wire n_0_2_128;
   wire n_0_2_129;
   wire n_0_2_130;
   wire n_0_2_131;
   wire n_0_2_132;
   wire n_0_2_133;
   wire n_0_2_134;
   wire n_0_2_135;
   wire n_0_2_136;
   wire n_0_2_137;
   wire n_0_2_138;
   wire n_0_2_139;
   wire n_0_2_140;

   datapath i_0_0 (.B(B), .p_0({n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, 
      n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, 
      n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, 
      n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, uc_0}));
   datapath__0_0 i_0_1 (.A(A), .p_0({n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, 
      n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, 
      n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, 
      n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, uc_1}));
   datapath__0_17 i_0_3 (.p_0({accumulator_A[30], uc_2, accumulator_A[29], 
      accumulator_A[28], accumulator_A[27], accumulator_A[26], accumulator_A[25], 
      accumulator_A[24], accumulator_A[23], accumulator_A[22], accumulator_A[21], 
      accumulator_A[20], accumulator_A[19], accumulator_A[18], accumulator_A[17], 
      accumulator_A[16], accumulator_A[15], accumulator_A[14], accumulator_A[13], 
      accumulator_A[12], accumulator_A[11], accumulator_A[10], accumulator_A[9], 
      accumulator_A[8], accumulator_A[7], accumulator_A[6], accumulator_A[5], 
      accumulator_A[4], accumulator_A[3], accumulator_A[2], accumulator_A[1], 
      accumulator_A[0], n_0_190, n_0_191, n_0_192, n_0_193, n_0_194, n_0_195, 
      n_0_196, n_0_197, n_0_198, n_0_199, n_0_200, n_0_201, n_0_202, n_0_203, 
      n_0_204, n_0_205, n_0_206, n_0_207, n_0_208, n_0_209, n_0_210, n_0_211, 
      n_0_212, n_0_213, n_0_214, n_0_215, n_0_216, n_0_217, n_0_218, n_0_219, 
      n_0_220, Res[0]}), .p_1({n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, 
      n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, 
      n_0_112, n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, 
      n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, 
      n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, 
      n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, 
      n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, 
      n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, uc_3}));
   DLH_X1 \isNeg_reg[1]  (.D(n_0_327), .G(n_0_325), .Q(isNeg[1]));
   DLH_X1 \isNeg_reg[0]  (.D(n_0_326), .G(n_0_325), .Q(isNeg[0]));
   datapath__0_4 i_0_12 (.multiplier_M(multiplier_M), .accumulator_A({uc_4, 
      accumulator_A[30], accumulator_A[29], accumulator_A[28], accumulator_A[27], 
      accumulator_A[26], accumulator_A[25], accumulator_A[24], accumulator_A[23], 
      accumulator_A[22], accumulator_A[21], accumulator_A[20], accumulator_A[19], 
      accumulator_A[18], accumulator_A[17], accumulator_A[16], accumulator_A[15], 
      accumulator_A[14], accumulator_A[13], accumulator_A[12], accumulator_A[11], 
      accumulator_A[10], accumulator_A[9], accumulator_A[8], accumulator_A[7], 
      accumulator_A[6], accumulator_A[5], accumulator_A[4], accumulator_A[3], 
      accumulator_A[2], accumulator_A[1], accumulator_A[0]}), .p_0({n_0_157, 
      n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, n_0_151, n_0_150, n_0_149, 
      n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, n_0_143, n_0_142, n_0_141, 
      n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, n_0_133, 
      n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, n_0_126}));
   datapath__0_5 i_0_13 (.accumulator_A({uc_5, accumulator_A[30], 
      accumulator_A[29], accumulator_A[28], accumulator_A[27], accumulator_A[26], 
      accumulator_A[25], accumulator_A[24], accumulator_A[23], accumulator_A[22], 
      accumulator_A[21], accumulator_A[20], accumulator_A[19], accumulator_A[18], 
      accumulator_A[17], accumulator_A[16], accumulator_A[15], accumulator_A[14], 
      accumulator_A[13], accumulator_A[12], accumulator_A[11], accumulator_A[10], 
      accumulator_A[9], accumulator_A[8], accumulator_A[7], accumulator_A[6], 
      accumulator_A[5], accumulator_A[4], accumulator_A[3], accumulator_A[2], 
      accumulator_A[1], accumulator_A[0]}), .p_0({n_0_189, n_0_188, n_0_187, 
      n_0_186, n_0_185, n_0_184, n_0_183, n_0_182, n_0_181, n_0_180, n_0_179, 
      n_0_178, n_0_177, n_0_176, n_0_175, n_0_174, n_0_173, n_0_172, n_0_171, 
      n_0_170, n_0_169, n_0_168, n_0_167, n_0_166, n_0_165, n_0_164, n_0_163, 
      n_0_162, n_0_161, n_0_160, n_0_159, n_0_158}), .multiplier_M(multiplier_M));
   DLH_X1 \accumulator_A_reg[30]  (.D(n_0_259), .G(n_0_228), .Q(
      accumulator_A[30]));
   DLH_X1 \accumulator_A_reg[29]  (.D(n_0_258), .G(n_0_228), .Q(
      accumulator_A[29]));
   DLH_X1 \accumulator_A_reg[28]  (.D(n_0_257), .G(n_0_228), .Q(
      accumulator_A[28]));
   DLH_X1 \accumulator_A_reg[27]  (.D(n_0_256), .G(n_0_228), .Q(
      accumulator_A[27]));
   DLH_X1 \accumulator_A_reg[26]  (.D(n_0_255), .G(n_0_228), .Q(
      accumulator_A[26]));
   DLH_X1 \accumulator_A_reg[25]  (.D(n_0_254), .G(n_0_228), .Q(
      accumulator_A[25]));
   DLH_X1 \accumulator_A_reg[24]  (.D(n_0_253), .G(n_0_228), .Q(
      accumulator_A[24]));
   DLH_X1 \accumulator_A_reg[23]  (.D(n_0_252), .G(n_0_228), .Q(
      accumulator_A[23]));
   DLH_X1 \accumulator_A_reg[22]  (.D(n_0_251), .G(n_0_228), .Q(
      accumulator_A[22]));
   DLH_X1 \accumulator_A_reg[21]  (.D(n_0_250), .G(n_0_228), .Q(
      accumulator_A[21]));
   DLH_X1 \accumulator_A_reg[20]  (.D(n_0_249), .G(n_0_228), .Q(
      accumulator_A[20]));
   DLH_X1 \accumulator_A_reg[19]  (.D(n_0_248), .G(n_0_228), .Q(
      accumulator_A[19]));
   DLH_X1 \accumulator_A_reg[18]  (.D(n_0_247), .G(n_0_228), .Q(
      accumulator_A[18]));
   DLH_X1 \accumulator_A_reg[17]  (.D(n_0_246), .G(n_0_228), .Q(
      accumulator_A[17]));
   DLH_X1 \accumulator_A_reg[16]  (.D(n_0_245), .G(n_0_228), .Q(
      accumulator_A[16]));
   DLH_X1 \accumulator_A_reg[15]  (.D(n_0_244), .G(n_0_228), .Q(
      accumulator_A[15]));
   DLH_X1 \accumulator_A_reg[14]  (.D(n_0_243), .G(n_0_228), .Q(
      accumulator_A[14]));
   DLH_X1 \accumulator_A_reg[13]  (.D(n_0_242), .G(n_0_228), .Q(
      accumulator_A[13]));
   DLH_X1 \accumulator_A_reg[12]  (.D(n_0_241), .G(n_0_228), .Q(
      accumulator_A[12]));
   DLH_X1 \accumulator_A_reg[11]  (.D(n_0_240), .G(n_0_228), .Q(
      accumulator_A[11]));
   DLH_X1 \accumulator_A_reg[10]  (.D(n_0_239), .G(n_0_228), .Q(
      accumulator_A[10]));
   DLH_X1 \accumulator_A_reg[9]  (.D(n_0_238), .G(n_0_228), .Q(accumulator_A[9]));
   DLH_X1 \accumulator_A_reg[8]  (.D(n_0_237), .G(n_0_228), .Q(accumulator_A[8]));
   DLH_X1 \accumulator_A_reg[7]  (.D(n_0_236), .G(n_0_228), .Q(accumulator_A[7]));
   DLH_X1 \accumulator_A_reg[6]  (.D(n_0_235), .G(n_0_228), .Q(accumulator_A[6]));
   DLH_X1 \accumulator_A_reg[5]  (.D(n_0_234), .G(n_0_228), .Q(accumulator_A[5]));
   DLH_X1 \accumulator_A_reg[4]  (.D(n_0_233), .G(n_0_228), .Q(accumulator_A[4]));
   DLH_X1 \accumulator_A_reg[3]  (.D(n_0_232), .G(n_0_228), .Q(accumulator_A[3]));
   DLH_X1 \accumulator_A_reg[2]  (.D(n_0_231), .G(n_0_228), .Q(accumulator_A[2]));
   DLH_X1 \accumulator_A_reg[1]  (.D(n_0_230), .G(n_0_228), .Q(accumulator_A[1]));
   DLH_X1 \accumulator_A_reg[0]  (.D(n_0_229), .G(n_0_228), .Q(accumulator_A[0]));
   DLH_X1 \multiplicand_Q_reg[32]  (.D(n_0_292), .G(n_0_228), .Q(n_0_190));
   DLH_X1 \multiplicand_Q_reg[31]  (.D(n_0_291), .G(n_0_228), .Q(n_0_191));
   DLH_X1 \multiplicand_Q_reg[30]  (.D(n_0_290), .G(n_0_228), .Q(n_0_192));
   DLH_X1 \multiplicand_Q_reg[29]  (.D(n_0_289), .G(n_0_228), .Q(n_0_193));
   DLH_X1 \multiplicand_Q_reg[28]  (.D(n_0_288), .G(n_0_228), .Q(n_0_194));
   DLH_X1 \multiplicand_Q_reg[27]  (.D(n_0_287), .G(n_0_228), .Q(n_0_195));
   DLH_X1 \multiplicand_Q_reg[26]  (.D(n_0_286), .G(n_0_228), .Q(n_0_196));
   DLH_X1 \multiplicand_Q_reg[25]  (.D(n_0_285), .G(n_0_228), .Q(n_0_197));
   DLH_X1 \multiplicand_Q_reg[24]  (.D(n_0_284), .G(n_0_228), .Q(n_0_198));
   DLH_X1 \multiplicand_Q_reg[23]  (.D(n_0_283), .G(n_0_228), .Q(n_0_199));
   DLH_X1 \multiplicand_Q_reg[22]  (.D(n_0_282), .G(n_0_228), .Q(n_0_200));
   DLH_X1 \multiplicand_Q_reg[21]  (.D(n_0_281), .G(n_0_228), .Q(n_0_201));
   DLH_X1 \multiplicand_Q_reg[20]  (.D(n_0_280), .G(n_0_228), .Q(n_0_202));
   DLH_X1 \multiplicand_Q_reg[19]  (.D(n_0_279), .G(n_0_228), .Q(n_0_203));
   DLH_X1 \multiplicand_Q_reg[18]  (.D(n_0_278), .G(n_0_228), .Q(n_0_204));
   DLH_X1 \multiplicand_Q_reg[17]  (.D(n_0_277), .G(n_0_228), .Q(n_0_205));
   DLH_X1 \multiplicand_Q_reg[16]  (.D(n_0_276), .G(n_0_228), .Q(n_0_206));
   DLH_X1 \multiplicand_Q_reg[15]  (.D(n_0_275), .G(n_0_228), .Q(n_0_207));
   DLH_X1 \multiplicand_Q_reg[14]  (.D(n_0_274), .G(n_0_228), .Q(n_0_208));
   DLH_X1 \multiplicand_Q_reg[13]  (.D(n_0_273), .G(n_0_228), .Q(n_0_209));
   DLH_X1 \multiplicand_Q_reg[12]  (.D(n_0_272), .G(n_0_228), .Q(n_0_210));
   DLH_X1 \multiplicand_Q_reg[11]  (.D(n_0_271), .G(n_0_228), .Q(n_0_211));
   DLH_X1 \multiplicand_Q_reg[10]  (.D(n_0_270), .G(n_0_228), .Q(n_0_212));
   DLH_X1 \multiplicand_Q_reg[9]  (.D(n_0_269), .G(n_0_228), .Q(n_0_213));
   DLH_X1 \multiplicand_Q_reg[8]  (.D(n_0_268), .G(n_0_228), .Q(n_0_214));
   DLH_X1 \multiplicand_Q_reg[7]  (.D(n_0_267), .G(n_0_228), .Q(n_0_215));
   DLH_X1 \multiplicand_Q_reg[6]  (.D(n_0_266), .G(n_0_228), .Q(n_0_216));
   DLH_X1 \multiplicand_Q_reg[5]  (.D(n_0_265), .G(n_0_228), .Q(n_0_217));
   DLH_X1 \multiplicand_Q_reg[4]  (.D(n_0_264), .G(n_0_228), .Q(n_0_218));
   DLH_X1 \multiplicand_Q_reg[3]  (.D(n_0_263), .G(n_0_228), .Q(n_0_219));
   DLH_X1 \multiplicand_Q_reg[2]  (.D(n_0_262), .G(n_0_228), .Q(n_0_220));
   DLH_X1 \multiplicand_Q_reg[1]  (.D(n_0_261), .G(n_0_228), .Q(Res[0]));
   DLH_X1 \multiplicand_Q_reg[0]  (.D(n_0_260), .G(n_0_228), .Q(n_0_0));
   DLH_X1 \multiplier_M_reg[31]  (.D(n_0_324), .G(n_0_325), .Q(multiplier_M[31]));
   DLH_X1 \multiplier_M_reg[30]  (.D(n_0_323), .G(n_0_325), .Q(multiplier_M[30]));
   DLH_X1 \multiplier_M_reg[29]  (.D(n_0_322), .G(n_0_325), .Q(multiplier_M[29]));
   DLH_X1 \multiplier_M_reg[28]  (.D(n_0_321), .G(n_0_325), .Q(multiplier_M[28]));
   DLH_X1 \multiplier_M_reg[27]  (.D(n_0_320), .G(n_0_325), .Q(multiplier_M[27]));
   DLH_X1 \multiplier_M_reg[26]  (.D(n_0_319), .G(n_0_325), .Q(multiplier_M[26]));
   DLH_X1 \multiplier_M_reg[25]  (.D(n_0_318), .G(n_0_325), .Q(multiplier_M[25]));
   DLH_X1 \multiplier_M_reg[24]  (.D(n_0_317), .G(n_0_325), .Q(multiplier_M[24]));
   DLH_X1 \multiplier_M_reg[23]  (.D(n_0_316), .G(n_0_325), .Q(multiplier_M[23]));
   DLH_X1 \multiplier_M_reg[22]  (.D(n_0_315), .G(n_0_325), .Q(multiplier_M[22]));
   DLH_X1 \multiplier_M_reg[21]  (.D(n_0_314), .G(n_0_325), .Q(multiplier_M[21]));
   DLH_X1 \multiplier_M_reg[20]  (.D(n_0_313), .G(n_0_325), .Q(multiplier_M[20]));
   DLH_X1 \multiplier_M_reg[19]  (.D(n_0_312), .G(n_0_325), .Q(multiplier_M[19]));
   DLH_X1 \multiplier_M_reg[18]  (.D(n_0_311), .G(n_0_325), .Q(multiplier_M[18]));
   DLH_X1 \multiplier_M_reg[17]  (.D(n_0_310), .G(n_0_325), .Q(multiplier_M[17]));
   DLH_X1 \multiplier_M_reg[16]  (.D(n_0_309), .G(n_0_325), .Q(multiplier_M[16]));
   DLH_X1 \multiplier_M_reg[15]  (.D(n_0_308), .G(n_0_325), .Q(multiplier_M[15]));
   DLH_X1 \multiplier_M_reg[14]  (.D(n_0_307), .G(n_0_325), .Q(multiplier_M[14]));
   DLH_X1 \multiplier_M_reg[13]  (.D(n_0_306), .G(n_0_325), .Q(multiplier_M[13]));
   DLH_X1 \multiplier_M_reg[12]  (.D(n_0_305), .G(n_0_325), .Q(multiplier_M[12]));
   DLH_X1 \multiplier_M_reg[11]  (.D(n_0_304), .G(n_0_325), .Q(multiplier_M[11]));
   DLH_X1 \multiplier_M_reg[10]  (.D(n_0_303), .G(n_0_325), .Q(multiplier_M[10]));
   DLH_X1 \multiplier_M_reg[9]  (.D(n_0_302), .G(n_0_325), .Q(multiplier_M[9]));
   DLH_X1 \multiplier_M_reg[8]  (.D(n_0_301), .G(n_0_325), .Q(multiplier_M[8]));
   DLH_X1 \multiplier_M_reg[7]  (.D(n_0_300), .G(n_0_325), .Q(multiplier_M[7]));
   DLH_X1 \multiplier_M_reg[6]  (.D(n_0_299), .G(n_0_325), .Q(multiplier_M[6]));
   DLH_X1 \multiplier_M_reg[5]  (.D(n_0_298), .G(n_0_325), .Q(multiplier_M[5]));
   DLH_X1 \multiplier_M_reg[4]  (.D(n_0_297), .G(n_0_325), .Q(multiplier_M[4]));
   DLH_X1 \multiplier_M_reg[3]  (.D(n_0_296), .G(n_0_325), .Q(multiplier_M[3]));
   DLH_X1 \multiplier_M_reg[2]  (.D(n_0_295), .G(n_0_325), .Q(multiplier_M[2]));
   DLH_X1 \multiplier_M_reg[1]  (.D(n_0_294), .G(n_0_325), .Q(multiplier_M[1]));
   DLH_X1 \multiplier_M_reg[0]  (.D(n_0_293), .G(n_0_325), .Q(multiplier_M[0]));
   DLH_X1 ready_reg (.D(n_0_221), .G(n_0_222), .Q(ready));
   DLH_X1 \counter_reg[4]  (.D(n_0_227), .G(n_0_228), .Q(counter[4]));
   DLH_X1 \counter_reg[3]  (.D(n_0_226), .G(n_0_228), .Q(counter[3]));
   DLH_X1 \counter_reg[2]  (.D(n_0_225), .G(n_0_228), .Q(counter[2]));
   DLH_X1 \counter_reg[1]  (.D(n_0_224), .G(n_0_228), .Q(counter[1]));
   DLH_X1 \counter_reg[0]  (.D(n_0_223), .G(n_0_228), .Q(counter[0]));
   OAI211_X1 i_0_2_0 (.A(n_0_2_137), .B(clk), .C1(ready), .C2(enable), .ZN(
      n_0_221));
   NAND2_X1 i_0_2_1 (.A1(n_0_2_0), .A2(n_0_2_110), .ZN(n_0_222));
   NAND4_X1 i_0_2_2 (.A1(counter[0]), .A2(n_0_2_8), .A3(n_0_2_7), .A4(n_0_2_139), 
      .ZN(n_0_2_0));
   NOR2_X1 i_0_2_3 (.A1(n_0_325), .A2(counter[0]), .ZN(n_0_223));
   NOR2_X1 i_0_2_4 (.A1(n_0_2_1), .A2(n_0_325), .ZN(n_0_224));
   XOR2_X1 i_0_2_5 (.A(counter[1]), .B(counter[0]), .Z(n_0_2_1));
   AOI21_X1 i_0_2_6 (.A(n_0_325), .B1(n_0_2_6), .B2(n_0_2_2), .ZN(n_0_225));
   OAI21_X1 i_0_2_7 (.A(counter[2]), .B1(counter[1]), .B2(counter[0]), .ZN(
      n_0_2_2));
   NOR2_X1 i_0_2_8 (.A1(n_0_2_3), .A2(n_0_325), .ZN(n_0_226));
   XOR2_X1 i_0_2_9 (.A(counter[3]), .B(n_0_2_6), .Z(n_0_2_3));
   NOR2_X1 i_0_2_10 (.A1(n_0_2_4), .A2(n_0_325), .ZN(n_0_227));
   XNOR2_X1 i_0_2_11 (.A(counter[4]), .B(n_0_2_5), .ZN(n_0_2_4));
   NOR2_X1 i_0_2_12 (.A1(n_0_2_6), .A2(counter[3]), .ZN(n_0_2_5));
   OR3_X1 i_0_2_13 (.A1(counter[2]), .A2(counter[1]), .A3(counter[0]), .ZN(
      n_0_2_6));
   NOR3_X1 i_0_2_14 (.A1(counter[3]), .A2(counter[2]), .A3(counter[1]), .ZN(
      n_0_2_7));
   OR2_X1 i_0_2_15 (.A1(n_0_325), .A2(n_0_2_8), .ZN(n_0_228));
   AOI21_X1 i_0_2_16 (.A(ready), .B1(enable), .B2(clk), .ZN(n_0_2_8));
   INV_X1 i_0_2_17 (.A(n_0_2_9), .ZN(n_0_229));
   AOI222_X1 i_0_2_18 (.A1(accumulator_A[1]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_159), .C1(n_0_2_73), .C2(n_0_127), .ZN(n_0_2_9));
   INV_X1 i_0_2_19 (.A(n_0_2_10), .ZN(n_0_230));
   AOI222_X1 i_0_2_20 (.A1(accumulator_A[2]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_160), .C1(n_0_2_73), .C2(n_0_128), .ZN(n_0_2_10));
   INV_X1 i_0_2_21 (.A(n_0_2_11), .ZN(n_0_231));
   AOI222_X1 i_0_2_22 (.A1(accumulator_A[3]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_161), .C1(n_0_2_73), .C2(n_0_129), .ZN(n_0_2_11));
   INV_X1 i_0_2_23 (.A(n_0_2_12), .ZN(n_0_232));
   AOI222_X1 i_0_2_24 (.A1(accumulator_A[4]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_162), .C1(n_0_2_73), .C2(n_0_130), .ZN(n_0_2_12));
   INV_X1 i_0_2_25 (.A(n_0_2_13), .ZN(n_0_233));
   AOI222_X1 i_0_2_26 (.A1(accumulator_A[5]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_163), .C1(n_0_2_73), .C2(n_0_131), .ZN(n_0_2_13));
   INV_X1 i_0_2_27 (.A(n_0_2_14), .ZN(n_0_234));
   AOI222_X1 i_0_2_28 (.A1(accumulator_A[6]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_164), .C1(n_0_2_73), .C2(n_0_132), .ZN(n_0_2_14));
   INV_X1 i_0_2_29 (.A(n_0_2_15), .ZN(n_0_235));
   AOI222_X1 i_0_2_30 (.A1(accumulator_A[7]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_165), .C1(n_0_2_73), .C2(n_0_133), .ZN(n_0_2_15));
   INV_X1 i_0_2_31 (.A(n_0_2_16), .ZN(n_0_236));
   AOI222_X1 i_0_2_32 (.A1(accumulator_A[8]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_166), .C1(n_0_2_73), .C2(n_0_134), .ZN(n_0_2_16));
   INV_X1 i_0_2_33 (.A(n_0_2_17), .ZN(n_0_237));
   AOI222_X1 i_0_2_34 (.A1(accumulator_A[9]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_167), .C1(n_0_2_73), .C2(n_0_135), .ZN(n_0_2_17));
   INV_X1 i_0_2_35 (.A(n_0_2_18), .ZN(n_0_238));
   AOI222_X1 i_0_2_36 (.A1(accumulator_A[10]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_168), .C1(n_0_2_73), .C2(n_0_136), .ZN(n_0_2_18));
   INV_X1 i_0_2_37 (.A(n_0_2_19), .ZN(n_0_239));
   AOI222_X1 i_0_2_38 (.A1(accumulator_A[11]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_169), .C1(n_0_2_73), .C2(n_0_137), .ZN(n_0_2_19));
   INV_X1 i_0_2_39 (.A(n_0_2_20), .ZN(n_0_240));
   AOI222_X1 i_0_2_40 (.A1(accumulator_A[12]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_170), .C1(n_0_2_73), .C2(n_0_138), .ZN(n_0_2_20));
   INV_X1 i_0_2_41 (.A(n_0_2_21), .ZN(n_0_241));
   AOI222_X1 i_0_2_42 (.A1(accumulator_A[13]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_171), .C1(n_0_2_73), .C2(n_0_139), .ZN(n_0_2_21));
   INV_X1 i_0_2_43 (.A(n_0_2_22), .ZN(n_0_242));
   AOI222_X1 i_0_2_44 (.A1(accumulator_A[14]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_172), .C1(n_0_2_73), .C2(n_0_140), .ZN(n_0_2_22));
   INV_X1 i_0_2_45 (.A(n_0_2_23), .ZN(n_0_243));
   AOI222_X1 i_0_2_46 (.A1(accumulator_A[15]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_173), .C1(n_0_2_73), .C2(n_0_141), .ZN(n_0_2_23));
   INV_X1 i_0_2_47 (.A(n_0_2_24), .ZN(n_0_244));
   AOI222_X1 i_0_2_48 (.A1(accumulator_A[16]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_174), .C1(n_0_2_73), .C2(n_0_142), .ZN(n_0_2_24));
   INV_X1 i_0_2_49 (.A(n_0_2_25), .ZN(n_0_245));
   AOI222_X1 i_0_2_50 (.A1(accumulator_A[17]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_175), .C1(n_0_2_73), .C2(n_0_143), .ZN(n_0_2_25));
   INV_X1 i_0_2_51 (.A(n_0_2_26), .ZN(n_0_246));
   AOI222_X1 i_0_2_52 (.A1(accumulator_A[18]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_176), .C1(n_0_2_73), .C2(n_0_144), .ZN(n_0_2_26));
   INV_X1 i_0_2_53 (.A(n_0_2_27), .ZN(n_0_247));
   AOI222_X1 i_0_2_54 (.A1(accumulator_A[19]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_177), .C1(n_0_2_73), .C2(n_0_145), .ZN(n_0_2_27));
   INV_X1 i_0_2_55 (.A(n_0_2_28), .ZN(n_0_248));
   AOI222_X1 i_0_2_56 (.A1(accumulator_A[20]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_178), .C1(n_0_2_73), .C2(n_0_146), .ZN(n_0_2_28));
   INV_X1 i_0_2_57 (.A(n_0_2_29), .ZN(n_0_249));
   AOI222_X1 i_0_2_58 (.A1(accumulator_A[21]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_179), .C1(n_0_2_73), .C2(n_0_147), .ZN(n_0_2_29));
   INV_X1 i_0_2_59 (.A(n_0_2_30), .ZN(n_0_250));
   AOI222_X1 i_0_2_60 (.A1(accumulator_A[22]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_180), .C1(n_0_2_73), .C2(n_0_148), .ZN(n_0_2_30));
   INV_X1 i_0_2_61 (.A(n_0_2_31), .ZN(n_0_251));
   AOI222_X1 i_0_2_62 (.A1(accumulator_A[23]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_181), .C1(n_0_2_73), .C2(n_0_149), .ZN(n_0_2_31));
   INV_X1 i_0_2_63 (.A(n_0_2_32), .ZN(n_0_252));
   AOI222_X1 i_0_2_64 (.A1(accumulator_A[24]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_182), .C1(n_0_2_73), .C2(n_0_150), .ZN(n_0_2_32));
   INV_X1 i_0_2_65 (.A(n_0_2_33), .ZN(n_0_253));
   AOI222_X1 i_0_2_66 (.A1(accumulator_A[25]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_183), .C1(n_0_2_73), .C2(n_0_151), .ZN(n_0_2_33));
   INV_X1 i_0_2_67 (.A(n_0_2_34), .ZN(n_0_254));
   AOI222_X1 i_0_2_68 (.A1(accumulator_A[26]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_184), .C1(n_0_2_73), .C2(n_0_152), .ZN(n_0_2_34));
   INV_X1 i_0_2_69 (.A(n_0_2_35), .ZN(n_0_255));
   AOI222_X1 i_0_2_70 (.A1(accumulator_A[27]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_185), .C1(n_0_2_73), .C2(n_0_153), .ZN(n_0_2_35));
   INV_X1 i_0_2_71 (.A(n_0_2_36), .ZN(n_0_256));
   AOI222_X1 i_0_2_72 (.A1(accumulator_A[28]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_186), .C1(n_0_2_73), .C2(n_0_154), .ZN(n_0_2_36));
   INV_X1 i_0_2_73 (.A(n_0_2_37), .ZN(n_0_257));
   AOI222_X1 i_0_2_74 (.A1(accumulator_A[29]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_187), .C1(n_0_2_73), .C2(n_0_155), .ZN(n_0_2_37));
   INV_X1 i_0_2_75 (.A(n_0_2_38), .ZN(n_0_258));
   AOI222_X1 i_0_2_76 (.A1(accumulator_A[30]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_188), .C1(n_0_2_73), .C2(n_0_156), .ZN(n_0_2_38));
   INV_X1 i_0_2_77 (.A(n_0_2_39), .ZN(n_0_259));
   AOI222_X1 i_0_2_78 (.A1(accumulator_A[30]), .A2(n_0_2_76), .B1(n_0_2_75), 
      .B2(n_0_189), .C1(n_0_2_73), .C2(n_0_157), .ZN(n_0_2_39));
   AND2_X1 i_0_2_79 (.A1(n_0_2_137), .A2(n_0_2_40), .ZN(n_0_261));
   MUX2_X1 i_0_2_80 (.A(B[0]), .B(n_0_220), .S(n_0_2_111), .Z(n_0_2_40));
   INV_X1 i_0_2_81 (.A(n_0_2_41), .ZN(n_0_262));
   AOI222_X1 i_0_2_82 (.A1(n_0_219), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_1), 
      .C1(n_0_2_71), .C2(B[1]), .ZN(n_0_2_41));
   INV_X1 i_0_2_83 (.A(n_0_2_42), .ZN(n_0_263));
   AOI222_X1 i_0_2_84 (.A1(n_0_218), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_2), 
      .C1(n_0_2_71), .C2(B[2]), .ZN(n_0_2_42));
   INV_X1 i_0_2_85 (.A(n_0_2_43), .ZN(n_0_264));
   AOI222_X1 i_0_2_86 (.A1(n_0_217), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_3), 
      .C1(n_0_2_71), .C2(B[3]), .ZN(n_0_2_43));
   INV_X1 i_0_2_87 (.A(n_0_2_44), .ZN(n_0_265));
   AOI222_X1 i_0_2_88 (.A1(n_0_216), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_4), 
      .C1(n_0_2_71), .C2(B[4]), .ZN(n_0_2_44));
   INV_X1 i_0_2_89 (.A(n_0_2_45), .ZN(n_0_266));
   AOI222_X1 i_0_2_90 (.A1(n_0_215), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_5), 
      .C1(n_0_2_71), .C2(B[5]), .ZN(n_0_2_45));
   INV_X1 i_0_2_91 (.A(n_0_2_46), .ZN(n_0_267));
   AOI222_X1 i_0_2_92 (.A1(n_0_214), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_6), 
      .C1(n_0_2_71), .C2(B[6]), .ZN(n_0_2_46));
   INV_X1 i_0_2_93 (.A(n_0_2_47), .ZN(n_0_268));
   AOI222_X1 i_0_2_94 (.A1(n_0_213), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_7), 
      .C1(n_0_2_71), .C2(B[7]), .ZN(n_0_2_47));
   INV_X1 i_0_2_95 (.A(n_0_2_48), .ZN(n_0_269));
   AOI222_X1 i_0_2_96 (.A1(n_0_212), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_8), 
      .C1(n_0_2_71), .C2(B[8]), .ZN(n_0_2_48));
   INV_X1 i_0_2_97 (.A(n_0_2_49), .ZN(n_0_270));
   AOI222_X1 i_0_2_98 (.A1(n_0_211), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_9), 
      .C1(n_0_2_71), .C2(B[9]), .ZN(n_0_2_49));
   INV_X1 i_0_2_99 (.A(n_0_2_50), .ZN(n_0_271));
   AOI222_X1 i_0_2_100 (.A1(n_0_210), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_10), 
      .C1(n_0_2_71), .C2(B[10]), .ZN(n_0_2_50));
   INV_X1 i_0_2_101 (.A(n_0_2_51), .ZN(n_0_272));
   AOI222_X1 i_0_2_102 (.A1(n_0_209), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_11), 
      .C1(n_0_2_71), .C2(B[11]), .ZN(n_0_2_51));
   INV_X1 i_0_2_103 (.A(n_0_2_52), .ZN(n_0_273));
   AOI222_X1 i_0_2_104 (.A1(n_0_208), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_12), 
      .C1(n_0_2_71), .C2(B[12]), .ZN(n_0_2_52));
   INV_X1 i_0_2_105 (.A(n_0_2_53), .ZN(n_0_274));
   AOI222_X1 i_0_2_106 (.A1(n_0_207), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_13), 
      .C1(n_0_2_71), .C2(B[13]), .ZN(n_0_2_53));
   INV_X1 i_0_2_107 (.A(n_0_2_54), .ZN(n_0_275));
   AOI222_X1 i_0_2_108 (.A1(n_0_206), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_14), 
      .C1(n_0_2_71), .C2(B[14]), .ZN(n_0_2_54));
   INV_X1 i_0_2_109 (.A(n_0_2_55), .ZN(n_0_276));
   AOI222_X1 i_0_2_110 (.A1(n_0_205), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_15), 
      .C1(n_0_2_71), .C2(B[15]), .ZN(n_0_2_55));
   INV_X1 i_0_2_111 (.A(n_0_2_56), .ZN(n_0_277));
   AOI222_X1 i_0_2_112 (.A1(n_0_204), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_16), 
      .C1(n_0_2_71), .C2(B[16]), .ZN(n_0_2_56));
   INV_X1 i_0_2_113 (.A(n_0_2_57), .ZN(n_0_278));
   AOI222_X1 i_0_2_114 (.A1(n_0_203), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_17), 
      .C1(n_0_2_71), .C2(B[17]), .ZN(n_0_2_57));
   INV_X1 i_0_2_115 (.A(n_0_2_58), .ZN(n_0_279));
   AOI222_X1 i_0_2_116 (.A1(n_0_202), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_18), 
      .C1(n_0_2_71), .C2(B[18]), .ZN(n_0_2_58));
   INV_X1 i_0_2_117 (.A(n_0_2_59), .ZN(n_0_280));
   AOI222_X1 i_0_2_118 (.A1(n_0_201), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_19), 
      .C1(n_0_2_71), .C2(B[19]), .ZN(n_0_2_59));
   INV_X1 i_0_2_119 (.A(n_0_2_60), .ZN(n_0_281));
   AOI222_X1 i_0_2_120 (.A1(n_0_200), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_20), 
      .C1(n_0_2_71), .C2(B[20]), .ZN(n_0_2_60));
   INV_X1 i_0_2_121 (.A(n_0_2_61), .ZN(n_0_282));
   AOI222_X1 i_0_2_122 (.A1(n_0_199), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_21), 
      .C1(n_0_2_71), .C2(B[21]), .ZN(n_0_2_61));
   INV_X1 i_0_2_123 (.A(n_0_2_62), .ZN(n_0_283));
   AOI222_X1 i_0_2_124 (.A1(n_0_198), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_22), 
      .C1(n_0_2_71), .C2(B[22]), .ZN(n_0_2_62));
   INV_X1 i_0_2_125 (.A(n_0_2_63), .ZN(n_0_284));
   AOI222_X1 i_0_2_126 (.A1(n_0_197), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_23), 
      .C1(n_0_2_71), .C2(B[23]), .ZN(n_0_2_63));
   INV_X1 i_0_2_127 (.A(n_0_2_64), .ZN(n_0_285));
   AOI222_X1 i_0_2_128 (.A1(n_0_196), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_24), 
      .C1(n_0_2_71), .C2(B[24]), .ZN(n_0_2_64));
   INV_X1 i_0_2_129 (.A(n_0_2_65), .ZN(n_0_286));
   AOI222_X1 i_0_2_130 (.A1(n_0_195), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_25), 
      .C1(n_0_2_71), .C2(B[25]), .ZN(n_0_2_65));
   INV_X1 i_0_2_131 (.A(n_0_2_66), .ZN(n_0_287));
   AOI222_X1 i_0_2_132 (.A1(n_0_194), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_26), 
      .C1(n_0_2_71), .C2(B[26]), .ZN(n_0_2_66));
   INV_X1 i_0_2_133 (.A(n_0_2_67), .ZN(n_0_288));
   AOI222_X1 i_0_2_134 (.A1(n_0_193), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_27), 
      .C1(n_0_2_71), .C2(B[27]), .ZN(n_0_2_67));
   INV_X1 i_0_2_135 (.A(n_0_2_68), .ZN(n_0_289));
   AOI222_X1 i_0_2_136 (.A1(n_0_192), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_28), 
      .C1(n_0_2_71), .C2(B[28]), .ZN(n_0_2_68));
   INV_X1 i_0_2_137 (.A(n_0_2_69), .ZN(n_0_290));
   AOI222_X1 i_0_2_138 (.A1(n_0_191), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_29), 
      .C1(n_0_2_71), .C2(B[29]), .ZN(n_0_2_69));
   INV_X1 i_0_2_139 (.A(n_0_2_70), .ZN(n_0_291));
   AOI222_X1 i_0_2_140 (.A1(n_0_190), .A2(n_0_2_110), .B1(n_0_2_78), .B2(n_0_30), 
      .C1(n_0_2_71), .C2(B[30]), .ZN(n_0_2_70));
   NOR3_X1 i_0_2_141 (.A1(n_0_2_111), .A2(reset), .A3(B[31]), .ZN(n_0_2_71));
   NAND2_X1 i_0_2_142 (.A1(n_0_2_72), .A2(n_0_2_74), .ZN(n_0_292));
   AOI222_X1 i_0_2_143 (.A1(accumulator_A[0]), .A2(n_0_2_76), .B1(n_0_2_73), 
      .B2(n_0_126), .C1(n_0_31), .C2(n_0_2_78), .ZN(n_0_2_72));
   NOR3_X1 i_0_2_144 (.A1(n_0_325), .A2(Res[0]), .A3(n_0_2_140), .ZN(n_0_2_73));
   NAND2_X1 i_0_2_145 (.A1(n_0_158), .A2(n_0_2_75), .ZN(n_0_2_74));
   AND2_X1 i_0_2_146 (.A1(n_0_260), .A2(n_0_2_140), .ZN(n_0_2_75));
   AND2_X1 i_0_2_147 (.A1(Res[0]), .A2(n_0_2_110), .ZN(n_0_260));
   NOR2_X1 i_0_2_148 (.A1(n_0_325), .A2(n_0_2_77), .ZN(n_0_2_76));
   XNOR2_X1 i_0_2_149 (.A(Res[0]), .B(n_0_2_140), .ZN(n_0_2_77));
   NOR3_X1 i_0_2_150 (.A1(n_0_2_138), .A2(n_0_2_111), .A3(reset), .ZN(n_0_2_78));
   AND2_X1 i_0_2_151 (.A1(n_0_2_137), .A2(A[0]), .ZN(n_0_293));
   INV_X1 i_0_2_152 (.A(n_0_2_79), .ZN(n_0_294));
   AOI22_X1 i_0_2_153 (.A1(n_0_32), .A2(n_0_327), .B1(n_0_2_109), .B2(A[1]), 
      .ZN(n_0_2_79));
   INV_X1 i_0_2_154 (.A(n_0_2_80), .ZN(n_0_295));
   AOI22_X1 i_0_2_155 (.A1(n_0_33), .A2(n_0_327), .B1(n_0_2_109), .B2(A[2]), 
      .ZN(n_0_2_80));
   INV_X1 i_0_2_156 (.A(n_0_2_81), .ZN(n_0_296));
   AOI22_X1 i_0_2_157 (.A1(n_0_34), .A2(n_0_327), .B1(n_0_2_109), .B2(A[3]), 
      .ZN(n_0_2_81));
   INV_X1 i_0_2_158 (.A(n_0_2_82), .ZN(n_0_297));
   AOI22_X1 i_0_2_159 (.A1(n_0_35), .A2(n_0_327), .B1(n_0_2_109), .B2(A[4]), 
      .ZN(n_0_2_82));
   INV_X1 i_0_2_160 (.A(n_0_2_83), .ZN(n_0_298));
   AOI22_X1 i_0_2_161 (.A1(n_0_36), .A2(n_0_327), .B1(n_0_2_109), .B2(A[5]), 
      .ZN(n_0_2_83));
   INV_X1 i_0_2_162 (.A(n_0_2_84), .ZN(n_0_299));
   AOI22_X1 i_0_2_163 (.A1(n_0_37), .A2(n_0_327), .B1(n_0_2_109), .B2(A[6]), 
      .ZN(n_0_2_84));
   INV_X1 i_0_2_164 (.A(n_0_2_85), .ZN(n_0_300));
   AOI22_X1 i_0_2_165 (.A1(n_0_38), .A2(n_0_327), .B1(n_0_2_109), .B2(A[7]), 
      .ZN(n_0_2_85));
   INV_X1 i_0_2_166 (.A(n_0_2_86), .ZN(n_0_301));
   AOI22_X1 i_0_2_167 (.A1(n_0_39), .A2(n_0_327), .B1(n_0_2_109), .B2(A[8]), 
      .ZN(n_0_2_86));
   INV_X1 i_0_2_168 (.A(n_0_2_87), .ZN(n_0_302));
   AOI22_X1 i_0_2_169 (.A1(n_0_40), .A2(n_0_327), .B1(n_0_2_109), .B2(A[9]), 
      .ZN(n_0_2_87));
   INV_X1 i_0_2_170 (.A(n_0_2_88), .ZN(n_0_303));
   AOI22_X1 i_0_2_171 (.A1(n_0_41), .A2(n_0_327), .B1(n_0_2_109), .B2(A[10]), 
      .ZN(n_0_2_88));
   INV_X1 i_0_2_172 (.A(n_0_2_89), .ZN(n_0_304));
   AOI22_X1 i_0_2_173 (.A1(n_0_42), .A2(n_0_327), .B1(n_0_2_109), .B2(A[11]), 
      .ZN(n_0_2_89));
   INV_X1 i_0_2_174 (.A(n_0_2_90), .ZN(n_0_305));
   AOI22_X1 i_0_2_175 (.A1(n_0_43), .A2(n_0_327), .B1(n_0_2_109), .B2(A[12]), 
      .ZN(n_0_2_90));
   INV_X1 i_0_2_176 (.A(n_0_2_91), .ZN(n_0_306));
   AOI22_X1 i_0_2_177 (.A1(n_0_44), .A2(n_0_327), .B1(n_0_2_109), .B2(A[13]), 
      .ZN(n_0_2_91));
   INV_X1 i_0_2_178 (.A(n_0_2_92), .ZN(n_0_307));
   AOI22_X1 i_0_2_179 (.A1(n_0_45), .A2(n_0_327), .B1(n_0_2_109), .B2(A[14]), 
      .ZN(n_0_2_92));
   INV_X1 i_0_2_180 (.A(n_0_2_93), .ZN(n_0_308));
   AOI22_X1 i_0_2_181 (.A1(n_0_46), .A2(n_0_327), .B1(n_0_2_109), .B2(A[15]), 
      .ZN(n_0_2_93));
   INV_X1 i_0_2_182 (.A(n_0_2_94), .ZN(n_0_309));
   AOI22_X1 i_0_2_183 (.A1(n_0_47), .A2(n_0_327), .B1(n_0_2_109), .B2(A[16]), 
      .ZN(n_0_2_94));
   INV_X1 i_0_2_184 (.A(n_0_2_95), .ZN(n_0_310));
   AOI22_X1 i_0_2_185 (.A1(n_0_48), .A2(n_0_327), .B1(n_0_2_109), .B2(A[17]), 
      .ZN(n_0_2_95));
   INV_X1 i_0_2_186 (.A(n_0_2_96), .ZN(n_0_311));
   AOI22_X1 i_0_2_187 (.A1(n_0_49), .A2(n_0_327), .B1(n_0_2_109), .B2(A[18]), 
      .ZN(n_0_2_96));
   INV_X1 i_0_2_188 (.A(n_0_2_97), .ZN(n_0_312));
   AOI22_X1 i_0_2_189 (.A1(n_0_50), .A2(n_0_327), .B1(n_0_2_109), .B2(A[19]), 
      .ZN(n_0_2_97));
   INV_X1 i_0_2_190 (.A(n_0_2_98), .ZN(n_0_313));
   AOI22_X1 i_0_2_191 (.A1(n_0_51), .A2(n_0_327), .B1(n_0_2_109), .B2(A[20]), 
      .ZN(n_0_2_98));
   INV_X1 i_0_2_192 (.A(n_0_2_99), .ZN(n_0_314));
   AOI22_X1 i_0_2_193 (.A1(n_0_52), .A2(n_0_327), .B1(n_0_2_109), .B2(A[21]), 
      .ZN(n_0_2_99));
   INV_X1 i_0_2_194 (.A(n_0_2_100), .ZN(n_0_315));
   AOI22_X1 i_0_2_195 (.A1(n_0_53), .A2(n_0_327), .B1(n_0_2_109), .B2(A[22]), 
      .ZN(n_0_2_100));
   INV_X1 i_0_2_196 (.A(n_0_2_101), .ZN(n_0_316));
   AOI22_X1 i_0_2_197 (.A1(n_0_54), .A2(n_0_327), .B1(n_0_2_109), .B2(A[23]), 
      .ZN(n_0_2_101));
   INV_X1 i_0_2_198 (.A(n_0_2_102), .ZN(n_0_317));
   AOI22_X1 i_0_2_199 (.A1(n_0_55), .A2(n_0_327), .B1(n_0_2_109), .B2(A[24]), 
      .ZN(n_0_2_102));
   INV_X1 i_0_2_200 (.A(n_0_2_103), .ZN(n_0_318));
   AOI22_X1 i_0_2_201 (.A1(n_0_56), .A2(n_0_327), .B1(n_0_2_109), .B2(A[25]), 
      .ZN(n_0_2_103));
   INV_X1 i_0_2_202 (.A(n_0_2_104), .ZN(n_0_319));
   AOI22_X1 i_0_2_203 (.A1(n_0_57), .A2(n_0_327), .B1(n_0_2_109), .B2(A[26]), 
      .ZN(n_0_2_104));
   INV_X1 i_0_2_204 (.A(n_0_2_105), .ZN(n_0_320));
   AOI22_X1 i_0_2_205 (.A1(n_0_58), .A2(n_0_327), .B1(n_0_2_109), .B2(A[27]), 
      .ZN(n_0_2_105));
   INV_X1 i_0_2_206 (.A(n_0_2_106), .ZN(n_0_321));
   AOI22_X1 i_0_2_207 (.A1(n_0_59), .A2(n_0_327), .B1(n_0_2_109), .B2(A[28]), 
      .ZN(n_0_2_106));
   INV_X1 i_0_2_208 (.A(n_0_2_107), .ZN(n_0_322));
   AOI22_X1 i_0_2_209 (.A1(n_0_60), .A2(n_0_327), .B1(n_0_2_109), .B2(A[29]), 
      .ZN(n_0_2_107));
   INV_X1 i_0_2_210 (.A(n_0_2_108), .ZN(n_0_323));
   AOI22_X1 i_0_2_211 (.A1(n_0_61), .A2(n_0_327), .B1(n_0_2_109), .B2(A[30]), 
      .ZN(n_0_2_108));
   NOR2_X1 i_0_2_212 (.A1(A[31]), .A2(reset), .ZN(n_0_2_109));
   AND2_X1 i_0_2_213 (.A1(n_0_62), .A2(n_0_327), .ZN(n_0_324));
   INV_X1 i_0_2_214 (.A(n_0_2_110), .ZN(n_0_325));
   AND2_X1 i_0_2_215 (.A1(n_0_2_137), .A2(n_0_2_111), .ZN(n_0_2_110));
   NAND3_X1 i_0_2_216 (.A1(clk), .A2(ready), .A3(enable), .ZN(n_0_2_111));
   NOR2_X1 i_0_2_217 (.A1(n_0_2_138), .A2(reset), .ZN(n_0_326));
   AND2_X1 i_0_2_218 (.A1(n_0_2_137), .A2(A[31]), .ZN(n_0_327));
   AOI21_X1 i_0_2_219 (.A(n_0_2_112), .B1(n_0_2_113), .B2(n_0_125), .ZN(OVF));
   AOI21_X1 i_0_2_220 (.A(isNeg[0]), .B1(n_0_2_114), .B2(accumulator_A[30]), 
      .ZN(n_0_2_112));
   MUX2_X1 i_0_2_221 (.A(n_0_63), .B(n_0_220), .S(n_0_2_114), .Z(Res[1]));
   MUX2_X1 i_0_2_222 (.A(n_0_64), .B(n_0_219), .S(n_0_2_114), .Z(Res[2]));
   MUX2_X1 i_0_2_223 (.A(n_0_65), .B(n_0_218), .S(n_0_2_114), .Z(Res[3]));
   MUX2_X1 i_0_2_224 (.A(n_0_66), .B(n_0_217), .S(n_0_2_114), .Z(Res[4]));
   MUX2_X1 i_0_2_225 (.A(n_0_67), .B(n_0_216), .S(n_0_2_114), .Z(Res[5]));
   MUX2_X1 i_0_2_226 (.A(n_0_68), .B(n_0_215), .S(n_0_2_114), .Z(Res[6]));
   MUX2_X1 i_0_2_227 (.A(n_0_69), .B(n_0_214), .S(n_0_2_114), .Z(Res[7]));
   MUX2_X1 i_0_2_228 (.A(n_0_70), .B(n_0_213), .S(n_0_2_114), .Z(Res[8]));
   MUX2_X1 i_0_2_229 (.A(n_0_71), .B(n_0_212), .S(n_0_2_114), .Z(Res[9]));
   MUX2_X1 i_0_2_230 (.A(n_0_72), .B(n_0_211), .S(n_0_2_114), .Z(Res[10]));
   MUX2_X1 i_0_2_231 (.A(n_0_73), .B(n_0_210), .S(n_0_2_114), .Z(Res[11]));
   MUX2_X1 i_0_2_232 (.A(n_0_74), .B(n_0_209), .S(n_0_2_114), .Z(Res[12]));
   MUX2_X1 i_0_2_233 (.A(n_0_75), .B(n_0_208), .S(n_0_2_114), .Z(Res[13]));
   MUX2_X1 i_0_2_234 (.A(n_0_76), .B(n_0_207), .S(n_0_2_114), .Z(Res[14]));
   MUX2_X1 i_0_2_235 (.A(n_0_77), .B(n_0_206), .S(n_0_2_114), .Z(Res[15]));
   MUX2_X1 i_0_2_236 (.A(n_0_78), .B(n_0_205), .S(n_0_2_114), .Z(Res[16]));
   MUX2_X1 i_0_2_237 (.A(n_0_79), .B(n_0_204), .S(n_0_2_114), .Z(Res[17]));
   MUX2_X1 i_0_2_238 (.A(n_0_80), .B(n_0_203), .S(n_0_2_114), .Z(Res[18]));
   MUX2_X1 i_0_2_239 (.A(n_0_81), .B(n_0_202), .S(n_0_2_114), .Z(Res[19]));
   MUX2_X1 i_0_2_240 (.A(n_0_82), .B(n_0_201), .S(n_0_2_114), .Z(Res[20]));
   MUX2_X1 i_0_2_241 (.A(n_0_83), .B(n_0_200), .S(n_0_2_114), .Z(Res[21]));
   MUX2_X1 i_0_2_242 (.A(n_0_84), .B(n_0_199), .S(n_0_2_114), .Z(Res[22]));
   MUX2_X1 i_0_2_243 (.A(n_0_85), .B(n_0_198), .S(n_0_2_114), .Z(Res[23]));
   MUX2_X1 i_0_2_244 (.A(n_0_86), .B(n_0_197), .S(n_0_2_114), .Z(Res[24]));
   MUX2_X1 i_0_2_245 (.A(n_0_87), .B(n_0_196), .S(n_0_2_114), .Z(Res[25]));
   MUX2_X1 i_0_2_246 (.A(n_0_88), .B(n_0_195), .S(n_0_2_114), .Z(Res[26]));
   MUX2_X1 i_0_2_247 (.A(n_0_89), .B(n_0_194), .S(n_0_2_114), .Z(Res[27]));
   MUX2_X1 i_0_2_248 (.A(n_0_90), .B(n_0_193), .S(n_0_2_114), .Z(Res[28]));
   MUX2_X1 i_0_2_249 (.A(n_0_91), .B(n_0_192), .S(n_0_2_114), .Z(Res[29]));
   MUX2_X1 i_0_2_250 (.A(n_0_92), .B(n_0_191), .S(n_0_2_114), .Z(Res[30]));
   MUX2_X1 i_0_2_251 (.A(n_0_93), .B(n_0_190), .S(n_0_2_114), .Z(Res[31]));
   MUX2_X1 i_0_2_252 (.A(n_0_94), .B(accumulator_A[0]), .S(n_0_2_114), .Z(
      Res[32]));
   MUX2_X1 i_0_2_253 (.A(n_0_95), .B(accumulator_A[1]), .S(n_0_2_114), .Z(
      Res[33]));
   MUX2_X1 i_0_2_254 (.A(n_0_96), .B(accumulator_A[2]), .S(n_0_2_114), .Z(
      Res[34]));
   MUX2_X1 i_0_2_255 (.A(n_0_97), .B(accumulator_A[3]), .S(n_0_2_114), .Z(
      Res[35]));
   MUX2_X1 i_0_2_256 (.A(n_0_98), .B(accumulator_A[4]), .S(n_0_2_114), .Z(
      Res[36]));
   MUX2_X1 i_0_2_257 (.A(n_0_99), .B(accumulator_A[5]), .S(n_0_2_114), .Z(
      Res[37]));
   MUX2_X1 i_0_2_258 (.A(n_0_100), .B(accumulator_A[6]), .S(n_0_2_114), .Z(
      Res[38]));
   MUX2_X1 i_0_2_259 (.A(n_0_101), .B(accumulator_A[7]), .S(n_0_2_114), .Z(
      Res[39]));
   MUX2_X1 i_0_2_260 (.A(n_0_102), .B(accumulator_A[8]), .S(n_0_2_114), .Z(
      Res[40]));
   MUX2_X1 i_0_2_261 (.A(n_0_103), .B(accumulator_A[9]), .S(n_0_2_114), .Z(
      Res[41]));
   MUX2_X1 i_0_2_262 (.A(n_0_104), .B(accumulator_A[10]), .S(n_0_2_114), 
      .Z(Res[42]));
   MUX2_X1 i_0_2_263 (.A(n_0_105), .B(accumulator_A[11]), .S(n_0_2_114), 
      .Z(Res[43]));
   MUX2_X1 i_0_2_264 (.A(n_0_106), .B(accumulator_A[12]), .S(n_0_2_114), 
      .Z(Res[44]));
   MUX2_X1 i_0_2_265 (.A(n_0_107), .B(accumulator_A[13]), .S(n_0_2_114), 
      .Z(Res[45]));
   MUX2_X1 i_0_2_266 (.A(n_0_108), .B(accumulator_A[14]), .S(n_0_2_114), 
      .Z(Res[46]));
   MUX2_X1 i_0_2_267 (.A(n_0_109), .B(accumulator_A[15]), .S(n_0_2_114), 
      .Z(Res[47]));
   MUX2_X1 i_0_2_268 (.A(n_0_110), .B(accumulator_A[16]), .S(n_0_2_114), 
      .Z(Res[48]));
   MUX2_X1 i_0_2_269 (.A(n_0_111), .B(accumulator_A[17]), .S(n_0_2_114), 
      .Z(Res[49]));
   MUX2_X1 i_0_2_270 (.A(n_0_112), .B(accumulator_A[18]), .S(n_0_2_114), 
      .Z(Res[50]));
   MUX2_X1 i_0_2_271 (.A(n_0_113), .B(accumulator_A[19]), .S(n_0_2_114), 
      .Z(Res[51]));
   MUX2_X1 i_0_2_272 (.A(n_0_114), .B(accumulator_A[20]), .S(n_0_2_114), 
      .Z(Res[52]));
   MUX2_X1 i_0_2_273 (.A(n_0_115), .B(accumulator_A[21]), .S(n_0_2_114), 
      .Z(Res[53]));
   MUX2_X1 i_0_2_274 (.A(n_0_116), .B(accumulator_A[22]), .S(n_0_2_114), 
      .Z(Res[54]));
   MUX2_X1 i_0_2_275 (.A(n_0_117), .B(accumulator_A[23]), .S(n_0_2_114), 
      .Z(Res[55]));
   MUX2_X1 i_0_2_276 (.A(n_0_118), .B(accumulator_A[24]), .S(n_0_2_114), 
      .Z(Res[56]));
   MUX2_X1 i_0_2_277 (.A(n_0_119), .B(accumulator_A[25]), .S(n_0_2_114), 
      .Z(Res[57]));
   MUX2_X1 i_0_2_278 (.A(n_0_120), .B(accumulator_A[26]), .S(n_0_2_114), 
      .Z(Res[58]));
   MUX2_X1 i_0_2_279 (.A(n_0_121), .B(accumulator_A[27]), .S(n_0_2_114), 
      .Z(Res[59]));
   MUX2_X1 i_0_2_280 (.A(n_0_122), .B(accumulator_A[28]), .S(n_0_2_114), 
      .Z(Res[60]));
   MUX2_X1 i_0_2_281 (.A(n_0_123), .B(accumulator_A[29]), .S(n_0_2_114), 
      .Z(Res[61]));
   MUX2_X1 i_0_2_282 (.A(n_0_124), .B(accumulator_A[30]), .S(n_0_2_114), 
      .Z(Res[62]));
   MUX2_X1 i_0_2_283 (.A(n_0_125), .B(accumulator_A[30]), .S(n_0_2_114), 
      .Z(Res[63]));
   INV_X1 i_0_2_284 (.A(n_0_2_114), .ZN(n_0_2_113));
   NAND2_X1 i_0_2_285 (.A1(n_0_2_116), .A2(n_0_2_115), .ZN(n_0_2_114));
   XOR2_X1 i_0_2_286 (.A(isNeg[1]), .B(isNeg[0]), .Z(n_0_2_115));
   OR4_X1 i_0_2_287 (.A1(n_0_2_132), .A2(n_0_2_127), .A3(n_0_2_122), .A4(
      n_0_2_117), .ZN(n_0_2_116));
   NAND4_X1 i_0_2_288 (.A1(n_0_2_121), .A2(n_0_2_120), .A3(n_0_2_119), .A4(
      n_0_2_118), .ZN(n_0_2_117));
   NOR4_X1 i_0_2_289 (.A1(accumulator_A[15]), .A2(accumulator_A[11]), .A3(
      accumulator_A[10]), .A4(accumulator_A[9]), .ZN(n_0_2_118));
   NOR4_X1 i_0_2_290 (.A1(accumulator_A[14]), .A2(accumulator_A[13]), .A3(
      accumulator_A[12]), .A4(accumulator_A[8]), .ZN(n_0_2_119));
   NOR4_X1 i_0_2_291 (.A1(accumulator_A[3]), .A2(accumulator_A[2]), .A3(
      accumulator_A[1]), .A4(accumulator_A[0]), .ZN(n_0_2_120));
   NOR4_X1 i_0_2_292 (.A1(accumulator_A[7]), .A2(accumulator_A[6]), .A3(
      accumulator_A[5]), .A4(accumulator_A[4]), .ZN(n_0_2_121));
   NAND4_X1 i_0_2_293 (.A1(n_0_2_126), .A2(n_0_2_125), .A3(n_0_2_124), .A4(
      n_0_2_123), .ZN(n_0_2_122));
   NOR4_X1 i_0_2_294 (.A1(accumulator_A[27]), .A2(accumulator_A[26]), .A3(
      accumulator_A[25]), .A4(accumulator_A[16]), .ZN(n_0_2_123));
   NOR4_X1 i_0_2_295 (.A1(accumulator_A[30]), .A2(accumulator_A[29]), .A3(
      accumulator_A[28]), .A4(accumulator_A[24]), .ZN(n_0_2_124));
   NOR4_X1 i_0_2_296 (.A1(accumulator_A[19]), .A2(accumulator_A[18]), .A3(
      accumulator_A[17]), .A4(Res[0]), .ZN(n_0_2_125));
   NOR4_X1 i_0_2_297 (.A1(accumulator_A[23]), .A2(accumulator_A[22]), .A3(
      accumulator_A[21]), .A4(accumulator_A[20]), .ZN(n_0_2_126));
   NAND4_X1 i_0_2_298 (.A1(n_0_2_131), .A2(n_0_2_130), .A3(n_0_2_129), .A4(
      n_0_2_128), .ZN(n_0_2_127));
   NOR3_X1 i_0_2_299 (.A1(n_0_202), .A2(n_0_203), .A3(n_0_204), .ZN(n_0_2_128));
   NOR4_X1 i_0_2_300 (.A1(n_0_198), .A2(n_0_199), .A3(n_0_200), .A4(n_0_201), 
      .ZN(n_0_2_129));
   NOR4_X1 i_0_2_301 (.A1(n_0_194), .A2(n_0_195), .A3(n_0_196), .A4(n_0_205), 
      .ZN(n_0_2_130));
   NOR4_X1 i_0_2_302 (.A1(n_0_191), .A2(n_0_192), .A3(n_0_193), .A4(n_0_197), 
      .ZN(n_0_2_131));
   NAND4_X1 i_0_2_303 (.A1(n_0_2_136), .A2(n_0_2_135), .A3(n_0_2_134), .A4(
      n_0_2_133), .ZN(n_0_2_132));
   NOR4_X1 i_0_2_304 (.A1(n_0_206), .A2(n_0_210), .A3(n_0_211), .A4(n_0_212), 
      .ZN(n_0_2_133));
   NOR4_X1 i_0_2_305 (.A1(n_0_207), .A2(n_0_208), .A3(n_0_209), .A4(n_0_213), 
      .ZN(n_0_2_134));
   NOR4_X1 i_0_2_306 (.A1(n_0_190), .A2(n_0_218), .A3(n_0_219), .A4(n_0_220), 
      .ZN(n_0_2_135));
   NOR4_X1 i_0_2_307 (.A1(n_0_214), .A2(n_0_215), .A3(n_0_216), .A4(n_0_217), 
      .ZN(n_0_2_136));
   INV_X1 i_0_2_308 (.A(reset), .ZN(n_0_2_137));
   INV_X1 i_0_2_309 (.A(B[31]), .ZN(n_0_2_138));
   INV_X1 i_0_2_310 (.A(counter[4]), .ZN(n_0_2_139));
   INV_X1 i_0_2_311 (.A(n_0_0), .ZN(n_0_2_140));
endmodule
