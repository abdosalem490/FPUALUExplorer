* SPICE NETLIST
***************************************

.SUBCKT MGC_via1_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT WELLTAP
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT FILLCELL_X2
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_2
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2_X1 A2 VSS A1 ZN VDD 6
** N=7 EP=6 IP=0 FDC=4
M0 7 A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN A1 7 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=2 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via1_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=2 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X4
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT via1_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT via2_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2_X1 A1 A2 VSS VDD ZN
** N=7 EP=5 IP=0 FDC=6
M0 6 A1 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 A1 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XNOR2_X1 VSS A ZN B VDD 6
** N=10 EP=6 IP=0 FDC=10
M0 10 A 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=155 $Y=90 $D=1
M1 VSS B 10 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=345 $Y=90 $D=1
M2 8 7 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=540 $Y=90 $D=1
M3 ZN A 8 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 8 B ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 7 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=155 $Y=995 $D=0
M6 VDD B 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=345 $Y=995 $D=0
M7 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=540 $Y=680 $D=0
M8 9 A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M9 VDD B 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI221_X1 B2 B1 VSS A C2 VDD C1 ZN 9
** N=13 EP=9 IP=0 FDC=10
M0 VSS B2 10 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 10 B1 VSS 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 11 A 10 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN C2 11 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 11 C1 ZN 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 12 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 ZN B1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 13 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 ZN C1 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV_X1 A VSS VDD ZN 5
** N=5 EP=5 IP=0 FDC=2
M0 ZN A VSS 5 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4
** N=4 EP=4 IP=8 FDC=2
X1 3 1 2 4 1 INV_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT NAND4_X1 A4 VSS A3 A2 A1 ZN VDD
** N=10 EP=7 IP=0 FDC=8
M0 8 A4 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 9 A3 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 10 A2 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN A4 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 VDD A3 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 ZN A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 VDD A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI22_X1 B2 B1 VSS ZN A1 A2 VDD 8
** N=11 EP=8 IP=0 FDC=8
M0 VSS B2 9 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 9 B1 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A1 9 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 9 A2 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 10 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 ZN B1 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 11 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 VDD A2 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT XOR2_X1 VDD A Z B VSS 6
** N=10 EP=6 IP=0 FDC=10
M0 7 A VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 7 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 10 A Z 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 10 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 9 A 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 8 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 8 B Z VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FILLCELL_X8
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_13
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4 5 6 7
** N=7 EP=7 IP=11 FDC=8
X1 3 4 1 5 6 7 2 1 OAI22_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_20
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4 5 6 7
** N=7 EP=7 IP=11 FDC=8
X1 3 4 1 5 6 7 2 1 OAI22_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT OAI21_X1 B2 B1 ZN A VSS VDD 7
** N=9 EP=7 IP=0 FDC=6
M0 ZN B2 8 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 8 B1 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS A 8 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=550 $Y=90 $D=1
M3 9 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M4 ZN B1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M5 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=550 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=6
X1 3 5 4 6 1 2 7 OAI21_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_23
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT AOI21_X1 B2 B1 ZN A VSS VDD
** N=8 EP=6 IP=0 FDC=6
M0 8 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN B1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M4 7 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M5 VDD A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR2_X1 A2 VDD A1 ZN VSS 6
** N=7 EP=6 IP=0 FDC=4
M0 ZN A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A1 ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 7 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 ZN A1 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_25
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT OR4_X1 A1 A2 A3 A4 VSS VDD ZN
** N=11 EP=7 IP=0 FDC=10
M0 8 A1 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 8 A3 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 VSS A4 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=715 $Y=90 $D=1
M4 ZN 8 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 9 A1 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 10 A2 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 11 A3 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M8 VDD A4 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=715 $Y=995 $D=0
M9 ZN 8 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=13 FDC=10
X0 1 2 3 4 2 INV_X1 $T=950 0 0 0 $X=835 $Y=-115
X1 5 6 2 7 8 9 3 2 OAI22_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=13 FDC=10
X0 1 2 3 4 2 INV_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 5 6 2 7 8 9 3 2 OAI22_X1 $T=380 0 0 0 $X=265 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_28
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_29
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_30
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_31
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=16 FDC=16
X0 1 2 3 4 5 6 7 3 OAI22_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 8 9 3 10 11 12 7 3 OAI22_X1 $T=950 0 0 0 $X=835 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_33
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FA_X1 CO CI B A VDD VSS S
** N=19 EP=7 IP=0 FDC=28
M0 VSS 8 CO VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 17 B VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06 $X=360 $Y=215 $D=1
M2 8 A 17 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=550 $Y=215 $D=1
M3 9 CI 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07 $X=740 $Y=215 $D=1
M4 VSS A 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07 $X=935 $Y=215 $D=1
M5 9 B VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1125 $Y=215 $D=1
M6 11 B VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1465 $Y=90 $D=1
M7 VSS CI 11 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1655 $Y=90 $D=1
M8 11 A VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1845 $Y=90 $D=1
M9 13 8 11 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07 $X=2035 $Y=90 $D=1
M10 18 CI 13 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.15e-14 PD=7e-07 PS=7.2e-07 $X=2235 $Y=90 $D=1
M11 19 B 18 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2425 $Y=90 $D=1
M12 VSS A 19 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=2615 $Y=90 $D=1
M13 S 13 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=2805 $Y=90 $D=1
M14 VDD 8 CO VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M15 14 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.54e-06 $X=360 $Y=870 $D=0
M16 8 A 14 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=550 $Y=870 $D=0
M17 10 CI 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06 PS=9.1e-07 $X=740 $Y=870 $D=0
M18 VDD A 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.53e-14 PD=9.1e-07 PS=1.07e-06 $X=935 $Y=945 $D=0
M19 10 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1125 $Y=945 $D=0
M20 12 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1465 $Y=995 $D=0
M21 VDD CI 12 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1655 $Y=995 $D=0
M22 12 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1845 $Y=995 $D=0
M23 13 8 12 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07 $X=2035 $Y=995 $D=0
M24 15 CI 13 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.725e-14 PD=9.1e-07 PS=9.3e-07 $X=2235 $Y=995 $D=0
M25 16 B 15 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=2425 $Y=995 $D=0
M26 VDD A 16 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2615 $Y=995 $D=0
M27 S 13 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2805 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI22_X1 B2 B1 VDD A1 ZN A2 VSS 8
** N=11 EP=8 IP=0 FDC=8
M0 10 B2 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN B1 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 11 A1 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 VSS A2 11 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 VDD B2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 9 B1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 ZN A1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 9 A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_34
** N=3 EP=0 IP=3 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_35
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_36
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_37
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT HA_X1 S B A VSS VDD CO
** N=12 EP=6 IP=0 FDC=16
M0 11 B VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 S A 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS 8 S VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.48e-14 AS=5.81e-14 PD=1.12e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 8 B VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.48e-14 PD=7e-07 PS=1.12e-06 $X=760 $Y=90 $D=1
M4 VSS A 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=950 $Y=90 $D=1
M5 12 A 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1320 $Y=90 $D=1
M6 VSS B 12 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=1510 $Y=90 $D=1
M7 CO 9 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1700 $Y=90 $D=1
M8 S B 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M9 7 A S VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M10 VDD 8 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.7725e-14 AS=8.82e-14 PD=1.55e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M11 10 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.7725e-14 PD=9.1e-07 PS=1.55e-06 $X=760 $Y=870 $D=0
M12 8 A 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=950 $Y=870 $D=0
M13 9 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1320 $Y=870 $D=0
M14 VDD B 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=1510 $Y=870 $D=0
M15 CO 9 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1700 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR2_X2 A1 ZN A2 VSS VDD
** N=7 EP=5 IP=0 FDC=8
M0 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 6 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN A1 6 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 7 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 VDD A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_38
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_39
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_40
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_41 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=2
X1 3 1 2 4 5 INV_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT NAND3_X1 A3 VSS A2 A1 VDD ZN
** N=8 EP=6 IP=0 FDC=6
M0 7 A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 8 A2 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 VDD A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_42
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X16
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT OAI33_X1 B3 B2 B1 VSS A1 A2 A3 ZN VDD
** N=14 EP=9 IP=0 FDC=12
M0 10 B3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS B2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 10 B1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 ZN A1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 10 A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 ZN A3 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1110 $Y=90 $D=1
M6 11 B3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M7 12 B2 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M8 ZN B1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M9 13 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M10 14 A2 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
M11 VDD A3 14 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1110 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_43
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_44
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_45
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_46
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT OAI222_X1 C2 C1 VSS B1 B2 A2 VDD A1 ZN
** N=14 EP=9 IP=0 FDC=12
M0 10 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=155 $Y=90 $D=1
M1 VSS C1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=345 $Y=90 $D=1
M2 10 B1 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=710 $Y=90 $D=1
M3 11 B2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=900 $Y=90 $D=1
M4 ZN A2 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1090 $Y=90 $D=1
M5 11 A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1280 $Y=90 $D=1
M6 12 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=155 $Y=680 $D=0
M7 ZN C1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=1.9845e-13 AS=8.82e-14 PD=1.89e-06 PS=1.54e-06 $X=345 $Y=680 $D=0
M8 13 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.9845e-13 PD=1.54e-06 PS=1.89e-06 $X=710 $Y=680 $D=0
M9 VDD B2 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=900 $Y=680 $D=0
M10 14 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1090 $Y=680 $D=0
M11 ZN A1 14 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1280 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI21_X2 A VDD B1 ZN B2 VSS
** N=9 EP=6 IP=0 FDC=12
M0 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 8 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 9 B1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=945 $Y=90 $D=1
M5 VSS B2 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1135 $Y=90 $D=1
M6 VDD A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M7 7 A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M8 ZN B2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M9 7 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
M10 ZN B1 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=945 $Y=680 $D=0
M11 7 B2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1135 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_47 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=4
X0 1 2 3 4 2 INV_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 5 2 3 6 2 INV_X1 $T=380 0 0 0 $X=265 $Y=-115
.ENDS
***************************************
.SUBCKT FILLCELL_X32
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_48 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=10
X0 1 2 3 5 6 7 8 4 9 OAI221_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT NOR3_X1 A3 VDD A2 A1 VSS ZN
** N=8 EP=6 IP=0 FDC=6
M0 ZN A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 8 A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI211_X1 C2 C1 A VDD B ZN VSS
** N=10 EP=7 IP=0 FDC=8
M0 ZN C2 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 8 C1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 10 A 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS B 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 9 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN C1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 ZN B VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AND2_X1 A1 A2 VSS VDD ZN
** N=7 EP=5 IP=0 FDC=6
M0 7 A1 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 6 A1 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OR3_X1 A1 A2 A3 VSS VDD ZN
** N=9 EP=6 IP=0 FDC=8
M0 VSS A1 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 7 A2 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 VSS A3 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=525 $Y=90 $D=1
M3 ZN 7 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 8 A1 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M5 9 A2 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M6 VDD A3 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=525 $Y=995 $D=0
M7 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_49 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=18
X0 1 2 3 4 5 6 7 11 OAI22_X1 $T=1140 0 0 0 $X=1025 $Y=-115
X1 7 8 9 10 3 11 XOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT CLKBUF_X2 A Z VSS VDD
** N=5 EP=4 IP=0 FDC=6
M0 VSS A 5 VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07 $X=145 $Y=90 $D=1
M1 Z 5 VSS VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=335 $Y=90 $D=1
M2 VSS 5 Z VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=525 $Y=90 $D=1
M3 VDD A 5 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 Z 5 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 VDD 5 Z VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI221_X1 B2 B1 VDD A C2 VSS C1 ZN
** N=12 EP=8 IP=0 FDC=10
M0 11 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN B1 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 12 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN C1 12 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 VDD B2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 9 B1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 10 A 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 ZN C2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 10 C1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FPU_VA B[31] B[24] A[25] SUM[20] A[27] A[23] B[28] B[30] SUM[9] A[30] A[20] B[3] SUM[19] SUM[15] B[27] SUM[2] A[28] B[17] B[11] A[14]
+ A[18] A[17] B[6] B[4] A[31] B[21] B[19] B[8] A[8] A[19] A[15] B[0] B[7] B[5] SUM[31] B[26] SUM[22] B[29] SUM[0] SUM[4]
+ B[23] SUM[29] SUM[8] SUM[10] SUM[30] A[26] SUM[5] B[16] B[14] A[12] A[11] B[18] B[13] A[22] B[2] A[10] B[1] A[9] A[21] B[22]
+ B[20] A[7] A[5] A[3] A[0] B[25] A[29] SUM[27] SUM[1] SUM[24] SUM[7] A[24] A[16] B[10] B[9] A[4] SUM[21] A[1] SUM[18] SUM[17]
+ A[6] A[2] B[15] SUM[16] SUM[26] SUM[25] SUM[23] SUM[28] SUM[12] SUM[11] B[12] SUM[14] A[13] SUM[6] SUM[13] SUM[3]
** N=996 EP=96 IP=14688 FDC=6266
M0 78 97 325 78 NMOS_VTL L=5e-08 W=9.5e-08 AD=2.03e-14 AS=9.975e-15 PD=6.7e-07 PS=4e-07 $X=15415 $Y=43160 $D=1
M1 33 325 78 78 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.03e-14 PD=6e-07 PS=6.7e-07 $X=15605 $Y=43160 $D=1
M2 78 5 327 78 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07 $X=16535 $Y=42700 $D=1
M3 97 327 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=16725 $Y=42495 $D=1
M4 989 167 332 78 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=27555 $Y=6300 $D=1
M5 990 180 989 78 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=27745 $Y=6300 $D=1
M6 991 266 990 78 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=27935 $Y=6300 $D=1
M7 78 211 991 78 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=28125 $Y=6300 $D=1
M8 333 332 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=28315 $Y=6095 $D=1
M9 992 334 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=28735 $Y=9490 $D=1
M10 339 182 992 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=28925 $Y=9490 $D=1
M11 78 187 339 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=29115 $Y=9490 $D=1
M12 339 338 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=29305 $Y=9490 $D=1
M13 993 347 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=34585 $Y=40290 $D=1
M14 351 245 993 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=1.2035e-13 AS=5.81e-14 PD=1.41e-06 PS=1.11e-06 $X=34775 $Y=40290 $D=1
M15 994 B[28] 351 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=1.2035e-13 PD=1.11e-06 PS=1.41e-06 $X=35115 $Y=40290 $D=1
M16 78 249 994 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=35305 $Y=40290 $D=1
M17 995 217 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=35495 $Y=40290 $D=1
M18 351 B[27] 995 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=35685 $Y=40290 $D=1
M19 78 270 357 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=37245 $Y=43090 $D=1
M20 357 270 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37435 $Y=43090 $D=1
M21 78 270 357 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37625 $Y=43090 $D=1
M22 357 270 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37815 $Y=43090 $D=1
M23 5 360 357 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38005 $Y=43090 $D=1
M24 357 B[30] 5 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38195 $Y=43090 $D=1
M25 5 B[30] 357 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38385 $Y=43090 $D=1
M26 357 360 5 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38575 $Y=43090 $D=1
M27 5 360 357 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38765 $Y=43090 $D=1
M28 357 B[30] 5 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38955 $Y=43090 $D=1
M29 5 B[30] 357 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=39145 $Y=43090 $D=1
M30 357 360 5 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=39335 $Y=43090 $D=1
M31 1 364 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=42565 $Y=39695 $D=1
M32 78 364 1 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=42755 $Y=39695 $D=1
M33 1 364 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=42945 $Y=39695 $D=1
M34 78 364 1 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43135 $Y=39695 $D=1
M35 1 369 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43325 $Y=39695 $D=1
M36 78 369 1 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43515 $Y=39695 $D=1
M37 1 369 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43705 $Y=39695 $D=1
M38 78 369 1 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=43895 $Y=39695 $D=1
M39 1 371 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=44270 $Y=39695 $D=1
M40 78 371 1 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=44460 $Y=39695 $D=1
M41 1 371 78 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=44650 $Y=39695 $D=1
M42 78 371 1 78 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=44840 $Y=39695 $D=1
M43 310 97 325 310 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=15415 $Y=43995 $D=0
M44 33 325 310 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=15605 $Y=43680 $D=0
M45 310 5 327 310 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=16535 $Y=41690 $D=0
M46 97 327 310 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=16725 $Y=41690 $D=0
M47 332 167 310 310 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=27555 $Y=5290 $D=0
M48 310 180 332 310 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=27745 $Y=5290 $D=0
M49 332 266 310 310 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=27935 $Y=5290 $D=0
M50 310 211 332 310 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=28125 $Y=5290 $D=0
M51 333 332 310 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=28315 $Y=5290 $D=0
M52 339 334 337 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=28735 $Y=10080 $D=0
M53 337 182 339 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=28925 $Y=10080 $D=0
M54 984 187 337 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=29115 $Y=10080 $D=0
M55 310 338 984 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=29305 $Y=10080 $D=0
M56 349 347 310 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=34585 $Y=40880 $D=0
M57 310 245 349 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=34775 $Y=40880 $D=0
M58 349 B[28] 352 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=35115 $Y=40880 $D=0
M59 352 249 349 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=35305 $Y=40880 $D=0
M60 351 217 352 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=35495 $Y=40880 $D=0
M61 352 B[27] 351 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=35685 $Y=40880 $D=0
M62 5 270 310 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=37245 $Y=43680 $D=0
M63 310 270 5 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37435 $Y=43680 $D=0
M64 5 270 310 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37625 $Y=43680 $D=0
M65 310 270 5 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37815 $Y=43680 $D=0
M66 985 360 310 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38005 $Y=43680 $D=0
M67 5 B[30] 985 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38195 $Y=43680 $D=0
M68 986 B[30] 5 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38385 $Y=43680 $D=0
M69 310 360 986 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38575 $Y=43680 $D=0
M70 987 360 310 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38765 $Y=43680 $D=0
M71 5 B[30] 987 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38955 $Y=43680 $D=0
M72 988 B[30] 5 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=39145 $Y=43680 $D=0
M73 310 360 988 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=39335 $Y=43680 $D=0
M74 1 364 370 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=42565 $Y=38890 $D=0
M75 370 364 1 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=42755 $Y=38890 $D=0
M76 1 364 370 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=42945 $Y=38890 $D=0
M77 370 364 1 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43135 $Y=38890 $D=0
M78 372 369 370 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43325 $Y=38890 $D=0
M79 370 369 372 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43515 $Y=38890 $D=0
M80 372 369 370 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43705 $Y=38890 $D=0
M81 370 369 372 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=43895 $Y=38890 $D=0
M82 372 371 310 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=44270 $Y=38890 $D=0
M83 310 371 372 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=44460 $Y=38890 $D=0
M84 372 371 310 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=44650 $Y=38890 $D=0
M85 310 371 372 310 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=44840 $Y=38890 $D=0
X5002 400 78 9 670 310 78 NAND2_X1 $T=1380 20600 0 0 $X=1265 $Y=20485
X5003 897 78 8 671 310 78 NAND2_X1 $T=2330 15000 1 0 $X=2215 $Y=13485
X5004 853 78 30 691 310 78 NAND2_X1 $T=5180 6600 0 0 $X=5065 $Y=6485
X5005 428 78 50 901 310 78 NAND2_X1 $T=7650 26200 1 0 $X=7535 $Y=24685
X5006 57 78 36 404 310 78 NAND2_X1 $T=8030 31800 1 0 $X=7915 $Y=30285
X5007 440 78 32 476 310 78 NAND2_X1 $T=12780 31800 1 0 $X=12665 $Y=30285
X5008 91 78 77 19 310 78 NAND2_X1 $T=13730 40200 0 0 $X=13615 $Y=40085
X5009 736 78 72 475 310 996 NAND2_X1 $T=14110 1000 0 0 $X=13995 $Y=885
X5010 506 78 136 937 310 78 NAND2_X1 $T=19810 9400 1 0 $X=19695 $Y=7885
X5011 507 78 122 505 310 78 NAND2_X1 $T=20000 6600 1 0 $X=19885 $Y=5085
X5012 329 78 134 758 310 78 NAND2_X1 $T=21140 15000 1 0 $X=21025 $Y=13485
X5013 211 78 253 549 310 78 NAND2_X1 $T=26650 9400 1 0 $X=26535 $Y=7885
X5014 266 78 220 776 310 78 NAND2_X1 $T=26650 12200 1 0 $X=26535 $Y=10685
X5015 180 78 780 171 310 78 NAND2_X1 $T=27980 12200 0 0 $X=27865 $Y=12085
X5016 242 78 297 200 310 78 NAND2_X1 $T=29500 15000 1 0 $X=29385 $Y=13485
X5017 570 78 583 275 310 78 NAND2_X1 $T=31970 20600 1 0 $X=31855 $Y=19085
X5018 229 78 797 955 310 78 NAND2_X1 $T=32920 26200 0 0 $X=32805 $Y=26085
X5019 218 78 225 348 310 78 NAND2_X1 $T=33110 9400 1 0 $X=32995 $Y=7885
X5020 607 78 275 233 310 78 NAND2_X1 $T=34440 15000 1 0 $X=34325 $Y=13485
X5021 260 78 793 811 310 78 NAND2_X1 $T=35770 23400 1 0 $X=35655 $Y=21885
X5022 256 78 250 361 310 78 NAND2_X1 $T=36910 20600 1 0 $X=36795 $Y=19085
X5023 603 78 618 SUM[27] 310 78 NAND2_X1 $T=37100 29000 0 0 $X=36985 $Y=28885
X5024 271 78 618 SUM[26] 310 78 NAND2_X1 $T=37480 31800 0 0 $X=37365 $Y=31685
X5025 272 78 618 SUM[25] 310 78 NAND2_X1 $T=37480 34600 1 0 $X=37365 $Y=33085
X5026 273 78 618 SUM[24] 310 78 NAND2_X1 $T=38810 31800 1 0 $X=38695 $Y=30285
X5027 225 78 265 630 310 78 NAND2_X1 $T=39950 9400 1 0 $X=39835 $Y=7885
X5028 225 78 250 615 310 78 NAND2_X1 $T=40330 6600 0 0 $X=40215 $Y=6485
X5029 296 78 618 SUM[23] 310 78 NAND2_X1 $T=40520 26200 0 0 $X=40405 $Y=26085
X5030 225 78 254 648 310 78 NAND2_X1 $T=41280 6600 0 0 $X=41165 $Y=6485
X5031 225 78 237 649 310 78 NAND2_X1 $T=42420 9400 1 0 $X=42305 $Y=7885
X5032 293 78 618 SUM[28] 310 78 NAND2_X1 $T=42420 26200 0 0 $X=42305 $Y=26085
X5033 295 78 618 SUM[29] 310 78 NAND2_X1 $T=42610 31800 1 0 $X=42495 $Y=30285
X5034 618 78 368 SUM[30] 310 78 NAND2_X1 $T=42990 29000 0 0 $X=42875 $Y=28885
X5035 A[30] 78 B[30] 663 310 78 NAND2_X1 $T=44510 43000 0 0 $X=44395 $Y=42885
X7347 670 4 78 310 678 OR2_X1 $T=2330 20600 1 0 $X=2215 $Y=19085
X7348 671 6 78 310 844 OR2_X1 $T=2520 12200 0 0 $X=2405 $Y=12085
X7349 691 15 78 310 414 OR2_X1 $T=4990 6600 1 0 $X=4875 $Y=5085
X7350 678 28 78 310 40 OR2_X1 $T=5750 20600 1 0 $X=5635 $Y=19085
X7351 901 31 78 310 311 OR2_X1 $T=5940 23400 0 0 $X=5825 $Y=23285
X7352 460 67 78 310 459 OR2_X1 $T=12590 34600 0 0 $X=12475 $Y=34485
X7353 88 90 78 310 86 OR2_X1 $T=15250 29000 1 0 $X=15135 $Y=27485
X7354 475 92 78 310 468 OR2_X1 $T=15440 3800 1 0 $X=15325 $Y=2285
X7355 399 93 78 310 485 OR2_X1 $T=15440 9400 0 0 $X=15325 $Y=9285
X7356 516 107 78 310 74 OR2_X1 $T=18100 20600 0 0 $X=17985 $Y=20485
X7357 912 116 78 310 106 OR2_X1 $T=19430 31800 0 0 $X=19315 $Y=31685
X7358 505 118 78 310 512 OR2_X1 $T=20380 3800 1 0 $X=20265 $Y=2285
X7359 509 123 78 310 912 OR2_X1 $T=20760 34600 1 0 $X=20645 $Y=33085
X7360 512 127 78 310 142 OR2_X1 $T=21140 3800 1 0 $X=21025 $Y=2285
X7361 772 146 78 310 124 OR2_X1 $T=24180 20600 1 0 $X=24065 $Y=19085
X7362 554 147 78 310 129 OR2_X1 $T=24180 23400 0 0 $X=24065 $Y=23285
X7363 SUM[31] 148 78 310 547 OR2_X1 $T=24370 15000 1 0 $X=24255 $Y=13485
X7364 173 154 78 310 541 OR2_X1 $T=24940 17800 1 0 $X=24825 $Y=16285
X7365 165 158 78 310 166 OR2_X1 $T=25510 15000 0 0 $X=25395 $Y=14885
X7366 557 169 78 310 554 OR2_X1 $T=27220 26200 0 0 $X=27105 $Y=26085
X7367 781 174 78 310 161 OR2_X1 $T=27790 23400 1 0 $X=27675 $Y=21885
X7368 336 184 78 310 781 OR2_X1 $T=28930 23400 0 0 $X=28815 $Y=23285
X7369 577 206 78 310 924 OR2_X1 $T=31020 20600 0 0 $X=30905 $Y=20485
X7370 275 218 78 310 231 OR2_X1 $T=32730 15000 1 0 $X=32615 $Y=13485
X7371 874 244 78 310 238 OR2_X1 $T=34630 23400 0 0 $X=34515 $Y=23285
X7372 250 269 78 310 622 OR2_X1 $T=37480 20600 1 0 $X=37365 $Y=19085
X7373 250 278 78 310 825 OR2_X1 $T=39000 17800 0 0 $X=38885 $Y=17685
X7374 366 282 78 310 285 OR2_X1 $T=39380 26200 1 0 $X=39265 $Y=24685
X7375 811 285 78 310 340 OR2_X1 $T=40140 26200 1 0 $X=40025 $Y=24685
X7376 B[30] A[30] 78 310 307 OR2_X1 $T=43940 37400 0 0 $X=43825 $Y=37285
X7377 78 395 682 7 310 78 XNOR2_X1 $T=3470 6600 1 180 $X=2215 $Y=6485
X7378 78 668 398 8 310 78 XNOR2_X1 $T=3470 15000 1 180 $X=2215 $Y=14885
X7379 78 899 685 9 310 78 XNOR2_X1 $T=3470 20600 1 180 $X=2215 $Y=20485
X7380 78 681 680 10 310 78 XNOR2_X1 $T=3470 26200 0 180 $X=2215 $Y=24685
X7381 78 410 702 22 310 996 XNOR2_X1 $T=5180 1000 0 0 $X=5065 $Y=885
X7382 78 466 717 30 310 78 XNOR2_X1 $T=5750 9400 1 0 $X=5635 $Y=7885
X7383 78 710 435 50 310 78 XNOR2_X1 $T=8220 26200 1 0 $X=8105 $Y=24685
X7384 78 455 463 69 310 78 XNOR2_X1 $T=12590 9400 0 0 $X=12475 $Y=9285
X7385 78 449 456 72 310 996 XNOR2_X1 $T=12970 1000 0 0 $X=12855 $Y=885
X7386 78 754 938 122 310 78 XNOR2_X1 $T=20570 6600 1 0 $X=20455 $Y=5085
X7387 78 525 940 134 310 78 XNOR2_X1 $T=22280 15000 1 0 $X=22165 $Y=13485
X7388 78 526 531 136 310 78 XNOR2_X1 $T=22470 9400 1 0 $X=22355 $Y=7885
X7389 78 752 769 138 310 78 XNOR2_X1 $T=22850 9400 0 0 $X=22735 $Y=9285
X7390 78 148 154 767 310 78 XNOR2_X1 $T=23800 12200 0 0 $X=23685 $Y=12085
X7391 78 SUM[31] 158 162 310 78 XNOR2_X1 $T=25700 15000 1 0 $X=25585 $Y=13485
X7392 78 141 555 172 310 996 XNOR2_X1 $T=27410 1000 0 0 $X=27295 $Y=885
X7393 78 633 302 287 310 78 XNOR2_X1 $T=39950 34600 0 0 $X=39835 $Y=34485
X7394 78 307 964 302 310 78 XNOR2_X1 $T=43560 34600 0 0 $X=43445 $Y=34485
X7395 78 837 953 307 310 78 XNOR2_X1 $T=43940 34600 1 0 $X=43825 $Y=33085
X7396 78 B[6] 78 3 5 310 A[6] 17 78 OAI221_X1 $T=1950 37400 1 0 $X=1835 $Y=35885
X7397 2 63 78 1 11 310 52 387 78 OAI221_X1 $T=2330 29000 1 0 $X=2215 $Y=27485
X7398 393 52 78 1 11 310 63 402 78 OAI221_X1 $T=2330 29000 0 0 $X=2215 $Y=28885
X7399 393 63 78 1 12 310 52 679 78 OAI221_X1 $T=3470 29000 0 0 $X=3355 $Y=28885
X7400 78 B[2] 78 3 5 310 A[2] 21 78 OAI221_X1 $T=3660 43000 0 0 $X=3545 $Y=42885
X7401 407 63 78 1 13 310 52 694 78 OAI221_X1 $T=4230 26200 0 0 $X=4115 $Y=26085
X7402 313 48 78 17 19 310 38 697 78 OAI221_X1 $T=4800 37400 0 0 $X=4685 $Y=37285
X7403 19 405 78 20 24 310 48 66 78 OAI221_X1 $T=4990 40200 1 0 $X=4875 $Y=38685
X7404 705 48 78 21 19 310 666 417 78 OAI221_X1 $T=4990 43000 1 0 $X=4875 $Y=41485
X7405 312 48 78 25 19 310 852 700 78 OAI221_X1 $T=5180 40200 0 0 $X=5065 $Y=40085
X7406 407 52 78 1 29 310 63 420 78 OAI221_X1 $T=5370 26200 0 0 $X=5255 $Y=26085
X7407 78 B[1] 78 3 33 310 A[1] 854 78 OAI221_X1 $T=5750 43000 0 0 $X=5635 $Y=42885
X7408 902 52 78 1 12 310 63 314 78 OAI221_X1 $T=6320 29000 1 0 $X=6205 $Y=27485
X7409 422 63 78 1 29 310 52 855 78 OAI221_X1 $T=6890 26200 0 0 $X=6775 $Y=26085
X7410 902 63 78 1 44 310 52 432 78 OAI221_X1 $T=7460 29000 1 0 $X=7345 $Y=27485
X7411 715 52 78 1 44 310 63 439 78 OAI221_X1 $T=9550 29000 1 0 $X=9435 $Y=27485
X7412 908 448 78 32 66 310 18 95 78 OAI221_X1 $T=12020 40200 1 0 $X=11905 $Y=38685
X7413 715 63 78 1 76 310 52 471 78 OAI221_X1 $T=13160 29000 1 0 $X=13045 $Y=27485
X7414 323 52 78 1 76 310 63 481 78 OAI221_X1 $T=14300 29000 0 0 $X=14185 $Y=28885
X7415 323 63 78 1 89 310 52 483 78 OAI221_X1 $T=14680 31800 1 0 $X=14565 $Y=30285
X7416 78 B[0] 78 3 33 310 A[0] 453 78 OAI221_X1 $T=15060 43000 1 0 $X=14945 $Y=41485
X7417 89 63 78 1 96 310 52 499 78 OAI221_X1 $T=15440 31800 0 0 $X=15325 $Y=31685
X7418 78 B[3] 78 3 97 310 A[3] 68 78 OAI221_X1 $T=15820 43000 0 0 $X=15705 $Y=42885
X7419 5 498 78 3 78 310 864 484 78 OAI221_X1 $T=17150 37400 1 0 $X=17035 $Y=35885
X7420 110 52 78 1 112 310 63 500 78 OAI221_X1 $T=18290 37400 1 0 $X=18175 $Y=35885
X7421 862 63 78 1 112 310 52 501 78 OAI221_X1 $T=18480 34600 1 0 $X=18365 $Y=33085
X7422 742 52 78 1 115 310 63 503 78 OAI221_X1 $T=18670 40200 1 0 $X=18555 $Y=38685
X7423 110 63 78 1 115 310 52 504 78 OAI221_X1 $T=18860 37400 0 0 $X=18745 $Y=37285
X7424 222 B[25] 78 195 198 310 B[26] 203 78 OAI221_X1 $T=29690 40200 0 0 $X=29575 $Y=40085
X7425 A[26] 216 78 203 A[27] 310 209 880 78 OAI221_X1 $T=30450 43000 1 0 $X=30335 $Y=41485
X7426 552 B[24] 78 219 222 310 B[25] 223 78 OAI221_X1 $T=32540 37400 0 0 $X=32425 $Y=37285
X7427 A[26] 216 78 223 A[25] 310 794 245 78 OAI221_X1 $T=32730 40200 1 0 $X=32615 $Y=38685
X7428 803 229 78 224 226 310 280 791 78 OAI221_X1 $T=32920 3800 1 0 $X=32805 $Y=2285
X7429 923 265 78 228 230 310 237 236 78 OAI221_X1 $T=33300 6600 1 0 $X=33185 $Y=5085
X7430 232 280 78 224 262 310 229 342 996 OAI221_X1 $T=36150 1000 0 0 $X=36035 $Y=885
X7431 817 229 78 224 262 310 280 619 996 OAI221_X1 $T=37290 1000 0 0 $X=37175 $Y=885
X7432 817 280 78 224 283 310 229 627 996 OAI221_X1 $T=39190 1000 0 0 $X=39075 $Y=885
X7433 298 229 78 224 283 310 280 832 996 OAI221_X1 $T=40330 1000 0 0 $X=40215 $Y=885
X7434 929 229 78 224 298 310 280 656 996 OAI221_X1 $T=42800 1000 0 0 $X=42685 $Y=885
X7435 308 280 78 224 300 310 229 841 78 OAI221_X1 $T=44700 3800 1 180 $X=43445 $Y=3685
X7436 365 229 78 224 300 310 280 572 78 OAI221_X1 $T=43560 6600 0 0 $X=43445 $Y=6485
X7437 365 280 78 224 304 310 229 830 78 OAI221_X1 $T=43560 9400 0 0 $X=43445 $Y=9285
X7438 304 280 78 224 301 310 229 657 78 OAI221_X1 $T=44700 12200 1 180 $X=43445 $Y=12085
X7439 301 280 78 224 305 310 229 643 78 OAI221_X1 $T=43560 15000 1 0 $X=43445 $Y=13485
X7440 929 280 78 224 308 310 229 343 996 OAI221_X1 $T=43940 1000 0 0 $X=43825 $Y=885
X7441 831 229 78 224 305 310 280 367 78 OAI221_X1 $T=43940 15000 0 0 $X=43825 $Y=14885
X7470 896 78 310 6 78 INV_X1 $T=2140 12200 0 0 $X=2025 $Y=12085
X7471 673 78 310 4 78 INV_X1 $T=2140 17800 0 0 $X=2025 $Y=17685
X7472 387 78 310 899 78 INV_X1 $T=2140 23400 1 0 $X=2025 $Y=21885
X7473 389 78 310 395 78 INV_X1 $T=2330 6600 1 0 $X=2215 $Y=5085
X7474 390 78 310 668 78 INV_X1 $T=2330 17800 1 0 $X=2215 $Y=16285
X7475 675 78 310 15 78 INV_X1 $T=2520 3800 0 0 $X=2405 $Y=3685
X7476 677 78 310 410 996 INV_X1 $T=2900 1000 0 0 $X=2785 $Y=885
X7477 385 78 310 396 78 INV_X1 $T=2900 17800 0 0 $X=2785 $Y=17685
X7478 847 78 310 397 78 INV_X1 $T=3090 9400 1 0 $X=2975 $Y=7885
X7479 679 78 310 381 78 INV_X1 $T=3470 23400 1 180 $X=2975 $Y=23285
X7480 899 78 310 400 78 INV_X1 $T=3850 20600 1 180 $X=3355 $Y=20485
X7481 680 78 310 684 78 INV_X1 $T=3470 23400 0 0 $X=3355 $Y=23285
X7482 402 78 310 681 78 INV_X1 $T=3850 26200 0 180 $X=3355 $Y=24685
X7483 685 78 310 693 78 INV_X1 $T=3850 20600 0 0 $X=3735 $Y=20485
X7484 408 78 310 849 78 INV_X1 $T=4610 12200 1 0 $X=4495 $Y=10685
X7485 692 78 310 850 78 INV_X1 $T=4990 12200 0 0 $X=4875 $Y=12085
X7486 411 78 310 695 78 INV_X1 $T=5180 17800 1 0 $X=5065 $Y=16285
X7487 413 78 310 973 78 INV_X1 $T=5370 9400 1 0 $X=5255 $Y=7885
X7488 694 78 310 28 78 INV_X1 $T=5370 17800 0 0 $X=5255 $Y=17685
X7489 314 78 310 31 78 INV_X1 $T=6130 26200 1 0 $X=6015 $Y=24685
X7490 903 78 310 315 78 INV_X1 $T=6510 34600 1 0 $X=6395 $Y=33085
X7491 423 78 310 930 78 INV_X1 $T=7080 6600 1 0 $X=6965 $Y=5085
X7492 855 78 310 43 78 INV_X1 $T=7460 23400 1 0 $X=7345 $Y=21885
X7493 401 78 310 907 78 INV_X1 $T=7650 15000 0 0 $X=7535 $Y=14885
X7494 433 78 310 59 78 INV_X1 $T=8410 17800 1 0 $X=8295 $Y=16285
X7495 710 78 310 428 78 INV_X1 $T=8410 23400 0 0 $X=8295 $Y=23285
X7496 711 78 310 852 78 INV_X1 $T=8410 29000 0 0 $X=8295 $Y=28885
X7497 57 78 310 35 78 INV_X1 $T=8600 31800 0 0 $X=8485 $Y=31685
X7498 55 78 310 932 78 INV_X1 $T=9550 23400 1 0 $X=9435 $Y=21885
X7499 A[21] 78 310 960 78 INV_X1 $T=10120 17800 0 0 $X=10005 $Y=17685
X7500 B[21] 78 310 436 78 INV_X1 $T=10120 20600 1 0 $X=10005 $Y=19085
X7501 439 78 310 447 78 INV_X1 $T=11070 26200 0 0 $X=10955 $Y=26085
X7502 430 78 310 18 78 INV_X1 $T=11070 37400 1 0 $X=10955 $Y=35885
X7503 730 78 310 60 78 INV_X1 $T=11260 23400 0 0 $X=11145 $Y=23285
X7504 B[15] 78 310 469 78 INV_X1 $T=12590 34600 1 0 $X=12475 $Y=33085
X7505 462 78 310 734 78 INV_X1 $T=13160 3800 0 0 $X=13045 $Y=3685
X7506 460 78 310 48 78 INV_X1 $T=13160 37400 1 0 $X=13045 $Y=35885
X7507 473 78 310 113 78 INV_X1 $T=14680 12200 0 0 $X=14565 $Y=12085
X7508 735 78 310 910 78 INV_X1 $T=14680 17800 1 0 $X=14565 $Y=16285
X7509 739 78 310 934 78 INV_X1 $T=15250 23400 0 0 $X=15135 $Y=23285
X7510 52 78 310 63 78 INV_X1 $T=15440 29000 0 0 $X=15325 $Y=28885
X7511 470 78 310 488 78 INV_X1 $T=16200 9400 0 0 $X=16085 $Y=9285
X7512 490 78 310 743 78 INV_X1 $T=16960 3800 1 0 $X=16845 $Y=2285
X7513 487 78 310 935 78 INV_X1 $T=17340 26200 1 0 $X=17225 $Y=24685
X7514 499 78 310 104 78 INV_X1 $T=17340 29000 0 0 $X=17225 $Y=28885
X7515 868 78 310 91 78 INV_X1 $T=17340 43000 1 0 $X=17225 $Y=41485
X7516 105 78 310 974 78 INV_X1 $T=18100 17800 1 0 $X=17985 $Y=16285
X7517 B[7] 78 310 864 78 INV_X1 $T=18100 34600 1 0 $X=17985 $Y=33085
X7518 755 78 310 103 78 INV_X1 $T=18480 31800 1 0 $X=18365 $Y=30285
X7519 A[7] 78 310 498 78 INV_X1 $T=18670 34600 0 0 $X=18555 $Y=34485
X7520 B[31] 78 310 399 78 INV_X1 $T=18860 15000 0 0 $X=18745 $Y=14885
X7521 496 78 310 914 78 INV_X1 $T=18860 20600 0 0 $X=18745 $Y=20485
X7522 5 78 310 78 78 INV_X1 $T=18860 43000 1 0 $X=18745 $Y=41485
X7523 754 78 310 507 78 INV_X1 $T=19050 6600 1 0 $X=18935 $Y=5085
X7524 526 78 310 506 78 INV_X1 $T=19430 9400 1 0 $X=19315 $Y=7885
X7525 501 78 310 116 78 INV_X1 $T=19810 31800 1 0 $X=19695 $Y=30285
X7526 525 78 310 329 78 INV_X1 $T=20570 15000 1 0 $X=20455 $Y=13485
X7527 865 78 310 130 78 INV_X1 $T=20570 40200 1 0 $X=20455 $Y=38685
X7528 764 78 310 510 78 INV_X1 $T=21140 23400 0 180 $X=20645 $Y=21885
X7529 500 78 310 123 78 INV_X1 $T=21140 34600 1 180 $X=20645 $Y=34485
X7530 504 78 310 511 78 INV_X1 $T=21140 37400 0 0 $X=21025 $Y=37285
X7531 762 78 310 137 78 INV_X1 $T=21520 20600 1 0 $X=21405 $Y=19085
X7532 514 78 310 942 78 INV_X1 $T=23040 34600 0 0 $X=22925 $Y=34485
X7533 766 78 310 135 78 INV_X1 $T=23610 20600 1 180 $X=23115 $Y=20485
X7534 503 78 310 121 78 INV_X1 $T=23420 37400 1 0 $X=23305 $Y=35885
X7535 SUM[31] 78 310 165 78 INV_X1 $T=23800 20600 1 0 $X=23685 $Y=19085
X7536 533 78 310 915 78 INV_X1 $T=24180 26200 0 0 $X=24065 $Y=26085
X7537 172 78 310 152 78 INV_X1 $T=24560 3800 1 0 $X=24445 $Y=2285
X7538 542 78 310 147 78 INV_X1 $T=26460 26200 1 0 $X=26345 $Y=24685
X7539 917 78 310 168 78 INV_X1 $T=26650 43000 0 0 $X=26535 $Y=42885
X7540 546 78 310 548 78 INV_X1 $T=26840 31800 1 0 $X=26725 $Y=30285
X7541 A[26] 78 310 198 78 INV_X1 $T=27030 40200 0 0 $X=26915 $Y=40085
X7542 550 78 310 177 78 INV_X1 $T=27600 17800 1 0 $X=27485 $Y=16285
X7543 173 78 310 565 78 INV_X1 $T=27980 17800 0 0 $X=27865 $Y=17685
X7544 918 78 310 169 78 INV_X1 $T=27980 26200 0 0 $X=27865 $Y=26085
X7545 266 78 310 178 996 INV_X1 $T=28550 1000 0 0 $X=28435 $Y=885
X7546 786 78 310 970 78 INV_X1 $T=28740 17800 1 0 $X=28625 $Y=16285
X7547 571 78 310 784 78 INV_X1 $T=28740 31800 0 0 $X=28625 $Y=31685
X7548 167 78 310 181 78 INV_X1 $T=29310 6600 1 0 $X=29195 $Y=5085
X7549 193 78 310 212 78 INV_X1 $T=29500 9400 0 0 $X=29385 $Y=9285
X7550 191 78 310 170 78 INV_X1 $T=29880 34600 1 0 $X=29765 $Y=33085
X7551 573 78 310 206 78 INV_X1 $T=30260 20600 1 0 $X=30145 $Y=19085
X7552 787 78 310 185 78 INV_X1 $T=30260 29000 0 0 $X=30145 $Y=28885
X7553 A[23] 78 310 568 78 INV_X1 $T=30260 37400 1 0 $X=30145 $Y=35885
X7554 792 78 310 563 78 INV_X1 $T=30450 29000 1 0 $X=30335 $Y=27485
X7555 190 78 310 812 78 INV_X1 $T=31210 12200 1 0 $X=31095 $Y=10685
X7556 569 78 310 962 78 INV_X1 $T=31210 12200 0 0 $X=31095 $Y=12085
X7557 199 78 310 338 78 INV_X1 $T=31400 9400 0 0 $X=31285 $Y=9285
X7558 A[25] 78 310 222 78 INV_X1 $T=31400 40200 1 0 $X=31285 $Y=38685
X7559 291 78 310 205 78 INV_X1 $T=31590 15000 1 0 $X=31475 $Y=13485
X7560 570 78 310 251 78 INV_X1 $T=32160 23400 1 0 $X=32045 $Y=21885
X7561 587 78 310 797 78 INV_X1 $T=33300 29000 1 0 $X=33185 $Y=27485
X7562 588 78 310 977 78 INV_X1 $T=33300 43000 1 0 $X=33185 $Y=41485
X7563 261 78 310 923 78 INV_X1 $T=33680 6600 0 0 $X=33565 $Y=6485
X7564 589 78 310 225 78 INV_X1 $T=33680 9400 1 0 $X=33565 $Y=7885
X7565 227 78 310 346 78 INV_X1 $T=34060 15000 0 0 $X=33945 $Y=14885
X7566 234 78 310 243 78 INV_X1 $T=34060 17800 1 0 $X=33945 $Y=16285
X7567 247 78 310 822 78 INV_X1 $T=34820 17800 0 0 $X=34705 $Y=17685
X7568 241 78 310 244 78 INV_X1 $T=34820 23400 1 0 $X=34705 $Y=21885
X7569 140 78 310 595 78 INV_X1 $T=35010 15000 1 0 $X=34895 $Y=13485
X7570 596 78 310 594 78 INV_X1 $T=35200 17800 1 0 $X=35085 $Y=16285
X7571 257 78 310 256 78 INV_X1 $T=36150 26200 1 0 $X=36035 $Y=24685
X7572 229 78 310 280 78 INV_X1 $T=36340 23400 1 0 $X=36225 $Y=21885
X7573 194 78 310 263 78 INV_X1 $T=36720 15000 0 0 $X=36605 $Y=14885
X7574 607 78 310 218 78 INV_X1 $T=37290 12200 0 0 $X=37175 $Y=12085
X7575 A[30] 78 310 360 78 INV_X1 $T=38240 43000 0 180 $X=37745 $Y=41485
X7576 B[28] 78 310 887 78 INV_X1 $T=38810 40200 1 0 $X=38695 $Y=38685
X7577 811 78 310 284 78 INV_X1 $T=39000 26200 1 0 $X=38885 $Y=24685
X7578 626 78 310 629 78 INV_X1 $T=39950 6600 1 0 $X=39835 $Y=5085
X7579 250 78 310 265 78 INV_X1 $T=40140 12200 0 0 $X=40025 $Y=12085
X7580 366 78 310 618 78 INV_X1 $T=41090 26200 0 0 $X=40975 $Y=26085
X7581 287 78 310 952 78 INV_X1 $T=41090 34600 0 0 $X=40975 $Y=34485
X7582 628 78 310 294 78 INV_X1 $T=41090 43000 0 0 $X=40975 $Y=42885
X7583 631 78 310 836 78 INV_X1 $T=41470 12200 1 0 $X=41355 $Y=10685
X7584 638 78 310 363 78 INV_X1 $T=41850 12200 0 0 $X=41735 $Y=12085
X7585 599 78 310 894 78 INV_X1 $T=43180 31800 1 0 $X=43065 $Y=30285
X7586 78 310 668 897 ICV_10 $T=1380 15000 0 0 $X=1265 $Y=14885
X7587 78 310 391 412 ICV_10 $T=2330 3800 1 0 $X=2215 $Y=2285
X7588 78 310 386 689 ICV_10 $T=4230 23400 1 0 $X=4115 $Y=21885
X7589 78 310 466 853 ICV_10 $T=6130 6600 0 0 $X=6015 $Y=6485
X7590 78 310 420 42 ICV_10 $T=6130 23400 1 0 $X=6015 $Y=21885
X7591 78 310 418 706 ICV_10 $T=7080 6600 0 0 $X=6965 $Y=6485
X7592 78 310 3 696 ICV_10 $T=7650 40200 1 0 $X=7535 $Y=38685
X7593 78 310 446 73 ICV_10 $T=11070 15000 1 0 $X=10955 $Y=13485
X7594 78 310 320 449 ICV_10 $T=11640 3800 1 0 $X=11525 $Y=2285
X7595 78 310 467 737 ICV_10 $T=14300 6600 0 0 $X=14185 $Y=6485
X7596 78 310 330 870 ICV_10 $T=22280 31800 1 0 $X=22165 $Y=30285
X7597 78 310 331 765 ICV_10 $T=22660 23400 0 0 $X=22545 $Y=23285
X7598 78 310 202 187 ICV_10 $T=28360 9400 1 0 $X=28245 $Y=7885
X7599 78 310 B[27] 209 ICV_10 $T=30260 43000 0 0 $X=30145 $Y=42885
X7600 78 310 259 602 ICV_10 $T=35960 17800 0 0 $X=35845 $Y=17685
X7601 78 310 613 286 ICV_10 $T=39570 37400 1 0 $X=39455 $Y=35885
X7602 78 310 637 299 ICV_10 $T=40520 6600 1 0 $X=40405 $Y=5085
X7603 78 310 237 254 ICV_10 $T=42040 3800 0 0 $X=41925 $Y=3685
X7604 78 310 661 368 ICV_10 $T=43750 29000 0 0 $X=43635 $Y=28885
X7605 335 78 561 180 780 214 310 NAND4_X1 $T=28930 12200 0 0 $X=28815 $Y=12085
X7606 583 78 922 972 586 570 310 NAND4_X1 $T=32540 20600 1 0 $X=32425 $Y=19085
X7607 B[27] 78 B[28] B[29] B[30] 644 310 NAND4_X1 $T=41470 26200 0 0 $X=41355 $Y=26085
X7608 B[23] 78 B[24] B[25] B[26] 654 310 NAND4_X1 $T=42610 26200 1 0 $X=42495 $Y=24685
X7609 A[27] 78 A[28] A[29] A[30] 967 310 NAND4_X1 $T=43750 23400 0 0 $X=43635 $Y=23285
X7610 A[23] 78 A[24] A[25] A[26] 895 310 NAND4_X1 $T=44700 29000 0 180 $X=43635 $Y=27485
X7611 376 36 78 2 32 383 310 78 OAI22_X1 $T=1000 31800 1 0 $X=885 $Y=30285
X7612 315 405 78 394 35 64 310 78 OAI22_X1 $T=3280 34600 0 180 $X=2215 $Y=33085
X7613 375 399 78 408 B[31] 397 310 78 OAI22_X1 $T=3090 12200 1 0 $X=2975 $Y=10685
X7614 673 A[31] 78 683 551 396 310 78 OAI22_X1 $T=3280 17800 0 0 $X=3165 $Y=17685
X7615 666 35 78 403 38 315 310 78 OAI22_X1 $T=4230 34600 0 180 $X=3165 $Y=33085
X7616 682 399 78 413 B[31] 395 310 78 OAI22_X1 $T=3660 6600 0 0 $X=3545 $Y=6485
X7617 387 A[31] 78 688 551 693 310 78 OAI22_X1 $T=4230 20600 0 0 $X=4115 $Y=20485
X7618 679 A[31] 78 425 551 689 310 78 OAI22_X1 $T=4800 23400 1 0 $X=4685 $Y=21885
X7619 848 399 78 423 B[31] 412 310 78 OAI22_X1 $T=5180 3800 0 0 $X=5065 $Y=3685
X7620 46 35 78 415 852 315 310 78 OAI22_X1 $T=5180 34600 1 0 $X=5065 $Y=33085
X7621 26 399 78 418 B[31] 15 310 78 OAI22_X1 $T=5750 6600 1 0 $X=5635 $Y=5085
X7622 404 852 78 29 36 416 310 78 OAI22_X1 $T=5940 31800 1 0 $X=5825 $Y=30285
X7623 48 405 78 322 696 24 310 78 OAI22_X1 $T=5940 37400 0 0 $X=5825 $Y=37285
X7624 702 399 78 714 B[31] 410 310 996 OAI22_X1 $T=6320 1000 0 0 $X=6205 $Y=885
X7625 419 399 78 433 B[31] 695 310 78 OAI22_X1 $T=6510 17800 1 0 $X=6395 $Y=16285
X7626 312 696 78 318 852 48 310 78 OAI22_X1 $T=6890 37400 0 0 $X=6775 $Y=37285
X7627 709 712 78 716 18 700 310 78 OAI22_X1 $T=8980 40200 0 0 $X=8865 $Y=40085
X7628 855 A[31] 78 718 551 932 310 78 OAI22_X1 $T=9360 20600 0 0 $X=9245 $Y=20485
X7629 432 A[31] 78 56 551 931 310 78 OAI22_X1 $T=9360 23400 0 0 $X=9245 $Y=23285
X7630 5 436 78 442 960 355 310 78 OAI22_X1 $T=10500 17800 0 0 $X=10385 $Y=17685
X7631 723 696 78 725 64 48 310 78 OAI22_X1 $T=10690 37400 0 0 $X=10575 $Y=37285
X7632 71 696 78 80 721 48 310 78 OAI22_X1 $T=10880 40200 0 0 $X=10765 $Y=40085
X7633 731 36 78 76 32 319 310 78 OAI22_X1 $T=12590 31800 0 0 $X=12475 $Y=31685
X7634 464 399 78 735 B[31] 75 310 78 OAI22_X1 $T=13540 15000 0 0 $X=13425 $Y=14885
X7635 80 18 78 478 430 933 310 78 OAI22_X1 $T=14110 37400 1 0 $X=13995 $Y=35885
X7636 321 32 78 96 36 857 310 78 OAI22_X1 $T=14490 34600 0 0 $X=14375 $Y=34485
X7637 738 36 78 110 32 860 310 78 OAI22_X1 $T=15820 40200 1 0 $X=15705 $Y=38685
X7638 740 36 78 112 32 857 310 78 OAI22_X1 $T=16770 37400 0 0 $X=16655 $Y=37285
X7639 481 A[31] 78 750 551 935 310 78 OAI22_X1 $T=16960 23400 0 0 $X=16845 $Y=23285
X7640 5 864 78 107 498 78 310 78 OAI22_X1 $T=17720 34600 0 0 $X=17605 $Y=34485
X7641 118 SUM[31] 78 253 165 760 310 78 OAI22_X1 $T=20950 3800 0 0 $X=20835 $Y=3685
X7642 754 SUM[31] 78 211 165 938 310 78 OAI22_X1 $T=21710 6600 1 0 $X=21595 $Y=5085
X7643 127 SUM[31] 78 266 165 517 310 996 OAI22_X1 $T=22280 1000 0 0 $X=22165 $Y=885
X7644 761 SUM[31] 78 199 165 757 310 78 OAI22_X1 $T=22280 6600 0 0 $X=22165 $Y=6485
X7645 756 SUM[31] 78 190 165 515 310 78 OAI22_X1 $T=22280 12200 0 0 $X=22165 $Y=12085
X7646 520 399 78 764 B[31] 135 310 78 OAI22_X1 $T=22280 23400 1 0 $X=22165 $Y=21885
X7647 500 A[31] 78 775 551 941 310 78 OAI22_X1 $T=22660 31800 0 0 $X=22545 $Y=31685
X7648 501 A[31] 78 524 551 870 310 78 OAI22_X1 $T=22850 31800 1 0 $X=22735 $Y=30285
X7649 529 399 78 331 B[31] 137 310 78 OAI22_X1 $T=24180 23400 0 180 $X=23115 $Y=21885
X7650 525 SUM[31] 78 140 165 940 310 78 OAI22_X1 $T=23420 15000 1 0 $X=23305 $Y=13485
X7651 526 SUM[31] 78 202 165 531 310 78 OAI22_X1 $T=23610 9400 1 0 $X=23495 $Y=7885
X7652 752 SUM[31] 78 193 165 769 310 78 OAI22_X1 $T=23990 9400 0 0 $X=23875 $Y=9285
X7653 144 399 78 533 B[31] 147 310 78 OAI22_X1 $T=24180 26200 1 0 $X=24065 $Y=24685
X7654 143 SUM[31] 78 167 165 771 310 78 OAI22_X1 $T=26080 6600 0 0 $X=25965 $Y=6485
X7655 768 SUM[31] 78 180 165 534 310 78 OAI22_X1 $T=26270 3800 0 0 $X=26155 $Y=3685
X7656 156 SUM[31] 78 234 165 774 310 78 OAI22_X1 $T=26650 20600 0 0 $X=26535 $Y=20485
X7657 141 SUM[31] 78 780 165 555 310 78 OAI22_X1 $T=27220 3800 1 0 $X=27105 $Y=2285
X7658 778 399 78 546 B[31] 563 310 78 OAI22_X1 $T=27220 29000 0 0 $X=27105 $Y=28885
X7659 779 552 78 164 213 562 310 78 OAI22_X1 $T=27410 37400 0 0 $X=27295 $Y=37285
X7660 5 216 78 267 198 355 310 78 OAI22_X1 $T=27410 40200 0 0 $X=27295 $Y=40085
X7661 5 213 78 248 552 355 310 78 OAI22_X1 $T=27600 37400 1 0 $X=27485 $Y=35885
X7662 779 568 78 149 578 562 310 78 OAI22_X1 $T=29500 37400 0 0 $X=29385 $Y=37285
X7663 174 SUM[31] 78 194 165 566 310 78 OAI22_X1 $T=29690 23400 1 0 $X=29575 $Y=21885
X7664 779 217 78 344 209 562 310 78 OAI22_X1 $T=30830 43000 0 0 $X=30715 $Y=42885
X7665 5 794 78 240 222 355 310 78 OAI22_X1 $T=31780 40200 1 0 $X=31665 $Y=38685
X7666 5 209 78 276 217 355 310 78 OAI22_X1 $T=31780 43000 0 0 $X=31665 $Y=42885
X7667 218 211 78 277 242 348 310 78 OAI22_X1 $T=32160 9400 1 0 $X=32045 $Y=7885
X7668 231 194 78 590 589 962 310 78 OAI22_X1 $T=33490 15000 1 0 $X=33375 $Y=13485
X7669 591 589 78 801 274 231 310 78 OAI22_X1 $T=34060 9400 1 0 $X=33945 $Y=7885
X7670 584 260 78 589 610 275 310 78 OAI22_X1 $T=34630 20600 0 0 $X=34515 $Y=20485
X7671 218 187 78 601 243 607 310 78 OAI22_X1 $T=35770 9400 1 0 $X=35655 $Y=7885
X7672 218 812 78 353 263 607 310 78 OAI22_X1 $T=36150 12200 1 0 $X=36035 $Y=10685
X7673 218 338 78 606 346 607 310 78 OAI22_X1 $T=36530 9400 0 0 $X=36415 $Y=9285
X7674 218 597 78 608 822 607 310 78 OAI22_X1 $T=36720 15000 1 0 $X=36605 $Y=13485
X7675 218 212 78 612 609 607 310 78 OAI22_X1 $T=37100 12200 1 0 $X=36985 $Y=10685
X7676 800 254 78 262 237 829 310 78 OAI22_X1 $T=37480 3800 0 0 $X=37365 $Y=3685
X7677 218 595 78 620 359 607 310 78 OAI22_X1 $T=37670 15000 1 0 $X=37555 $Y=13485
X7678 622 221 78 624 247 825 310 78 OAI22_X1 $T=38050 23400 1 0 $X=37935 $Y=21885
X7679 622 194 78 358 259 825 310 78 OAI22_X1 $T=38240 20600 0 0 $X=38125 $Y=20485
X7680 821 254 78 817 237 965 310 78 OAI22_X1 $T=38430 3800 0 0 $X=38315 $Y=3685
X7681 620 615 78 626 606 630 310 78 OAI22_X1 $T=39000 9400 1 0 $X=38885 $Y=7885
X7682 827 616 78 SUM[2] 221 340 310 78 OAI22_X1 $T=39190 23400 0 0 $X=39075 $Y=23285
X7683 361 274 78 635 250 608 310 78 OAI22_X1 $T=40140 15000 1 0 $X=40025 $Y=13485
X7684 265 194 78 833 242 250 310 78 OAI22_X1 $T=40710 15000 0 0 $X=40595 $Y=14885
X7685 636 278 78 301 649 363 310 78 OAI22_X1 $T=42230 15000 1 0 $X=42115 $Y=13485
X7686 629 254 78 929 237 840 310 78 OAI22_X1 $T=42610 3800 0 0 $X=42495 $Y=3685
X7687 646 648 78 308 254 299 310 78 OAI22_X1 $T=42610 6600 1 0 $X=42495 $Y=5085
X7688 363 648 78 365 646 649 310 78 OAI22_X1 $T=42610 9400 0 0 $X=42495 $Y=9285
X7689 644 654 78 366 895 967 310 78 OAI22_X1 $T=42990 26200 0 0 $X=42875 $Y=26085
X7690 953 811 78 661 894 964 310 78 OAI22_X1 $T=43560 31800 1 0 $X=43445 $Y=30285
X7691 968 616 78 SUM[7] 242 340 310 78 OAI22_X1 $T=43750 17800 0 0 $X=43635 $Y=17685
X7692 658 616 78 SUM[5] 234 340 310 78 OAI22_X1 $T=43750 23400 1 0 $X=43635 $Y=21885
X7757 310 397 375 844 78 78 XOR2_X1 $T=2140 9400 0 180 $X=885 $Y=7885
X7758 310 6 384 671 78 78 XOR2_X1 $T=1000 12200 0 0 $X=885 $Y=12085
X7759 310 4 385 670 78 78 XOR2_X1 $T=1000 17800 0 0 $X=885 $Y=17685
X7760 310 381 386 311 78 78 XOR2_X1 $T=1000 23400 1 0 $X=885 $Y=21885
X7761 310 412 848 414 78 78 XOR2_X1 $T=2900 3800 0 0 $X=2785 $Y=3685
X7762 310 15 26 691 78 78 XOR2_X1 $T=3850 6600 1 0 $X=3735 $Y=5085
X7763 310 28 703 678 78 78 XOR2_X1 $T=4610 20600 1 0 $X=4495 $Y=19085
X7764 310 31 699 901 78 78 XOR2_X1 $T=4990 26200 1 0 $X=4875 $Y=24685
X7765 310 695 419 732 78 78 XOR2_X1 $T=5180 15000 1 0 $X=5065 $Y=13485
X7766 310 60 443 61 78 78 XOR2_X1 $T=9930 23400 1 0 $X=9815 $Y=21885
X7767 310 447 452 450 78 78 XOR2_X1 $T=11260 26200 1 0 $X=11145 $Y=24685
X7768 310 81 487 86 78 78 XOR2_X1 $T=15060 26200 1 0 $X=14945 $Y=24685
X7769 310 92 491 475 78 996 XOR2_X1 $T=15630 1000 0 0 $X=15515 $Y=885
X7770 310 90 744 88 78 78 XOR2_X1 $T=16010 29000 1 0 $X=15895 $Y=27485
X7771 310 103 748 106 78 78 XOR2_X1 $T=18480 29000 0 0 $X=18365 $Y=28885
X7772 310 118 760 505 78 78 XOR2_X1 $T=19050 3800 0 0 $X=18935 $Y=3685
X7773 310 123 753 509 78 78 XOR2_X1 $T=19620 34600 1 0 $X=19505 $Y=33085
X7774 310 116 330 912 78 78 XOR2_X1 $T=20190 31800 0 0 $X=20075 $Y=31685
X7775 310 756 515 758 78 78 XOR2_X1 $T=20380 12200 0 0 $X=20265 $Y=12085
X7776 310 761 757 937 78 78 XOR2_X1 $T=20570 6600 0 0 $X=20455 $Y=6485
X7777 310 127 517 512 78 996 XOR2_X1 $T=21140 1000 0 0 $X=21025 $Y=885
X7778 310 147 144 554 78 78 XOR2_X1 $T=23040 26200 1 0 $X=22925 $Y=24685
X7779 310 137 529 129 78 78 XOR2_X1 $T=23800 20600 0 0 $X=23685 $Y=20485
X7780 310 121 770 130 78 78 XOR2_X1 $T=23990 34600 0 0 $X=23875 $Y=34485
X7781 310 169 537 557 78 78 XOR2_X1 $T=26080 26200 0 0 $X=25965 $Y=26085
X7782 310 174 566 781 78 78 XOR2_X1 $T=28550 23400 1 0 $X=28435 $Y=21885
X7783 310 184 581 336 78 78 XOR2_X1 $T=30830 23400 0 0 $X=30715 $Y=23285
X7784 310 197 592 201 78 78 XOR2_X1 $T=33110 26200 1 0 $X=32995 $Y=24685
X7785 310 663 927 660 78 78 XOR2_X1 $T=44700 43000 0 180 $X=43445 $Y=41485
X8081 78 310 376 32 393 36 39 ICV_19 $T=2330 31800 1 0 $X=2215 $Y=30285
X8082 78 310 384 399 692 B[31] 6 ICV_19 $T=3280 12200 0 0 $X=3165 $Y=12085
X8083 78 310 361 227 631 250 620 ICV_19 $T=39760 12200 1 0 $X=39645 $Y=10685
X8084 78 310 269 292 632 278 963 ICV_19 $T=39760 17800 0 0 $X=39645 $Y=17685
X8085 78 310 965 254 298 237 299 ICV_19 $T=40330 3800 0 0 $X=40215 $Y=3685
X8086 78 310 255 615 637 601 630 ICV_19 $T=40520 9400 1 0 $X=40405 $Y=7885
X8087 78 310 292 278 305 649 892 ICV_19 $T=42230 15000 0 0 $X=42115 $Y=14885
X8088 78 310 652 616 SUM[6] 227 340 ICV_19 $T=42990 20600 1 0 $X=42875 $Y=19085
X8097 78 310 398 399 401 B[31] 668 ICV_21 $T=3090 17800 1 0 $X=2975 $Y=16285
X8098 78 310 402 A[31] 406 551 684 ICV_21 $T=3850 26200 1 0 $X=3735 $Y=24685
X8099 78 310 313 696 14 38 48 ICV_21 $T=4800 37400 1 0 $X=4685 $Y=35885
X8100 78 310 5 960 711 436 355 ICV_21 $T=8980 20600 1 0 $X=8865 $Y=19085
X8101 78 310 486 551 489 A[31] 82 ICV_21 $T=15820 20600 1 0 $X=15705 $Y=19085
X8102 78 310 779 222 785 794 562 ICV_21 $T=28550 40200 0 0 $X=28435 $Y=40085
X8103 78 310 608 615 828 612 630 ICV_21 $T=39190 6600 0 0 $X=39075 $Y=6485
X8104 78 310 645 616 SUM[4] 274 340 ICV_21 $T=40710 20600 0 0 $X=40595 $Y=20485
X8105 78 310 892 648 304 836 649 ICV_21 $T=42230 12200 1 0 $X=42115 $Y=10685
X8106 78 310 634 229 658 280 640 ICV_21 $T=42610 20600 0 0 $X=42495 $Y=20485
X8107 42 40 51 43 78 310 78 OAI21_X1 $T=6890 20600 0 0 $X=6775 $Y=20485
X8108 19 46 709 854 78 310 78 OAI21_X1 $T=7650 43000 1 0 $X=7535 $Y=41485
X8109 317 48 712 18 78 310 78 OAI21_X1 $T=8220 40200 0 0 $X=8105 $Y=40085
X8110 905 35 54 52 78 310 78 OAI21_X1 $T=8790 29000 0 0 $X=8675 $Y=28885
X8111 60 61 65 62 78 310 78 OAI21_X1 $T=11070 23400 1 0 $X=10955 $Y=21885
X8112 723 48 908 453 78 310 78 OAI21_X1 $T=11640 43000 1 0 $X=11525 $Y=41485
X8113 451 63 729 440 78 310 78 OAI21_X1 $T=12020 31800 1 0 $X=11905 $Y=30285
X8114 73 74 70 75 78 310 78 OAI21_X1 $T=13160 12200 0 0 $X=13045 $Y=12085
X8115 81 86 85 83 78 310 78 OAI21_X1 $T=14300 26200 0 0 $X=14185 $Y=26085
X8116 67 91 324 484 78 310 78 OAI21_X1 $T=15060 37400 1 0 $X=14945 $Y=35885
X8117 103 106 111 104 78 310 78 OAI21_X1 $T=17720 29000 0 0 $X=17605 $Y=28885
X8118 130 121 132 511 78 310 78 OAI21_X1 $T=20190 37400 1 0 $X=20075 $Y=35885
X8119 117 124 128 119 78 310 78 OAI21_X1 $T=20760 17800 0 0 $X=20645 $Y=17685
X8120 137 129 131 135 78 310 78 OAI21_X1 $T=20950 20600 0 0 $X=20835 $Y=20485
X8121 527 142 150 768 78 310 78 OAI21_X1 $T=23800 3800 0 0 $X=23685 $Y=3685
X8122 141 152 157 143 78 310 78 OAI21_X1 $T=24560 6600 0 0 $X=24445 $Y=6485
X8123 155 161 163 156 78 310 78 OAI21_X1 $T=25510 23400 1 0 $X=25395 $Y=21885
X8124 166 154 871 547 78 310 78 OAI21_X1 $T=25700 17800 1 0 $X=25585 $Y=16285
X8125 541 165 550 547 78 310 78 OAI21_X1 $T=26270 15000 0 0 $X=26155 $Y=14885
X8126 541 166 543 547 78 310 78 OAI21_X1 $T=26460 17800 1 0 $X=26345 $Y=16285
X8127 782 171 179 561 78 310 78 OAI21_X1 $T=27220 12200 0 0 $X=27105 $Y=12085
X8128 158 173 559 SUM[31] 78 310 78 OAI21_X1 $T=27600 15000 0 0 $X=27485 $Y=14885
X8129 556 177 874 559 78 310 78 OAI21_X1 $T=27980 17800 1 0 $X=27865 $Y=16285
X8130 253 178 875 220 78 310 78 OAI21_X1 $T=28170 3800 1 0 $X=28055 $Y=2285
X8131 945 181 876 208 78 310 78 OAI21_X1 $T=28550 6600 1 0 $X=28435 $Y=5085
X8132 170 185 176 563 78 310 78 OAI21_X1 $T=28740 29000 1 0 $X=28625 $Y=27485
X8133 919 187 175 199 78 310 78 OAI21_X1 $T=28930 9400 1 0 $X=28815 $Y=7885
X8134 920 189 786 335 78 310 78 OAI21_X1 $T=29120 17800 1 0 $X=29005 $Y=16285
X8135 565 165 793 543 78 310 78 OAI21_X1 $T=29120 17800 0 0 $X=29005 $Y=17685
X8136 340 193 SUM[12] 572 78 310 78 OAI21_X1 $T=29690 9400 1 0 $X=29575 $Y=7885
X8137 340 780 SUM[20] 788 78 310 996 OAI21_X1 $T=29880 1000 0 0 $X=29765 $Y=885
X8138 607 190 569 180 78 310 78 OAI21_X1 $T=29880 12200 0 0 $X=29765 $Y=12085
X8139 970 196 573 543 78 310 78 OAI21_X1 $T=29880 17800 1 0 $X=29765 $Y=16285
X8140 607 199 574 208 78 310 78 OAI21_X1 $T=30070 6600 0 0 $X=29955 $Y=6485
X8141 586 200 334 789 78 310 78 OAI21_X1 $T=30070 15000 0 0 $X=29955 $Y=14885
X8142 201 197 207 582 78 310 78 OAI21_X1 $T=30260 26200 0 0 $X=30145 $Y=26085
X8143 340 180 SUM[19] 342 78 310 996 OAI21_X1 $T=30640 1000 0 0 $X=30525 $Y=885
X8144 340 199 SUM[14] 343 78 310 78 OAI21_X1 $T=30640 3800 1 0 $X=30525 $Y=2285
X8145 921 205 576 140 78 310 78 OAI21_X1 $T=30830 15000 1 0 $X=30715 $Y=13485
X8146 340 208 SUM[22] 580 78 310 78 OAI21_X1 $T=31020 6600 1 0 $X=30905 $Y=5085
X8147 340 211 SUM[15] 656 78 310 78 OAI21_X1 $T=31400 3800 0 0 $X=31285 $Y=3685
X8148 922 214 257 584 78 310 78 OAI21_X1 $T=31780 20600 0 0 $X=31665 $Y=20485
X8149 231 227 796 229 78 310 78 OAI21_X1 $T=33110 9400 0 0 $X=32995 $Y=9285
X8150 229 241 237 238 78 310 78 OAI21_X1 $T=34250 20600 1 0 $X=34135 $Y=19085
X8151 594 243 946 227 78 310 78 OAI21_X1 $T=34440 17800 1 0 $X=34325 $Y=16285
X8152 351 252 270 598 78 310 78 OAI21_X1 $T=35200 43000 1 0 $X=35085 $Y=41485
X8153 810 252 600 598 78 310 78 OAI21_X1 $T=35580 43000 0 0 $X=35465 $Y=42885
X8154 360 B[30] 779 600 78 310 78 OAI21_X1 $T=36340 43000 0 0 $X=36225 $Y=42885
X8155 925 263 596 274 78 310 78 OAI21_X1 $T=37100 15000 0 0 $X=36985 $Y=14885
X8156 622 259 819 280 78 310 78 OAI21_X1 $T=37290 23400 1 0 $X=37175 $Y=21885
X8157 340 266 SUM[17] 627 78 310 996 OAI21_X1 $T=38430 1000 0 0 $X=38315 $Y=885
X8158 624 280 827 819 78 310 78 OAI21_X1 $T=39000 23400 1 0 $X=38885 $Y=21885
X8159 340 190 SUM[11] 830 78 310 78 OAI21_X1 $T=39760 9400 0 0 $X=39645 $Y=9285
X8160 340 253 SUM[16] 832 78 310 78 OAI21_X1 $T=40330 3800 1 0 $X=40215 $Y=2285
X8161 340 291 SUM[9] 643 78 310 78 OAI21_X1 $T=41090 15000 1 0 $X=40975 $Y=13485
X8162 78 310 19 448 64 18 78 ICV_22 $T=11070 40200 1 0 $X=10955 $Y=38685
X8163 78 310 79 87 84 82 78 ICV_22 $T=14110 20600 0 0 $X=13995 $Y=20485
X8164 78 310 565 577 165 570 78 ICV_22 $T=29310 20600 1 0 $X=29195 $Y=19085
X8165 78 310 340 SUM[13] 202 841 78 ICV_22 $T=30070 6600 1 0 $X=29955 $Y=5085
X8166 78 310 340 SUM[21] 167 791 78 ICV_22 $T=30450 3800 0 0 $X=30335 $Y=3685
X8167 78 310 340 SUM[18] 220 619 996 ICV_22 $T=32540 1000 0 0 $X=32425 $Y=885
X8168 78 310 340 SUM[10] 140 657 78 ICV_22 $T=42610 12200 0 0 $X=42495 $Y=12085
X8169 78 310 340 SUM[8] 297 367 78 ICV_22 $T=42610 17800 1 0 $X=42495 $Y=16285
X8193 14 18 39 409 78 310 AOI21_X1 $T=4990 34600 0 0 $X=4875 $Y=34485
X8194 322 18 704 316 78 310 AOI21_X1 $T=6890 37400 1 0 $X=6775 $Y=35885
X8195 318 18 719 856 78 310 AOI21_X1 $T=8410 34600 0 0 $X=8295 $Y=34485
X8196 905 63 62 729 78 310 AOI21_X1 $T=11260 29000 0 0 $X=11145 $Y=28885
X8197 38 63 79 476 78 310 AOI21_X1 $T=12400 29000 1 0 $X=12285 $Y=27485
X8198 785 153 911 773 78 310 AOI21_X1 $T=24560 40200 0 0 $X=24445 $Y=40085
X8199 539 160 913 917 78 310 AOI21_X1 $T=25320 43000 1 0 $X=25205 $Y=41485
X8200 149 164 540 873 78 310 AOI21_X1 $T=25890 40200 1 0 $X=25775 $Y=38685
X8201 344 168 916 558 78 310 AOI21_X1 $T=27030 43000 0 0 $X=26915 $Y=42885
X8202 333 175 556 876 78 310 AOI21_X1 $T=27790 6600 0 0 $X=27675 $Y=6485
X8203 871 179 241 577 78 310 AOI21_X1 $T=28360 17800 0 0 $X=28245 $Y=17685
X8204 875 180 945 877 78 310 AOI21_X1 $T=28550 3800 0 0 $X=28435 $Y=3685
X8205 576 190 919 212 78 310 AOI21_X1 $T=29500 12200 1 0 $X=29385 $Y=10685
X8206 218 187 239 181 78 310 AOI21_X1 $T=30830 6600 0 0 $X=30715 $Y=6485
X8207 795 210 920 575 78 310 AOI21_X1 $T=31210 17800 1 0 $X=31095 $Y=16285
X8208 218 212 591 877 78 310 AOI21_X1 $T=31400 9400 1 0 $X=31285 $Y=7885
X8209 A[26] 216 347 588 78 310 AOI21_X1 $T=32350 40200 0 0 $X=32235 $Y=40085
X8210 259 221 585 798 78 310 AOI21_X1 $T=32730 17800 0 0 $X=32615 $Y=17685
X8211 574 225 228 796 78 310 AOI21_X1 $T=32920 6600 0 0 $X=32805 $Y=6485
X8212 946 242 921 597 78 310 AOI21_X1 $T=34440 15000 0 0 $X=34325 $Y=14885
X8213 268 250 230 801 78 310 AOI21_X1 $T=35010 6600 0 0 $X=34895 $Y=6485
X8214 816 250 947 802 78 310 AOI21_X1 $T=35010 9400 1 0 $X=34895 $Y=7885
X8215 806 254 226 947 78 310 AOI21_X1 $T=35770 6600 1 0 $X=35655 $Y=5085
X8216 261 265 800 948 78 310 AOI21_X1 $T=36530 6600 1 0 $X=36415 $Y=5085
X8217 816 265 821 886 78 310 AOI21_X1 $T=36720 9400 1 0 $X=36605 $Y=7885
X8218 268 265 829 820 78 310 AOI21_X1 $T=37290 6600 1 0 $X=37175 $Y=5085
X8219 822 259 925 359 78 310 AOI21_X1 $T=37860 15000 0 0 $X=37745 $Y=14885
X8220 277 265 965 625 78 310 AOI21_X1 $T=39190 6600 1 0 $X=39075 $Y=5085
X8221 251 286 639 362 78 310 AOI21_X1 $T=39950 31800 1 0 $X=39835 $Y=30285
X8222 354 288 926 628 78 310 AOI21_X1 $T=40330 43000 0 0 $X=40215 $Y=42885
X8223 604 294 928 660 78 310 AOI21_X1 $T=42230 43000 0 0 $X=42115 $Y=42885
X8224 381 310 311 10 78 78 NOR2_X1 $T=1380 26200 1 0 $X=1265 $Y=24685
X8225 397 310 844 7 78 78 NOR2_X1 $T=2330 9400 0 0 $X=2215 $Y=9285
X8226 666 310 315 409 78 78 NOR2_X1 $T=4420 34600 0 0 $X=4305 $Y=34485
X8227 412 310 414 22 78 996 NOR2_X1 $T=4610 1000 0 0 $X=4495 $Y=885
X8228 695 310 732 8 78 78 NOR2_X1 $T=5180 15000 0 0 $X=5065 $Y=14885
X8229 696 310 18 903 78 78 NOR2_X1 $T=5750 34600 0 0 $X=5635 $Y=34485
X8230 903 310 859 416 78 78 NOR2_X1 $T=6890 34600 1 0 $X=6775 $Y=33085
X8231 64 310 315 316 78 78 NOR2_X1 $T=7080 34600 0 0 $X=6965 $Y=34485
X8232 46 310 315 856 78 78 NOR2_X1 $T=7460 34600 1 0 $X=7345 $Y=33085
X8233 696 310 430 57 78 78 NOR2_X1 $T=9170 34600 0 0 $X=9055 $Y=34485
X8234 711 310 36 905 78 78 NOR2_X1 $T=9550 29000 0 0 $X=9435 $Y=28885
X8235 721 310 696 859 78 78 NOR2_X1 $T=10120 37400 0 0 $X=10005 $Y=37285
X8236 38 310 36 451 78 78 NOR2_X1 $T=11450 31800 1 0 $X=11335 $Y=30285
X8237 447 310 450 50 78 78 NOR2_X1 $T=11640 23400 0 0 $X=11525 $Y=23285
X8238 442 310 468 69 78 78 NOR2_X1 $T=13160 9400 1 0 $X=13045 $Y=7885
X8239 91 310 77 460 78 78 NOR2_X1 $T=13540 37400 1 0 $X=13425 $Y=35885
X8240 476 310 52 82 78 78 NOR2_X1 $T=14300 29000 1 0 $X=14185 $Y=27485
X8241 868 310 77 3 78 78 NOR2_X1 $T=17720 43000 1 0 $X=17605 $Y=41485
X8242 761 310 937 122 78 78 NOR2_X1 $T=20000 6600 0 0 $X=19885 $Y=6485
X8243 749 310 513 134 78 78 NOR2_X1 $T=20000 15000 0 0 $X=19885 $Y=14885
X8244 756 310 758 138 78 78 NOR2_X1 $T=21140 9400 0 0 $X=21025 $Y=9285
X8245 528 310 532 767 78 78 NOR2_X1 $T=23990 12200 1 0 $X=23875 $Y=10685
X8246 162 310 SUM[31] 173 78 78 NOR2_X1 $T=25130 15000 1 0 $X=25015 $Y=13485
X8247 785 310 153 773 78 78 NOR2_X1 $T=25320 40200 0 0 $X=25205 $Y=40085
X8248 539 310 160 917 78 78 NOR2_X1 $T=26080 43000 1 0 $X=25965 $Y=41485
X8249 149 310 164 873 78 78 NOR2_X1 $T=26650 40200 1 0 $X=26535 $Y=38685
X8250 339 310 549 553 78 78 NOR2_X1 $T=26840 9400 0 0 $X=26725 $Y=9285
X8251 549 310 776 335 78 78 NOR2_X1 $T=27220 12200 1 0 $X=27105 $Y=10685
X8252 553 310 776 782 78 78 NOR2_X1 $T=27790 12200 1 0 $X=27675 $Y=10685
X8253 344 310 168 558 78 78 NOR2_X1 $T=27790 43000 0 0 $X=27675 $Y=42885
X8254 575 310 189 922 78 78 NOR2_X1 $T=30640 17800 1 0 $X=30525 $Y=16285
X8255 812 310 212 182 78 78 NOR2_X1 $T=30830 9400 0 0 $X=30715 $Y=9285
X8256 214 310 793 583 78 78 NOR2_X1 $T=31400 17800 0 0 $X=31285 $Y=17685
X8257 205 310 595 789 78 78 NOR2_X1 $T=32160 15000 1 0 $X=32045 $Y=13485
X8258 251 310 793 584 78 78 NOR2_X1 $T=32540 20600 0 0 $X=32425 $Y=20485
X8259 243 310 346 795 78 78 NOR2_X1 $T=32730 15000 0 0 $X=32615 $Y=14885
X8260 217 310 B[27] 588 78 78 NOR2_X1 $T=32730 43000 1 0 $X=32615 $Y=41485
X8261 206 310 238 260 78 78 NOR2_X1 $T=34060 20600 0 0 $X=33945 $Y=20485
X8262 263 310 609 210 78 78 NOR2_X1 $T=36720 17800 1 0 $X=36605 $Y=16285
X8263 256 310 260 610 78 78 NOR2_X1 $T=37480 20600 1 180 $X=36795 $Y=20485
X8264 606 310 615 948 78 78 NOR2_X1 $T=37100 6600 0 0 $X=36985 $Y=6485
X8265 601 310 615 886 78 78 NOR2_X1 $T=37480 9400 1 0 $X=37365 $Y=7885
X8266 612 310 615 820 78 78 NOR2_X1 $T=38050 6600 1 0 $X=37935 $Y=5085
X8267 353 310 615 625 78 78 NOR2_X1 $T=38620 6600 1 0 $X=38505 $Y=5085
X8268 839 310 949 282 78 78 NOR2_X1 $T=39190 29000 0 0 $X=39075 $Y=28885
X8269 284 310 251 599 78 78 NOR2_X1 $T=39380 31800 1 0 $X=39265 $Y=30285
X8270 354 310 288 628 78 78 NOR2_X1 $T=39760 43000 0 0 $X=39645 $Y=42885
X8271 251 310 286 362 78 78 NOR2_X1 $T=39950 31800 0 0 $X=39835 $Y=31685
X8272 604 310 294 660 78 78 NOR2_X1 $T=42230 43000 1 0 $X=42115 $Y=41485
X8287 603 271 272 273 78 310 949 OR4_X1 $T=37670 31800 1 0 $X=37555 $Y=30285
X8288 368 296 295 293 78 310 839 OR4_X1 $T=43370 29000 0 180 $X=42115 $Y=27485
X8289 415 78 310 851 687 36 11 32 851 ICV_26 $T=4040 31800 0 0 $X=3925 $Y=31685
X8290 722 78 310 906 717 399 722 B[31] 466 ICV_26 $T=9550 9400 0 0 $X=9435 $Y=9285
X8291 452 78 310 454 439 A[31] 58 551 454 ICV_26 $T=11450 26200 0 0 $X=11335 $Y=26085
X8292 449 78 310 736 456 399 462 B[31] 449 ICV_26 $T=12970 3800 1 0 $X=12855 $Y=2285
X8293 A[15] 78 310 474 5 469 466 474 78 ICV_26 $T=12970 34600 1 0 $X=12855 $Y=33085
X8294 A[31] 78 310 551 471 A[31] 480 551 934 ICV_26 $T=14680 23400 1 0 $X=14565 $Y=21885
X8295 866 78 310 92 491 399 490 B[31] 92 ICV_26 $T=17340 3800 1 0 $X=17225 $Y=2285
X8296 508 78 310 751 499 A[31] 502 551 751 ICV_26 $T=19050 29000 1 0 $X=18935 $Y=27485
X8297 748 78 310 518 755 A[31] 521 551 518 ICV_26 $T=20760 29000 0 0 $X=20645 $Y=28885
X8298 544 78 310 777 537 399 544 B[31] 169 ICV_26 $T=25700 29000 1 0 $X=25585 $Y=27485
X8299 B[26] 78 310 216 779 198 539 216 562 ICV_26 $T=28360 43000 1 0 $X=28245 $Y=41485
X8300 B[23] 78 310 578 5 578 587 568 355 ICV_26 $T=29880 34600 0 0 $X=29765 $Y=34485
X8301 835 78 310 646 361 242 835 250 353 ICV_26 $T=40520 9400 0 0 $X=40405 $Y=9285
X8302 635 78 310 892 361 234 638 250 255 ICV_26 $T=40520 12200 0 0 $X=40405 $Y=12085
X8303 833 78 310 636 269 636 831 278 614 ICV_26 $T=40520 17800 1 0 $X=40405 $Y=16285
X8304 224 78 310 616 642 616 SUM[3] 194 340 ICV_26 $T=42230 23400 0 0 $X=42115 $Y=23285
X8305 703 78 310 421 694 A[31] 424 551 421 ICV_27 $T=6320 17800 0 0 $X=6205 $Y=17685
X8306 699 78 310 708 314 A[31] 707 551 708 ICV_27 $T=6700 23400 0 0 $X=6585 $Y=23285
X8307 36 78 310 32 45 32 323 36 321 ICV_27 $T=10500 34600 1 0 $X=10385 $Y=33085
X8308 443 78 310 728 730 A[31] 733 551 728 ICV_27 $T=12210 23400 0 0 $X=12095 $Y=23285
X8309 976 78 310 455 463 399 470 B[31] 455 ICV_27 $T=12970 12200 1 0 $X=12855 $Y=10685
X8310 324 78 310 933 479 36 115 32 740 ICV_27 $T=15440 37400 0 0 $X=15325 $Y=37285
X8311 744 78 310 746 483 A[31] 494 551 746 ICV_27 $T=17340 26200 0 0 $X=17225 $Y=26085
X8312 297 78 310 597 218 205 255 602 607 ICV_27 $T=35390 15000 1 0 $X=35275 $Y=13485
X8313 B[29] 78 310 814 5 814 287 809 355 ICV_27 $T=36340 37400 0 0 $X=36225 $Y=37285
X8314 828 78 310 840 836 648 300 254 840 ICV_27 $T=42230 6600 0 0 $X=42115 $Y=6485
X8379 404 405 78 407 36 383 310 851 36 13 32 416 ICV_32 $T=4040 31800 1 0 $X=3925 $Y=30285
X8380 704 36 78 902 32 39 310 687 32 12 36 719 ICV_32 $T=6320 31800 0 0 $X=6205 $Y=31685
X8381 705 696 78 434 666 48 310 317 696 724 46 48 ICV_32 $T=6320 40200 0 0 $X=6205 $Y=40085
X8382 45 36 78 715 32 704 310 719 32 44 36 319 ICV_32 $T=8980 31800 0 0 $X=8865 $Y=31685
X8383 504 A[31] 78 538 551 942 310 503 A[31] 535 551 944 ICV_32 $T=23800 34600 1 0 $X=23685 $Y=33085
X8384 800 237 78 803 254 230 310 806 254 232 237 821 ICV_32 $T=34440 3800 0 0 $X=34325 $Y=3685
X8385 809 B[29] 78 252 B[28] 249 310 779 249 354 887 562 ICV_32 $T=35960 40200 0 0 $X=35845 $Y=40085
X8386 779 809 78 604 814 562 310 5 887 613 249 355 ICV_32 $T=36150 40200 1 0 $X=36035 $Y=38685
X8387 963 269 78 634 221 825 310 269 614 640 194 825 ICV_32 $T=39950 20600 1 0 $X=39835 $Y=19085
X8388 624 229 78 642 280 358 310 358 229 645 280 634 ICV_32 $T=40900 23400 1 0 $X=40785 $Y=21885
X8389 640 229 78 652 280 632 310 632 229 968 280 831 ICV_32 $T=41850 17800 0 0 $X=41735 $Y=17685
X8398 41 16 406 973 310 78 526 FA_X1 $T=5940 9400 1 180 $X=2785 $Y=9285
X8399 16 23 425 849 310 78 752 FA_X1 $T=4990 12200 1 0 $X=4875 $Y=10685
X8400 23 27 707 850 310 78 756 FA_X1 $T=5370 12200 0 0 $X=5255 $Y=12085
X8401 698 34 431 904 310 78 127 FA_X1 $T=5940 3800 1 0 $X=5825 $Y=2285
X8402 34 37 424 930 310 78 118 FA_X1 $T=6130 3800 0 0 $X=6015 $Y=3685
X8403 47 41 688 906 310 78 761 FA_X1 $T=6890 9400 1 0 $X=6775 $Y=7885
X8404 37 47 683 706 310 78 754 FA_X1 $T=7650 6600 0 0 $X=7535 $Y=6485
X8405 27 49 56 907 310 78 525 FA_X1 $T=8030 15000 0 0 $X=7915 $Y=14885
X8406 49 53 58 59 310 78 749 FA_X1 $T=8790 17800 1 0 $X=8675 $Y=16285
X8407 98 698 718 734 310 78 527 FA_X1 $T=9170 3800 0 0 $X=9055 $Y=3685
X8408 53 94 480 910 310 78 119 FA_X1 $T=15060 17800 1 0 $X=14945 $Y=16285
X8409 101 98 733 743 310 78 768 FA_X1 $T=16010 3800 0 0 $X=15895 $Y=3685
X8410 863 99 497 488 310 78 143 FA_X1 $T=16390 9400 1 0 $X=16275 $Y=7885
X8411 981 100 867 B[31] 310 78 328 FA_X1 $T=16770 15000 1 0 $X=16655 $Y=13485
X8412 99 101 113 737 310 78 141 FA_X1 $T=16960 6600 0 0 $X=16845 $Y=6485
X8413 145 102 267 913 310 78 868 FA_X1 $T=16960 43000 0 0 $X=16845 $Y=42885
X8414 492 863 936 485 310 78 528 FA_X1 $T=17340 9400 0 0 $X=17225 $Y=9285
X8415 100 492 867 B[31] 310 78 148 FA_X1 $T=17340 12200 0 0 $X=17225 $Y=12085
X8416 94 109 750 974 310 78 117 FA_X1 $T=17720 17800 0 0 $X=17605 $Y=17685
X8417 109 939 494 914 310 78 146 FA_X1 $T=18480 20600 1 0 $X=18365 $Y=19085
X8418 939 125 502 510 310 78 156 FA_X1 $T=21900 23400 1 180 $X=18745 $Y=23285
X8419 102 126 240 911 310 78 430 FA_X1 $T=21900 40200 1 180 $X=18745 $Y=40085
X8420 125 120 521 765 310 78 155 FA_X1 $T=20000 26200 1 0 $X=19885 $Y=24685
X8421 126 133 248 540 310 78 36 FA_X1 $T=20950 40200 1 0 $X=20835 $Y=38685
X8422 133 149 587 78 310 78 52 FA_X1 $T=25320 37400 1 180 $X=22165 $Y=37285
X8423 120 139 524 915 310 78 174 FA_X1 $T=22660 29000 1 0 $X=22545 $Y=27485
X8424 289 145 276 916 310 78 77 FA_X1 $T=23610 43000 0 0 $X=23495 $Y=42885
X8425 151 943 538 548 310 78 582 FA_X1 $T=23800 31800 1 0 $X=23685 $Y=30285
X8426 139 151 775 777 310 78 184 FA_X1 $T=24180 29000 0 0 $X=24065 $Y=28885
X8427 943 159 535 784 310 78 197 FA_X1 $T=25130 31800 0 0 $X=25015 $Y=31685
X8428 159 170 130 78 310 78 201 FA_X1 $T=26840 34600 0 0 $X=26725 $Y=34485
X8429 235 954 240 924 310 78 804 FA_X1 $T=32160 31800 0 0 $X=32045 $Y=31685
X8430 954 955 248 244 310 78 884 FA_X1 $T=33110 29000 0 0 $X=32995 $Y=28885
X8431 258 235 256 267 310 78 885 FA_X1 $T=33490 34600 1 0 $X=33375 $Y=33085
X8432 279 258 617 257 310 78 605 FA_X1 $T=35580 29000 1 0 $X=35465 $Y=27485
X8433 281 279 639 889 310 78 891 FA_X1 $T=38620 29000 1 0 $X=38505 $Y=27485
X8434 633 281 952 362 310 78 893 FA_X1 $T=38810 34600 1 0 $X=38695 $Y=33085
X8435 303 289 613 926 310 78 371 FA_X1 $T=41850 43000 0 180 $X=38695 $Y=41485
X8436 982 78 307 927 310 78 364 FA_X1 $T=44700 37400 0 180 $X=41545 $Y=35885
X8437 78 303 287 928 310 78 369 FA_X1 $T=44700 40200 1 180 $X=41545 $Y=40085
X8438 355 B[17] 310 A[17] 391 5 78 996 AOI22_X1 $T=1000 1000 0 0 $X=885 $Y=885
X8439 355 B[16] 310 A[16] 675 5 78 78 AOI22_X1 $T=1000 3800 0 0 $X=885 $Y=3685
X8440 355 B[14] 310 A[14] 389 5 78 78 AOI22_X1 $T=1000 6600 1 0 $X=885 $Y=5085
X8441 355 B[12] 310 A[12] 896 5 78 78 AOI22_X1 $T=1000 12200 1 0 $X=885 $Y=10685
X8442 355 B[11] 310 A[11] 390 5 78 78 AOI22_X1 $T=1000 17800 1 0 $X=885 $Y=16285
X8443 78 A[20] 310 B[20] 405 5 78 78 AOI22_X1 $T=1000 34600 0 0 $X=885 $Y=34485
X8444 78 A[14] 310 B[14] 313 5 78 78 AOI22_X1 $T=1000 37400 1 0 $X=885 $Y=35885
X8445 78 A[16] 310 B[16] 64 5 78 78 AOI22_X1 $T=1000 37400 0 0 $X=885 $Y=37285
X8446 78 A[13] 310 B[13] 312 5 78 78 AOI22_X1 $T=1000 40200 1 0 $X=885 $Y=38685
X8447 78 A[18] 310 B[18] 666 5 78 78 AOI22_X1 $T=1000 40200 0 0 $X=885 $Y=40085
X8448 78 A[10] 310 B[10] 705 5 78 78 AOI22_X1 $T=1000 43000 0 0 $X=885 $Y=42885
X8449 355 B[18] 310 A[18] 677 5 78 996 AOI22_X1 $T=1950 1000 0 0 $X=1835 $Y=885
X8450 355 B[13] 310 A[13] 847 5 78 78 AOI22_X1 $T=2140 9400 1 0 $X=2025 $Y=7885
X8451 78 A[22] 310 B[22] 38 5 78 78 AOI22_X1 $T=2330 34600 0 0 $X=2215 $Y=34485
X8452 78 A[12] 310 B[12] 24 5 78 78 AOI22_X1 $T=2330 40200 1 0 $X=2215 $Y=38685
X8453 355 B[10] 310 A[10] 411 5 78 78 AOI22_X1 $T=4230 17800 1 0 $X=4115 $Y=16285
X8454 78 A[17] 310 B[17] 46 5 78 78 AOI22_X1 $T=4800 43000 0 0 $X=4685 $Y=42885
X8455 14 430 310 18 45 434 78 78 AOI22_X1 $T=7650 37400 1 0 $X=7535 $Y=35885
X8456 434 430 310 18 857 697 78 78 AOI22_X1 $T=7840 37400 0 0 $X=7725 $Y=37285
X8457 697 430 310 18 479 417 78 78 AOI22_X1 $T=8220 40200 1 0 $X=8105 $Y=38685
X8458 78 A[9] 310 B[9] 317 33 78 78 AOI22_X1 $T=8600 43000 0 0 $X=8485 $Y=42885
X8459 724 18 310 430 731 318 78 78 AOI22_X1 $T=9550 37400 1 0 $X=9435 $Y=35885
X8460 78 A[19] 310 B[19] 721 33 78 78 AOI22_X1 $T=9550 43000 0 0 $X=9435 $Y=42885
X8461 859 430 310 18 687 459 78 78 AOI22_X1 $T=9740 34600 0 0 $X=9625 $Y=34485
X8462 700 18 310 430 860 724 78 78 AOI22_X1 $T=9930 40200 0 0 $X=9815 $Y=40085
X8463 355 B[19] 310 A[19] 320 5 78 996 AOI22_X1 $T=10500 1000 0 0 $X=10385 $Y=885
X8464 355 B[8] 310 A[8] 446 5 78 78 AOI22_X1 $T=10500 12200 0 0 $X=10385 $Y=12085
X8465 78 A[8] 310 B[8] 723 33 78 78 AOI22_X1 $T=10690 43000 1 0 $X=10575 $Y=41485
X8466 355 B[22] 310 A[22] 976 5 78 78 AOI22_X1 $T=11070 12200 1 0 $X=10955 $Y=10685
X8467 355 B[9] 310 A[9] 727 5 78 78 AOI22_X1 $T=11450 12200 0 0 $X=11335 $Y=12085
X8468 725 18 310 430 321 322 78 78 AOI22_X1 $T=11450 37400 1 0 $X=11335 $Y=35885
X8469 459 430 310 18 319 80 78 78 AOI22_X1 $T=11640 34600 0 0 $X=11525 $Y=34485
X8470 78 A[11] 310 B[11] 71 33 78 78 AOI22_X1 $T=12970 43000 0 0 $X=12855 $Y=42885
X8471 66 18 310 430 740 725 78 78 AOI22_X1 $T=13160 37400 0 0 $X=13045 $Y=37285
X8472 62 551 310 A[31] 473 477 78 78 AOI22_X1 $T=13730 23400 1 0 $X=13615 $Y=21885
X8473 933 430 310 18 738 461 78 78 AOI22_X1 $T=14300 40200 0 0 $X=14185 $Y=40085
X8474 731 36 310 32 89 478 78 78 AOI22_X1 $T=14490 31800 0 0 $X=14375 $Y=31685
X8475 860 32 310 36 862 478 78 78 AOI22_X1 $T=15440 34600 1 0 $X=15325 $Y=33085
X8476 738 36 310 32 742 716 78 78 AOI22_X1 $T=16580 40200 0 0 $X=16465 $Y=40085
X8477 355 B[20] 310 A[20] 866 5 78 996 AOI22_X1 $T=18290 1000 0 0 $X=18175 $Y=885
X8478 355 B[5] 310 A[5] 762 5 78 78 AOI22_X1 $T=21900 20600 1 0 $X=21785 $Y=19085
X8479 869 SUM[31] 310 165 297 119 78 78 AOI22_X1 $T=22660 15000 0 0 $X=22545 $Y=14885
X8480 355 B[6] 310 A[6] 766 5 78 78 AOI22_X1 $T=22850 20600 1 0 $X=22735 $Y=19085
X8481 355 B[4] 310 A[4] 542 5 78 78 AOI22_X1 $T=26080 23400 0 0 $X=25965 $Y=23285
X8482 A[31] 399 310 B[31] 356 551 78 78 AOI22_X1 $T=26840 26200 1 0 $X=26725 $Y=24685
X8483 355 B[3] 310 A[3] 918 5 78 78 AOI22_X1 $T=27790 26200 1 0 $X=27675 $Y=24685
X8484 355 B[0] 310 A[0] 191 5 78 78 AOI22_X1 $T=30260 34600 1 0 $X=30145 $Y=33085
X8485 355 B[1] 310 A[1] 787 5 78 78 AOI22_X1 $T=30640 29000 0 0 $X=30525 $Y=28885
X8486 355 B[2] 310 A[2] 792 5 78 78 AOI22_X1 $T=30830 29000 1 0 $X=30715 $Y=27485
X8487 881 SUM[31] 310 165 259 582 78 78 AOI22_X1 $T=31020 26200 1 0 $X=30905 $Y=24685
X8488 581 SUM[31] 310 165 221 184 78 78 AOI22_X1 $T=31970 23400 0 0 $X=31855 $Y=23285
X8489 874 587 310 797 296 229 78 78 AOI22_X1 $T=33490 26200 0 0 $X=33375 $Y=26085
X8490 880 977 310 B[28] 810 249 78 78 AOI22_X1 $T=33490 43000 0 0 $X=33375 $Y=42885
X8491 277 250 310 265 806 590 78 78 AOI22_X1 $T=34060 6600 0 0 $X=33945 $Y=6485
X8492 592 SUM[31] 310 165 247 197 78 78 AOI22_X1 $T=34250 26200 1 0 $X=34135 $Y=24685
X8493 284 807 310 884 273 599 78 78 AOI22_X1 $T=35200 31800 1 0 $X=35085 $Y=30285
X8494 284 808 310 804 272 599 78 78 AOI22_X1 $T=35200 31800 0 0 $X=35085 $Y=31685
X8495 241 602 310 822 813 280 78 78 AOI22_X1 $T=35960 20600 1 0 $X=35845 $Y=19085
X8496 284 621 310 605 603 599 78 78 AOI22_X1 $T=36150 29000 0 0 $X=36035 $Y=28885
X8497 284 815 310 885 271 599 78 78 AOI22_X1 $T=36530 34600 1 0 $X=36415 $Y=33085
X8498 809 B[29] 310 B[30] 598 360 78 78 AOI22_X1 $T=36910 43000 1 0 $X=36795 $Y=41485
X8499 250 602 310 243 614 265 78 78 AOI22_X1 $T=37290 17800 1 0 $X=37175 $Y=16285
X8500 250 822 310 609 963 265 78 78 AOI22_X1 $T=38240 17800 1 0 $X=38125 $Y=16285
X8501 629 254 310 237 283 829 78 78 AOI22_X1 $T=39380 3800 0 0 $X=39265 $Y=3685
X8502 250 359 310 346 292 265 78 78 AOI22_X1 $T=39760 15000 0 0 $X=39645 $Y=14885
X8503 284 834 310 891 293 599 78 78 AOI22_X1 $T=40900 31800 1 0 $X=40785 $Y=30285
X8504 284 838 310 893 295 599 78 78 AOI22_X1 $T=41660 31800 0 0 $X=41545 $Y=31685
X8584 808 593 240 78 310 883 HA_X1 $T=33490 37400 1 0 $X=33375 $Y=35885
X8585 807 587 248 78 310 593 HA_X1 $T=34250 34600 0 0 $X=34135 $Y=34485
X8586 815 883 267 78 310 824 HA_X1 $T=36150 34600 0 0 $X=36035 $Y=34485
X8587 617 276 275 78 310 889 HA_X1 $T=37670 26200 0 0 $X=37555 $Y=26085
X8588 621 824 276 78 310 890 HA_X1 $T=38050 34600 0 0 $X=37935 $Y=34485
X8589 838 950 287 78 310 837 HA_X1 $T=39950 37400 0 0 $X=39835 $Y=37285
X8590 834 890 613 78 310 950 HA_X1 $T=41850 40200 0 180 $X=39835 $Y=38685
X8591 251 229 874 78 310 NOR2_X2 $T=35200 26200 1 0 $X=35085 $Y=24685
X8592 284 224 285 78 310 NOR2_X2 $T=39570 26200 0 0 $X=39455 $Y=26085
X8625 78 310 714 904 996 ICV_41 $T=8980 1000 0 0 $X=8865 $Y=885
X8626 78 310 429 431 78 ICV_41 $T=9550 12200 1 0 $X=9435 $Y=10685
X8627 78 310 483 90 78 ICV_41 $T=16200 29000 0 0 $X=16085 $Y=28885
X8628 78 310 489 936 78 ICV_41 $T=18480 17800 1 0 $X=18365 $Y=16285
X8629 78 310 753 941 78 ICV_41 $T=22660 34600 1 0 $X=22545 $Y=33085
X8630 78 310 770 944 78 ICV_41 $T=25130 34600 0 0 $X=25015 $Y=34485
X8631 78 310 780 877 78 ICV_41 $T=29310 3800 0 0 $X=29195 $Y=3685
X8632 78 310 210 798 78 ICV_41 $T=33490 17800 0 0 $X=33375 $Y=17685
X8633 78 310 B[25] 794 78 ICV_41 $T=33680 37400 0 0 $X=33565 $Y=37285
X8634 78 310 A[28] 249 78 ICV_41 $T=34630 40200 1 0 $X=34515 $Y=38685
X8635 78 310 274 609 78 ICV_41 $T=38620 15000 1 0 $X=38505 $Y=13485
X8636 78 310 221 359 78 ICV_41 $T=38620 15000 0 0 $X=38505 $Y=14885
X8637 182 78 202 199 310 189 NAND3_X1 $T=28740 12200 1 0 $X=28625 $Y=10685
X8638 561 78 180 780 310 196 NAND3_X1 $T=28740 15000 1 0 $X=28625 $Y=13485
X8639 789 78 242 297 310 575 NAND3_X1 $T=30830 15000 0 0 $X=30715 $Y=14885
X8640 254 78 607 275 310 278 NAND3_X1 $T=38240 12200 0 0 $X=38125 $Y=12085
X8641 237 78 607 275 310 269 NAND3_X1 $T=38240 17800 0 0 $X=38125 $Y=17685
X8671 282 356 618 78 811 285 247 SUM[0] 310 OAI33_X1 $T=37670 26200 1 0 $X=37555 $Y=24685
X8672 616 813 622 78 811 285 259 SUM[1] 310 OAI33_X1 $T=37860 23400 0 0 $X=37745 $Y=23285
X8724 348 140 78 221 231 233 310 220 261 OAI222_X1 $T=33110 12200 1 0 $X=32995 $Y=10685
X8725 348 297 78 247 231 233 310 253 268 OAI222_X1 $T=34630 12200 1 0 $X=34515 $Y=10685
X8726 348 291 78 259 231 233 310 266 816 OAI222_X1 $T=35770 12200 0 0 $X=35655 $Y=12085
X8727 260 310 238 250 924 78 AOI21_X2 $T=33490 23400 1 0 $X=33375 $Y=21885
X8728 610 310 260 607 256 78 AOI21_X2 $T=35580 20600 0 0 $X=35465 $Y=20485
X8729 394 78 310 376 403 383 ICV_47 $T=1760 31800 0 0 $X=1645 $Y=31685
X8730 435 78 310 931 432 710 ICV_47 $T=9360 26200 1 0 $X=9245 $Y=24685
X8731 727 78 310 75 465 497 ICV_47 $T=13920 12200 0 0 $X=13805 $Y=12085
X8732 471 78 310 83 481 81 ICV_47 $T=15060 26200 0 0 $X=14945 $Y=26085
X8733 873 78 310 153 773 160 ICV_47 $T=25890 40200 0 0 $X=25775 $Y=40085
X8734 A[24] 78 310 552 B[24] 213 ICV_47 $T=26840 37400 1 0 $X=26725 $Y=35885
X8735 A[27] 78 310 217 558 288 ICV_47 $T=32730 43000 0 0 $X=32615 $Y=42885
X8736 779 78 310 562 A[29] 809 ICV_47 $T=34820 37400 0 0 $X=34705 $Y=37285
X8741 13 63 78 673 1 2 310 52 78 ICV_48 $T=1000 26200 0 0 $X=885 $Y=26085
X8742 78 B[5] 78 25 3 5 310 A[5] 78 ICV_48 $T=1950 40200 0 0 $X=1835 $Y=40085
X8743 78 B[4] 78 20 3 5 310 A[4] 78 ICV_48 $T=2330 43000 1 0 $X=2215 $Y=41485
X8744 19 721 78 461 68 71 310 48 78 ICV_48 $T=12400 43000 1 0 $X=12285 $Y=41485
X8745 862 52 78 755 1 96 310 63 78 ICV_48 $T=16580 31800 0 0 $X=16465 $Y=31685
X8746 A[24] 213 78 195 186 A[25] 310 794 78 ICV_48 $T=28740 40200 1 0 $X=28625 $Y=38685
X8747 803 280 78 788 224 232 310 229 996 ICV_48 $T=33490 1000 0 0 $X=33375 $Y=885
X8748 231 234 78 802 237 239 310 589 78 ICV_48 $T=33870 9400 0 0 $X=33755 $Y=9285
X8749 681 310 381 311 78 9 NOR3_X1 $T=2330 23400 0 0 $X=2215 $Y=23285
X8750 395 310 397 844 78 30 NOR3_X1 $T=3470 9400 1 0 $X=3355 $Y=7885
X8751 410 310 412 414 78 72 NOR3_X1 $T=5180 3800 1 0 $X=5065 $Y=2285
X8752 455 310 442 468 78 93 NOR3_X1 $T=13730 9400 1 0 $X=13615 $Y=7885
X8753 752 310 756 758 78 136 NOR3_X1 $T=20380 9400 0 0 $X=20265 $Y=9285
X8754 768 310 527 142 78 172 NOR3_X1 $T=23800 3800 1 0 $X=23685 $Y=2285
X8755 148 310 528 532 78 162 NOR3_X1 $T=24560 12200 1 0 $X=24445 $Y=10685
X8756 585 310 243 346 78 586 NOR3_X1 $T=33300 17800 1 0 $X=33185 $Y=16285
X8757 798 310 822 201 78 972 NOR3_X1 $T=33490 20600 1 0 $X=33375 $Y=19085
X8758 422 52 1 310 54 730 78 OAI211_X1 $T=8600 29000 1 0 $X=8485 $Y=27485
X8759 479 32 63 310 95 861 78 OAI211_X1 $T=14870 40200 1 0 $X=14755 $Y=38685
X8760 742 63 1 310 861 865 78 OAI211_X1 $T=18860 40200 1 180 $X=17795 $Y=40085
X8761 552 B[24] B[23] 310 568 186 78 OAI211_X1 $T=28550 37400 1 0 $X=28435 $Y=35885
X8762 A[24] 213 578 310 A[23] 219 78 OAI211_X1 $T=31590 37400 0 0 $X=31475 $Y=37285
X8763 226 229 224 310 236 580 78 OAI211_X1 $T=33490 3800 0 0 $X=33375 $Y=3685
X8764 61 51 78 310 55 AND2_X1 $T=8600 20600 0 0 $X=8485 $Y=20485
X8765 1 57 78 310 440 AND2_X1 $T=9930 31800 1 0 $X=9815 $Y=30285
X8766 84 65 78 310 477 AND2_X1 $T=12210 20600 0 0 $X=12095 $Y=20485
X8767 732 70 78 310 464 AND2_X1 $T=12780 15000 0 0 $X=12665 $Y=14885
X8768 450 85 78 310 739 AND2_X1 $T=14490 23400 0 0 $X=14375 $Y=23285
X8769 108 87 78 310 486 AND2_X1 $T=15060 20600 0 0 $X=14945 $Y=20485
X8770 A[31] 108 78 310 867 AND2_X1 $T=18100 15000 0 0 $X=17985 $Y=14885
X8771 88 111 78 310 508 AND2_X1 $T=18290 29000 1 0 $X=18175 $Y=27485
X8772 513 128 78 310 869 AND2_X1 $T=21140 17800 1 0 $X=21025 $Y=16285
X8773 516 131 78 310 520 AND2_X1 $T=21900 23400 0 180 $X=21025 $Y=21885
X8774 509 132 78 310 514 AND2_X1 $T=21900 34600 1 180 $X=21025 $Y=34485
X8775 152 150 78 310 534 AND2_X1 $T=24560 3800 0 0 $X=24445 $Y=3685
X8776 532 157 78 310 771 AND2_X1 $T=25320 6600 0 0 $X=25205 $Y=6485
X8777 772 163 78 310 774 AND2_X1 $T=25890 20600 0 0 $X=25775 $Y=20485
X8778 208 167 78 310 561 AND2_X1 $T=27030 6600 0 0 $X=26915 $Y=6485
X8779 557 176 78 310 778 AND2_X1 $T=27980 29000 1 0 $X=27865 $Y=27485
X8780 336 207 78 310 881 AND2_X1 $T=31020 26200 0 0 $X=30905 $Y=26085
X8781 40 42 43 78 310 61 OR3_X1 $T=7650 20600 0 0 $X=7535 $Y=20485
X8782 61 60 62 78 310 84 OR3_X1 $T=11260 20600 0 0 $X=11145 $Y=20485
X8783 74 73 75 78 310 732 OR3_X1 $T=13160 15000 1 0 $X=13045 $Y=13485
X8784 84 79 82 78 310 108 OR3_X1 $T=13920 20600 1 0 $X=13805 $Y=19085
X8785 86 81 83 78 310 450 OR3_X1 $T=14110 26200 1 0 $X=13995 $Y=24685
X8786 106 103 104 78 310 88 OR3_X1 $T=17530 31800 1 0 $X=17415 $Y=30285
X8787 124 117 119 78 310 513 OR3_X1 $T=20190 17800 1 0 $X=20075 $Y=16285
X8788 511 121 130 78 310 509 OR3_X1 $T=20950 37400 1 0 $X=20835 $Y=35885
X8789 129 137 135 78 310 516 OR3_X1 $T=23230 20600 1 180 $X=22165 $Y=20485
X8790 152 141 143 78 310 532 OR3_X1 $T=23800 6600 1 0 $X=23685 $Y=5085
X8791 161 155 156 78 310 772 OR3_X1 $T=24940 20600 0 0 $X=24825 $Y=20485
X8792 563 185 170 78 310 557 OR3_X1 $T=29500 29000 1 0 $X=29385 $Y=27485
X8793 582 197 201 78 310 336 OR3_X1 $T=30070 26200 1 0 $X=29955 $Y=24685
X8794 427 551 78 429 A[31] 42 310 42 427 40 78 ICV_49 $T=6510 20600 1 0 $X=6395 $Y=19085
X8795 458 551 78 465 A[31] 79 310 79 458 84 78 ICV_49 $T=11830 20600 1 0 $X=11715 $Y=19085
X8796 457 399 78 467 B[31] 442 310 442 457 468 78 ICV_49 $T=12020 6600 0 0 $X=11905 $Y=6485
X8797 741 399 78 105 B[31] 73 310 73 741 74 78 ICV_49 $T=16010 15000 0 0 $X=15895 $Y=14885
X8798 493 399 78 496 B[31] 107 310 107 493 516 78 ICV_49 $T=16770 23400 1 0 $X=16655 $Y=21885
X8799 749 SUM[31] 78 291 165 759 310 749 759 513 78 ICV_49 $T=20570 15000 0 0 $X=20455 $Y=14885
X8800 117 SUM[31] 78 242 165 523 310 117 523 124 78 ICV_49 $T=22470 17800 0 0 $X=22355 $Y=17685
X8801 527 SUM[31] 78 220 165 530 310 527 530 142 996 ICV_49 $T=23230 1000 0 0 $X=23115 $Y=885
X8802 528 SUM[31] 78 208 165 536 310 528 536 532 78 ICV_49 $T=24560 9400 1 0 $X=24445 $Y=7885
X8803 146 SUM[31] 78 227 165 545 310 146 545 772 78 ICV_49 $T=24940 20600 1 0 $X=24825 $Y=19085
X8804 155 SUM[31] 78 274 165 560 310 155 560 161 78 ICV_49 $T=27600 20600 0 0 $X=27485 $Y=20485
X8805 567 399 78 571 B[31] 185 310 185 567 170 78 ICV_49 $T=28550 31800 1 0 $X=28435 $Y=30285
X8806 328 SUM[31] 78 310 CLKBUF_X2 $T=19810 15000 1 0 $X=19695 $Y=13485
X8807 78 355 78 310 CLKBUF_X2 $T=28360 37400 0 0 $X=28245 $Y=37285
X8808 405 32 310 35 38 78 36 422 AOI221_X1 $T=6130 29000 0 0 $X=6015 $Y=28885
X8809 5 469 310 77 78 78 474 67 AOI221_X1 $T=13350 34600 0 0 $X=13235 $Y=34485
.ENDS
***************************************
