/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Dec 17 20:47:37 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 387956002 */

module datapath(p_0, accumulator, p_1);
   input [31:0]p_0;
   input [31:0]accumulator;
   output [31:0]p_1;

   INV_X1 i_0 (.A(n_0), .ZN(p_1[0]));
   OAI21_X1 i_1 (.A(n_159), .B1(p_0[0]), .B2(accumulator[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_159), .B(n_1), .Z(p_1[1]));
   OAI21_X1 i_3 (.A(n_158), .B1(p_0[1]), .B2(accumulator[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_157), .B(n_2), .ZN(p_1[2]));
   OAI21_X1 i_5 (.A(n_162), .B1(p_0[2]), .B2(accumulator[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_156), .B(n_3), .Z(p_1[3]));
   OAI21_X1 i_7 (.A(n_163), .B1(n_168), .B2(n_165), .ZN(n_3));
   XOR2_X1 i_8 (.A(n_154), .B(n_10), .Z(p_1[4]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_1[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_1[6]));
   NOR2_X1 i_11 (.A1(n_151), .A2(n_142), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_1[7]));
   OAI22_X1 i_13 (.A1(p_0[6]), .A2(accumulator[6]), .B1(n_142), .B2(n_7), 
      .ZN(n_5));
   AOI21_X1 i_14 (.A(n_152), .B1(p_0[5]), .B2(accumulator[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_152), .B1(n_146), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_149), .B1(n_154), .B2(n_147), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_147), .B1(p_0[4]), .B2(accumulator[4]), .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_153), .A2(n_144), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_140), .B(n_18), .ZN(p_1[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_1[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_1[10]));
   NOR2_X1 i_23 (.A1(n_137), .A2(n_128), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_1[11]));
   OAI22_X1 i_25 (.A1(p_0[10]), .A2(accumulator[10]), .B1(n_128), .B2(n_15), 
      .ZN(n_13));
   AOI21_X1 i_26 (.A(n_138), .B1(p_0[9]), .B2(accumulator[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_138), .B1(n_132), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_135), .B1(n_140), .B2(n_133), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_135), .B1(p_0[8]), .B2(accumulator[8]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_139), .A2(n_130), .ZN(n_19));
   XOR2_X1 i_32 (.A(n_126), .B(n_26), .Z(p_1[12]));
   XOR2_X1 i_33 (.A(n_25), .B(n_22), .Z(p_1[13]));
   XOR2_X1 i_34 (.A(n_23), .B(n_20), .Z(p_1[14]));
   NOR2_X1 i_35 (.A1(n_123), .A2(n_114), .ZN(n_20));
   XNOR2_X1 i_36 (.A(n_27), .B(n_21), .ZN(p_1[15]));
   OAI22_X1 i_37 (.A1(p_0[14]), .A2(accumulator[14]), .B1(n_114), .B2(n_23), 
      .ZN(n_21));
   AOI21_X1 i_38 (.A(n_124), .B1(p_0[13]), .B2(accumulator[13]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_124), .B1(n_118), .B2(n_24), .ZN(n_23));
   INV_X1 i_40 (.A(n_25), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_121), .B1(n_126), .B2(n_119), .ZN(n_25));
   OAI21_X1 i_42 (.A(n_119), .B1(p_0[12]), .B2(accumulator[12]), .ZN(n_26));
   NOR2_X1 i_43 (.A1(n_125), .A2(n_116), .ZN(n_27));
   XOR2_X1 i_44 (.A(n_112), .B(n_34), .Z(p_1[16]));
   XOR2_X1 i_45 (.A(n_33), .B(n_30), .Z(p_1[17]));
   XOR2_X1 i_46 (.A(n_31), .B(n_28), .Z(p_1[18]));
   NOR2_X1 i_47 (.A1(n_109), .A2(n_100), .ZN(n_28));
   XNOR2_X1 i_48 (.A(n_35), .B(n_29), .ZN(p_1[19]));
   OAI22_X1 i_49 (.A1(p_0[18]), .A2(accumulator[18]), .B1(n_100), .B2(n_31), 
      .ZN(n_29));
   AOI21_X1 i_50 (.A(n_110), .B1(p_0[17]), .B2(accumulator[17]), .ZN(n_30));
   AOI21_X1 i_51 (.A(n_110), .B1(n_104), .B2(n_32), .ZN(n_31));
   INV_X1 i_52 (.A(n_33), .ZN(n_32));
   AOI21_X1 i_53 (.A(n_107), .B1(n_112), .B2(n_105), .ZN(n_33));
   OAI21_X1 i_54 (.A(n_105), .B1(p_0[16]), .B2(accumulator[16]), .ZN(n_34));
   NOR2_X1 i_55 (.A1(n_111), .A2(n_102), .ZN(n_35));
   XOR2_X1 i_56 (.A(n_98), .B(n_42), .Z(p_1[20]));
   XOR2_X1 i_57 (.A(n_41), .B(n_38), .Z(p_1[21]));
   XOR2_X1 i_58 (.A(n_39), .B(n_36), .Z(p_1[22]));
   NOR2_X1 i_59 (.A1(n_87), .A2(n_77), .ZN(n_36));
   XNOR2_X1 i_60 (.A(n_43), .B(n_37), .ZN(p_1[23]));
   OAI21_X1 i_61 (.A(n_86), .B1(n_77), .B2(n_39), .ZN(n_37));
   NOR2_X1 i_62 (.A1(n_89), .A2(n_79), .ZN(n_38));
   INV_X1 i_63 (.A(n_40), .ZN(n_39));
   OAI21_X1 i_64 (.A(n_88), .B1(n_79), .B2(n_41), .ZN(n_40));
   AOI21_X1 i_65 (.A(n_84), .B1(n_98), .B2(n_81), .ZN(n_41));
   OAI21_X1 i_66 (.A(n_81), .B1(p_0[20]), .B2(accumulator[20]), .ZN(n_42));
   AOI21_X1 i_67 (.A(n_91), .B1(p_0[23]), .B2(accumulator[23]), .ZN(n_43));
   XNOR2_X1 i_68 (.A(n_52), .B(n_51), .ZN(p_1[24]));
   XOR2_X1 i_69 (.A(n_49), .B(n_48), .Z(p_1[25]));
   XNOR2_X1 i_70 (.A(n_45), .B(n_44), .ZN(p_1[26]));
   OAI22_X1 i_71 (.A1(p_0[25]), .A2(accumulator[25]), .B1(n_72), .B2(n_49), 
      .ZN(n_44));
   NOR2_X1 i_72 (.A1(n_95), .A2(n_68), .ZN(n_45));
   XNOR2_X1 i_73 (.A(n_53), .B(n_46), .ZN(p_1[27]));
   OAI21_X1 i_74 (.A(n_47), .B1(n_94), .B2(n_68), .ZN(n_46));
   NAND3_X1 i_75 (.A1(n_69), .A2(n_48), .A3(n_50), .ZN(n_47));
   NOR2_X1 i_76 (.A1(n_96), .A2(n_72), .ZN(n_48));
   INV_X1 i_77 (.A(n_50), .ZN(n_49));
   OAI22_X1 i_78 (.A1(p_0[24]), .A2(accumulator[24]), .B1(n_73), .B2(n_52), 
      .ZN(n_50));
   OAI21_X1 i_79 (.A(n_74), .B1(p_0[24]), .B2(accumulator[24]), .ZN(n_51));
   OAI21_X1 i_80 (.A(n_76), .B1(n_98), .B2(n_83), .ZN(n_52));
   AOI21_X1 i_81 (.A(n_97), .B1(p_0[27]), .B2(accumulator[27]), .ZN(n_53));
   XNOR2_X1 i_82 (.A(n_66), .B(n_65), .ZN(p_1[28]));
   AOI22_X1 i_83 (.A1(n_63), .A2(n_59), .B1(n_64), .B2(n_58), .ZN(p_1[29]));
   XOR2_X1 i_84 (.A(n_55), .B(n_54), .Z(p_1[30]));
   AOI22_X1 i_85 (.A1(p_0[29]), .A2(accumulator[29]), .B1(n_64), .B2(n_60), 
      .ZN(n_54));
   OAI21_X1 i_86 (.A(n_62), .B1(p_0[30]), .B2(accumulator[30]), .ZN(n_55));
   XNOR2_X1 i_87 (.A(p_0[31]), .B(n_56), .ZN(p_1[31]));
   OAI221_X1 i_88 (.A(n_57), .B1(p_0[30]), .B2(accumulator[30]), .C1(n_61), 
      .C2(n_60), .ZN(n_56));
   NAND3_X1 i_89 (.A1(n_62), .A2(n_58), .A3(n_63), .ZN(n_57));
   INV_X1 i_90 (.A(n_59), .ZN(n_58));
   OAI21_X1 i_91 (.A(n_60), .B1(n_170), .B2(n_167), .ZN(n_59));
   NAND2_X1 i_92 (.A1(n_170), .A2(n_167), .ZN(n_60));
   INV_X1 i_93 (.A(n_62), .ZN(n_61));
   NAND2_X1 i_94 (.A1(p_0[30]), .A2(accumulator[30]), .ZN(n_62));
   INV_X1 i_95 (.A(n_64), .ZN(n_63));
   AOI21_X1 i_96 (.A(n_164), .B1(n_66), .B2(n_65), .ZN(n_64));
   AOI21_X1 i_97 (.A(n_164), .B1(p_0[28]), .B2(accumulator[28]), .ZN(n_65));
   NOR4_X1 i_98 (.A1(n_70), .A2(n_67), .A3(n_75), .A4(n_82), .ZN(n_66));
   OAI22_X1 i_99 (.A1(n_169), .A2(n_166), .B1(n_97), .B2(n_69), .ZN(n_67));
   INV_X1 i_100 (.A(n_69), .ZN(n_68));
   NAND2_X1 i_101 (.A1(p_0[26]), .A2(accumulator[26]), .ZN(n_69));
   INV_X1 i_102 (.A(n_71), .ZN(n_70));
   OAI21_X1 i_103 (.A(n_93), .B1(n_73), .B2(n_72), .ZN(n_71));
   AND2_X1 i_104 (.A1(p_0[25]), .A2(accumulator[25]), .ZN(n_72));
   INV_X1 i_105 (.A(n_74), .ZN(n_73));
   NAND2_X1 i_106 (.A1(p_0[24]), .A2(accumulator[24]), .ZN(n_74));
   NOR2_X1 i_107 (.A1(n_92), .A2(n_76), .ZN(n_75));
   AOI221_X1 i_108 (.A(n_78), .B1(p_0[23]), .B2(accumulator[23]), .C1(n_90), 
      .C2(n_77), .ZN(n_76));
   AND2_X1 i_109 (.A1(p_0[22]), .A2(accumulator[22]), .ZN(n_77));
   AOI21_X1 i_110 (.A(n_85), .B1(n_81), .B2(n_80), .ZN(n_78));
   INV_X1 i_111 (.A(n_80), .ZN(n_79));
   NAND2_X1 i_112 (.A1(p_0[21]), .A2(accumulator[21]), .ZN(n_80));
   NAND2_X1 i_113 (.A1(p_0[20]), .A2(accumulator[20]), .ZN(n_81));
   NOR3_X1 i_114 (.A1(n_92), .A2(n_83), .A3(n_98), .ZN(n_82));
   OR2_X1 i_115 (.A1(n_85), .A2(n_84), .ZN(n_83));
   NOR2_X1 i_116 (.A1(p_0[20]), .A2(accumulator[20]), .ZN(n_84));
   NAND3_X1 i_117 (.A1(n_90), .A2(n_86), .A3(n_88), .ZN(n_85));
   INV_X1 i_118 (.A(n_87), .ZN(n_86));
   NOR2_X1 i_119 (.A1(p_0[22]), .A2(accumulator[22]), .ZN(n_87));
   INV_X1 i_120 (.A(n_89), .ZN(n_88));
   NOR2_X1 i_121 (.A1(p_0[21]), .A2(accumulator[21]), .ZN(n_89));
   INV_X1 i_122 (.A(n_91), .ZN(n_90));
   NOR2_X1 i_123 (.A1(p_0[23]), .A2(accumulator[23]), .ZN(n_91));
   OAI21_X1 i_124 (.A(n_93), .B1(p_0[24]), .B2(accumulator[24]), .ZN(n_92));
   NOR3_X1 i_125 (.A1(n_97), .A2(n_95), .A3(n_96), .ZN(n_93));
   NOR2_X1 i_126 (.A1(n_96), .A2(n_95), .ZN(n_94));
   NOR2_X1 i_127 (.A1(p_0[26]), .A2(accumulator[26]), .ZN(n_95));
   NOR2_X1 i_128 (.A1(p_0[25]), .A2(accumulator[25]), .ZN(n_96));
   NOR2_X1 i_129 (.A1(p_0[27]), .A2(accumulator[27]), .ZN(n_97));
   NOR4_X1 i_130 (.A1(n_102), .A2(n_99), .A3(n_103), .A4(n_106), .ZN(n_98));
   NOR2_X1 i_131 (.A1(n_111), .A2(n_101), .ZN(n_99));
   INV_X1 i_132 (.A(n_101), .ZN(n_100));
   NAND2_X1 i_133 (.A1(p_0[18]), .A2(accumulator[18]), .ZN(n_101));
   AND2_X1 i_134 (.A1(p_0[19]), .A2(accumulator[19]), .ZN(n_102));
   AOI21_X1 i_135 (.A(n_108), .B1(n_105), .B2(n_104), .ZN(n_103));
   NAND2_X1 i_136 (.A1(p_0[17]), .A2(accumulator[17]), .ZN(n_104));
   NAND2_X1 i_137 (.A1(p_0[16]), .A2(accumulator[16]), .ZN(n_105));
   NOR3_X1 i_138 (.A1(n_108), .A2(n_107), .A3(n_112), .ZN(n_106));
   NOR2_X1 i_139 (.A1(p_0[16]), .A2(accumulator[16]), .ZN(n_107));
   OR3_X1 i_140 (.A1(n_111), .A2(n_109), .A3(n_110), .ZN(n_108));
   NOR2_X1 i_141 (.A1(p_0[18]), .A2(accumulator[18]), .ZN(n_109));
   NOR2_X1 i_142 (.A1(p_0[17]), .A2(accumulator[17]), .ZN(n_110));
   NOR2_X1 i_143 (.A1(p_0[19]), .A2(accumulator[19]), .ZN(n_111));
   NOR4_X1 i_144 (.A1(n_116), .A2(n_113), .A3(n_117), .A4(n_120), .ZN(n_112));
   NOR2_X1 i_145 (.A1(n_125), .A2(n_115), .ZN(n_113));
   INV_X1 i_146 (.A(n_115), .ZN(n_114));
   NAND2_X1 i_147 (.A1(p_0[14]), .A2(accumulator[14]), .ZN(n_115));
   AND2_X1 i_148 (.A1(p_0[15]), .A2(accumulator[15]), .ZN(n_116));
   AOI21_X1 i_149 (.A(n_122), .B1(n_119), .B2(n_118), .ZN(n_117));
   NAND2_X1 i_150 (.A1(p_0[13]), .A2(accumulator[13]), .ZN(n_118));
   NAND2_X1 i_151 (.A1(p_0[12]), .A2(accumulator[12]), .ZN(n_119));
   NOR3_X1 i_152 (.A1(n_122), .A2(n_121), .A3(n_126), .ZN(n_120));
   NOR2_X1 i_153 (.A1(p_0[12]), .A2(accumulator[12]), .ZN(n_121));
   OR3_X1 i_154 (.A1(n_125), .A2(n_123), .A3(n_124), .ZN(n_122));
   NOR2_X1 i_155 (.A1(p_0[14]), .A2(accumulator[14]), .ZN(n_123));
   NOR2_X1 i_156 (.A1(p_0[13]), .A2(accumulator[13]), .ZN(n_124));
   NOR2_X1 i_157 (.A1(p_0[15]), .A2(accumulator[15]), .ZN(n_125));
   NOR4_X1 i_158 (.A1(n_130), .A2(n_127), .A3(n_131), .A4(n_134), .ZN(n_126));
   NOR2_X1 i_159 (.A1(n_139), .A2(n_129), .ZN(n_127));
   INV_X1 i_160 (.A(n_129), .ZN(n_128));
   NAND2_X1 i_161 (.A1(p_0[10]), .A2(accumulator[10]), .ZN(n_129));
   AND2_X1 i_162 (.A1(p_0[11]), .A2(accumulator[11]), .ZN(n_130));
   AOI21_X1 i_163 (.A(n_136), .B1(n_133), .B2(n_132), .ZN(n_131));
   NAND2_X1 i_164 (.A1(p_0[9]), .A2(accumulator[9]), .ZN(n_132));
   NAND2_X1 i_165 (.A1(p_0[8]), .A2(accumulator[8]), .ZN(n_133));
   NOR3_X1 i_166 (.A1(n_136), .A2(n_135), .A3(n_140), .ZN(n_134));
   NOR2_X1 i_167 (.A1(p_0[8]), .A2(accumulator[8]), .ZN(n_135));
   OR3_X1 i_168 (.A1(n_139), .A2(n_137), .A3(n_138), .ZN(n_136));
   NOR2_X1 i_169 (.A1(p_0[10]), .A2(accumulator[10]), .ZN(n_137));
   NOR2_X1 i_170 (.A1(p_0[9]), .A2(accumulator[9]), .ZN(n_138));
   NOR2_X1 i_171 (.A1(p_0[11]), .A2(accumulator[11]), .ZN(n_139));
   NOR4_X1 i_172 (.A1(n_144), .A2(n_141), .A3(n_145), .A4(n_148), .ZN(n_140));
   NOR2_X1 i_173 (.A1(n_153), .A2(n_143), .ZN(n_141));
   INV_X1 i_174 (.A(n_143), .ZN(n_142));
   NAND2_X1 i_175 (.A1(p_0[6]), .A2(accumulator[6]), .ZN(n_143));
   AND2_X1 i_176 (.A1(p_0[7]), .A2(accumulator[7]), .ZN(n_144));
   AOI21_X1 i_177 (.A(n_150), .B1(n_147), .B2(n_146), .ZN(n_145));
   NAND2_X1 i_178 (.A1(p_0[5]), .A2(accumulator[5]), .ZN(n_146));
   NAND2_X1 i_179 (.A1(p_0[4]), .A2(accumulator[4]), .ZN(n_147));
   NOR3_X1 i_180 (.A1(n_150), .A2(n_149), .A3(n_154), .ZN(n_148));
   NOR2_X1 i_181 (.A1(p_0[4]), .A2(accumulator[4]), .ZN(n_149));
   OR3_X1 i_182 (.A1(n_153), .A2(n_151), .A3(n_152), .ZN(n_150));
   NOR2_X1 i_183 (.A1(p_0[6]), .A2(accumulator[6]), .ZN(n_151));
   NOR2_X1 i_184 (.A1(p_0[5]), .A2(accumulator[5]), .ZN(n_152));
   NOR2_X1 i_185 (.A1(p_0[7]), .A2(accumulator[7]), .ZN(n_153));
   NAND2_X1 i_186 (.A1(n_163), .A2(n_155), .ZN(n_154));
   OAI21_X1 i_187 (.A(n_156), .B1(n_168), .B2(n_165), .ZN(n_155));
   OAI22_X1 i_188 (.A1(p_0[2]), .A2(accumulator[2]), .B1(n_161), .B2(n_157), 
      .ZN(n_156));
   AOI21_X1 i_189 (.A(n_160), .B1(n_159), .B2(n_158), .ZN(n_157));
   NAND2_X1 i_190 (.A1(p_0[1]), .A2(accumulator[1]), .ZN(n_158));
   NAND2_X1 i_191 (.A1(p_0[0]), .A2(accumulator[0]), .ZN(n_159));
   NOR2_X1 i_192 (.A1(p_0[1]), .A2(accumulator[1]), .ZN(n_160));
   INV_X1 i_193 (.A(n_162), .ZN(n_161));
   NAND2_X1 i_194 (.A1(p_0[2]), .A2(accumulator[2]), .ZN(n_162));
   NAND2_X1 i_195 (.A1(n_168), .A2(n_165), .ZN(n_163));
   NOR2_X1 i_196 (.A1(p_0[28]), .A2(accumulator[28]), .ZN(n_164));
   INV_X1 i_197 (.A(accumulator[3]), .ZN(n_165));
   INV_X1 i_198 (.A(accumulator[27]), .ZN(n_166));
   INV_X1 i_199 (.A(accumulator[29]), .ZN(n_167));
   INV_X1 i_200 (.A(p_0[3]), .ZN(n_168));
   INV_X1 i_201 (.A(p_0[27]), .ZN(n_169));
   INV_X1 i_202 (.A(p_0[29]), .ZN(n_170));
endmodule

module datapath__0_4(p_0, A);
   output [31:0]p_0;
   input [31:0]A;

   XOR2_X1 i_0 (.A(A[1]), .B(A[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(A[2]), .B1(A[1]), .B2(A[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(A[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(A[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(A[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(A[6]), .B1(n_27), .B2(A[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(A[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(A[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(A[9]), .B1(n_25), .B2(A[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(A[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(A[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(A[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(A[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(A[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(A[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(A[16]), .B1(n_19), .B2(A[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(A[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(A[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(A[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(A[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(A[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(A[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(A[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(A[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(A[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(A[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(A[27]), .B1(n_9), .B2(A[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(A[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(A[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(A[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(A[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(A[28]), .A3(A[29]), .A4(A[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(A[28]), .A3(A[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(A[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(A[26]), .A3(A[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(A[23]), .A3(A[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(A[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(A[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(A[18]), .A3(A[19]), .A4(A[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(A[18]), .A3(A[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(A[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(A[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(A[15]), .A3(A[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(A[12]), .A3(A[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(A[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(A[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(A[8]), .A3(A[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(A[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(A[5]), .A3(A[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(A[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(A[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(A[2]), .A2(A[1]), .A3(A[0]), .ZN(n_29));
   INV_X1 i_61 (.A(A[11]), .ZN(n_30));
   INV_X1 i_62 (.A(A[14]), .ZN(n_31));
   INV_X1 i_63 (.A(A[21]), .ZN(n_32));
   INV_X1 i_64 (.A(A[25]), .ZN(n_33));
endmodule

module datapath__0_6(p_0, B);
   output [31:0]p_0;
   input [31:0]B;

   XOR2_X1 i_0 (.A(B[1]), .B(B[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(B[2]), .B1(B[1]), .B2(B[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(B[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(B[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(B[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(B[6]), .B1(n_27), .B2(B[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(B[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(B[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(B[9]), .B1(n_25), .B2(B[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(B[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(B[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(B[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(B[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(B[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(B[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(B[16]), .B1(n_19), .B2(B[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(B[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(B[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(B[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(B[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(B[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(B[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(B[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(B[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(B[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(B[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(B[27]), .B1(n_9), .B2(B[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(B[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(B[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(B[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(B[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(B[28]), .A3(B[29]), .A4(B[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(B[28]), .A3(B[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(B[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(B[26]), .A3(B[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(B[23]), .A3(B[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(B[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(B[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(B[18]), .A3(B[19]), .A4(B[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(B[18]), .A3(B[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(B[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(B[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(B[15]), .A3(B[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(B[12]), .A3(B[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(B[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(B[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(B[8]), .A3(B[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(B[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(B[5]), .A3(B[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(B[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(B[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(B[2]), .A2(B[1]), .A3(B[0]), .ZN(n_29));
   INV_X1 i_61 (.A(B[11]), .ZN(n_30));
   INV_X1 i_62 (.A(B[14]), .ZN(n_31));
   INV_X1 i_63 (.A(B[21]), .ZN(n_32));
   INV_X1 i_64 (.A(B[25]), .ZN(n_33));
endmodule

module datapath__0_13(Res_imm, p_0);
   input [63:0]Res_imm;
   output [63:0]p_0;

   XOR2_X1 i_0 (.A(Res_imm[1]), .B(Res_imm[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_60), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(Res_imm[2]), .B1(Res_imm[1]), .B2(Res_imm[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(Res_imm[3]), .B(n_60), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(Res_imm[4]), .B(n_59), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(Res_imm[5]), .B(n_58), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_57), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(Res_imm[6]), .B1(n_58), .B2(Res_imm[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(Res_imm[7]), .B(n_57), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(Res_imm[8]), .B(n_56), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_55), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(Res_imm[9]), .B1(n_56), .B2(Res_imm[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(Res_imm[10]), .B(n_55), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(Res_imm[11]), .B(n_54), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(Res_imm[12]), .B(n_53), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(Res_imm[13]), .B(n_52), .ZN(p_0[13]));
   XOR2_X1 i_16 (.A(Res_imm[14]), .B(n_51), .Z(p_0[14]));
   AND2_X1 i_17 (.A1(n_50), .A2(n_3), .ZN(p_0[15]));
   OAI21_X1 i_18 (.A(Res_imm[15]), .B1(n_51), .B2(Res_imm[14]), .ZN(n_3));
   XOR2_X1 i_19 (.A(Res_imm[16]), .B(n_50), .Z(p_0[16]));
   XOR2_X1 i_20 (.A(Res_imm[17]), .B(n_49), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(Res_imm[18]), .B(n_48), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(Res_imm[19]), .B(n_47), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(Res_imm[20]), .B(n_46), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(Res_imm[21]), .B(n_45), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(Res_imm[22]), .B(n_44), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(Res_imm[23]), .B(n_43), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(Res_imm[24]), .B(n_42), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(Res_imm[25]), .B(n_41), .ZN(p_0[25]));
   XNOR2_X1 i_29 (.A(Res_imm[26]), .B(n_40), .ZN(p_0[26]));
   XOR2_X1 i_30 (.A(Res_imm[27]), .B(n_39), .Z(p_0[27]));
   XOR2_X1 i_31 (.A(Res_imm[28]), .B(n_38), .Z(p_0[28]));
   XNOR2_X1 i_32 (.A(Res_imm[29]), .B(n_37), .ZN(p_0[29]));
   XNOR2_X1 i_33 (.A(Res_imm[30]), .B(n_36), .ZN(p_0[30]));
   XNOR2_X1 i_34 (.A(Res_imm[31]), .B(n_35), .ZN(p_0[31]));
   XOR2_X1 i_35 (.A(Res_imm[32]), .B(n_34), .Z(p_0[32]));
   XOR2_X1 i_36 (.A(Res_imm[33]), .B(n_33), .Z(p_0[33]));
   XNOR2_X1 i_37 (.A(Res_imm[34]), .B(n_32), .ZN(p_0[34]));
   XNOR2_X1 i_38 (.A(Res_imm[35]), .B(n_31), .ZN(p_0[35]));
   XNOR2_X1 i_39 (.A(Res_imm[36]), .B(n_30), .ZN(p_0[36]));
   XOR2_X1 i_40 (.A(Res_imm[37]), .B(n_29), .Z(p_0[37]));
   XOR2_X1 i_41 (.A(Res_imm[38]), .B(n_28), .Z(p_0[38]));
   XNOR2_X1 i_42 (.A(Res_imm[39]), .B(n_27), .ZN(p_0[39]));
   XNOR2_X1 i_43 (.A(Res_imm[40]), .B(n_26), .ZN(p_0[40]));
   XOR2_X1 i_44 (.A(Res_imm[41]), .B(n_25), .Z(p_0[41]));
   XNOR2_X1 i_45 (.A(Res_imm[42]), .B(n_24), .ZN(p_0[42]));
   XOR2_X1 i_46 (.A(Res_imm[43]), .B(n_23), .Z(p_0[43]));
   AND2_X1 i_47 (.A1(n_22), .A2(n_4), .ZN(p_0[44]));
   OAI21_X1 i_48 (.A(Res_imm[44]), .B1(n_23), .B2(Res_imm[43]), .ZN(n_4));
   XOR2_X1 i_49 (.A(Res_imm[45]), .B(n_22), .Z(p_0[45]));
   XOR2_X1 i_50 (.A(Res_imm[46]), .B(n_21), .Z(p_0[46]));
   XOR2_X1 i_51 (.A(Res_imm[47]), .B(n_20), .Z(p_0[47]));
   XOR2_X1 i_52 (.A(Res_imm[48]), .B(n_19), .Z(p_0[48]));
   XNOR2_X1 i_53 (.A(Res_imm[49]), .B(n_18), .ZN(p_0[49]));
   XNOR2_X1 i_54 (.A(Res_imm[50]), .B(n_17), .ZN(p_0[50]));
   XNOR2_X1 i_55 (.A(Res_imm[51]), .B(n_16), .ZN(p_0[51]));
   XOR2_X1 i_56 (.A(Res_imm[52]), .B(n_15), .Z(p_0[52]));
   XNOR2_X1 i_57 (.A(Res_imm[53]), .B(n_14), .ZN(p_0[53]));
   XNOR2_X1 i_58 (.A(Res_imm[54]), .B(n_13), .ZN(p_0[54]));
   XNOR2_X1 i_59 (.A(Res_imm[55]), .B(n_12), .ZN(p_0[55]));
   XOR2_X1 i_60 (.A(Res_imm[56]), .B(n_11), .Z(p_0[56]));
   AND2_X1 i_61 (.A1(n_10), .A2(n_5), .ZN(p_0[57]));
   OAI21_X1 i_62 (.A(Res_imm[57]), .B1(n_11), .B2(Res_imm[56]), .ZN(n_5));
   XOR2_X1 i_63 (.A(Res_imm[58]), .B(n_10), .Z(p_0[58]));
   XNOR2_X1 i_64 (.A(Res_imm[59]), .B(n_9), .ZN(p_0[59]));
   XNOR2_X1 i_65 (.A(Res_imm[60]), .B(n_8), .ZN(p_0[60]));
   XOR2_X1 i_66 (.A(Res_imm[61]), .B(n_7), .Z(p_0[61]));
   XNOR2_X1 i_67 (.A(Res_imm[62]), .B(n_6), .ZN(p_0[62]));
   NAND2_X1 i_68 (.A1(n_6), .A2(n_72), .ZN(p_0[63]));
   NOR2_X1 i_69 (.A1(n_7), .A2(Res_imm[61]), .ZN(n_6));
   NAND2_X1 i_70 (.A1(n_8), .A2(n_71), .ZN(n_7));
   NOR3_X1 i_71 (.A1(n_10), .A2(Res_imm[58]), .A3(Res_imm[59]), .ZN(n_8));
   NOR2_X1 i_72 (.A1(n_10), .A2(Res_imm[58]), .ZN(n_9));
   OR3_X1 i_73 (.A1(n_11), .A2(Res_imm[56]), .A3(Res_imm[57]), .ZN(n_10));
   NAND2_X1 i_74 (.A1(n_12), .A2(n_70), .ZN(n_11));
   NOR4_X1 i_75 (.A1(n_15), .A2(Res_imm[52]), .A3(Res_imm[53]), .A4(Res_imm[54]), 
      .ZN(n_12));
   NOR3_X1 i_76 (.A1(n_15), .A2(Res_imm[52]), .A3(Res_imm[53]), .ZN(n_13));
   NOR2_X1 i_77 (.A1(n_15), .A2(Res_imm[52]), .ZN(n_14));
   NAND2_X1 i_78 (.A1(n_16), .A2(n_69), .ZN(n_15));
   NOR4_X1 i_79 (.A1(n_19), .A2(Res_imm[48]), .A3(Res_imm[49]), .A4(Res_imm[50]), 
      .ZN(n_16));
   NOR3_X1 i_80 (.A1(n_19), .A2(Res_imm[48]), .A3(Res_imm[49]), .ZN(n_17));
   NOR2_X1 i_81 (.A1(n_19), .A2(Res_imm[48]), .ZN(n_18));
   OR2_X1 i_82 (.A1(n_20), .A2(Res_imm[47]), .ZN(n_19));
   OR2_X1 i_83 (.A1(n_21), .A2(Res_imm[46]), .ZN(n_20));
   OR2_X1 i_84 (.A1(n_22), .A2(Res_imm[45]), .ZN(n_21));
   OR3_X1 i_85 (.A1(n_23), .A2(Res_imm[43]), .A3(Res_imm[44]), .ZN(n_22));
   NAND2_X1 i_86 (.A1(n_24), .A2(n_68), .ZN(n_23));
   NOR2_X1 i_87 (.A1(n_25), .A2(Res_imm[41]), .ZN(n_24));
   NAND2_X1 i_88 (.A1(n_26), .A2(n_67), .ZN(n_25));
   NOR3_X1 i_89 (.A1(n_28), .A2(Res_imm[38]), .A3(Res_imm[39]), .ZN(n_26));
   NOR2_X1 i_90 (.A1(n_28), .A2(Res_imm[38]), .ZN(n_27));
   OR2_X1 i_91 (.A1(n_29), .A2(Res_imm[37]), .ZN(n_28));
   NAND2_X1 i_92 (.A1(n_30), .A2(n_66), .ZN(n_29));
   NOR4_X1 i_93 (.A1(n_33), .A2(Res_imm[33]), .A3(Res_imm[34]), .A4(Res_imm[35]), 
      .ZN(n_30));
   NOR3_X1 i_94 (.A1(n_33), .A2(Res_imm[33]), .A3(Res_imm[34]), .ZN(n_31));
   NOR2_X1 i_95 (.A1(n_33), .A2(Res_imm[33]), .ZN(n_32));
   OR2_X1 i_96 (.A1(n_34), .A2(Res_imm[32]), .ZN(n_33));
   NAND2_X1 i_97 (.A1(n_35), .A2(n_65), .ZN(n_34));
   NOR4_X1 i_98 (.A1(n_38), .A2(Res_imm[28]), .A3(Res_imm[29]), .A4(Res_imm[30]), 
      .ZN(n_35));
   NOR3_X1 i_99 (.A1(n_38), .A2(Res_imm[28]), .A3(Res_imm[29]), .ZN(n_36));
   NOR2_X1 i_100 (.A1(n_38), .A2(Res_imm[28]), .ZN(n_37));
   OR2_X1 i_101 (.A1(n_39), .A2(Res_imm[27]), .ZN(n_38));
   NAND2_X1 i_102 (.A1(n_40), .A2(n_64), .ZN(n_39));
   NOR4_X1 i_103 (.A1(n_43), .A2(Res_imm[23]), .A3(Res_imm[24]), .A4(Res_imm[25]), 
      .ZN(n_40));
   NOR3_X1 i_104 (.A1(n_43), .A2(Res_imm[23]), .A3(Res_imm[24]), .ZN(n_41));
   NOR2_X1 i_105 (.A1(n_43), .A2(Res_imm[23]), .ZN(n_42));
   OR2_X1 i_106 (.A1(n_44), .A2(Res_imm[22]), .ZN(n_43));
   NAND2_X1 i_107 (.A1(n_45), .A2(n_63), .ZN(n_44));
   NOR4_X1 i_108 (.A1(n_48), .A2(Res_imm[18]), .A3(Res_imm[19]), .A4(Res_imm[20]), 
      .ZN(n_45));
   NOR3_X1 i_109 (.A1(n_48), .A2(Res_imm[18]), .A3(Res_imm[19]), .ZN(n_46));
   NOR2_X1 i_110 (.A1(n_48), .A2(Res_imm[18]), .ZN(n_47));
   OR2_X1 i_111 (.A1(n_49), .A2(Res_imm[17]), .ZN(n_48));
   OR2_X1 i_112 (.A1(n_50), .A2(Res_imm[16]), .ZN(n_49));
   OR3_X1 i_113 (.A1(n_51), .A2(Res_imm[14]), .A3(Res_imm[15]), .ZN(n_50));
   NAND2_X1 i_114 (.A1(n_52), .A2(n_62), .ZN(n_51));
   NOR2_X1 i_115 (.A1(n_53), .A2(Res_imm[12]), .ZN(n_52));
   NAND2_X1 i_116 (.A1(n_54), .A2(n_61), .ZN(n_53));
   NOR2_X1 i_117 (.A1(n_55), .A2(Res_imm[10]), .ZN(n_54));
   OR3_X1 i_118 (.A1(n_56), .A2(Res_imm[8]), .A3(Res_imm[9]), .ZN(n_55));
   OR2_X1 i_119 (.A1(n_57), .A2(Res_imm[7]), .ZN(n_56));
   OR3_X1 i_120 (.A1(n_58), .A2(Res_imm[5]), .A3(Res_imm[6]), .ZN(n_57));
   OR2_X1 i_121 (.A1(n_59), .A2(Res_imm[4]), .ZN(n_58));
   OR2_X1 i_122 (.A1(n_60), .A2(Res_imm[3]), .ZN(n_59));
   OR3_X1 i_123 (.A1(Res_imm[2]), .A2(Res_imm[1]), .A3(Res_imm[0]), .ZN(n_60));
   INV_X1 i_124 (.A(Res_imm[11]), .ZN(n_61));
   INV_X1 i_125 (.A(Res_imm[13]), .ZN(n_62));
   INV_X1 i_126 (.A(Res_imm[21]), .ZN(n_63));
   INV_X1 i_127 (.A(Res_imm[26]), .ZN(n_64));
   INV_X1 i_128 (.A(Res_imm[31]), .ZN(n_65));
   INV_X1 i_129 (.A(Res_imm[36]), .ZN(n_66));
   INV_X1 i_130 (.A(Res_imm[40]), .ZN(n_67));
   INV_X1 i_131 (.A(Res_imm[42]), .ZN(n_68));
   INV_X1 i_132 (.A(Res_imm[51]), .ZN(n_69));
   INV_X1 i_133 (.A(Res_imm[55]), .ZN(n_70));
   INV_X1 i_134 (.A(Res_imm[60]), .ZN(n_71));
   INV_X1 i_135 (.A(Res_imm[62]), .ZN(n_72));
endmodule

module sequentialMultiplier(Res, OVF, A, B, clk, reset, enable);
   output [63:0]Res;
   output OVF;
   input [31:0]A;
   input [31:0]B;
   input clk;
   input reset;
   input enable;

   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire [1:0]isNeg;
   wire [31:0]accumulator;
   wire [31:0]multiplier;
   wire [31:0]multiplicand;
   wire ready;
   wire n_0_159;
   wire [4:0]counter;
   wire n_0_0;
   wire n_0_1;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire [4:0]counter_in;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_160;
   wire n_0_161;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire [31:0]multiplicand_in;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_162;
   wire n_0_163;
   wire n_0_0_65;
   wire n_0_164;
   wire n_0_0_66;
   wire n_0_165;
   wire n_0_0_67;
   wire n_0_166;
   wire n_0_0_68;
   wire n_0_167;
   wire n_0_0_69;
   wire n_0_168;
   wire n_0_0_70;
   wire n_0_169;
   wire n_0_0_71;
   wire n_0_170;
   wire n_0_0_72;
   wire n_0_171;
   wire n_0_0_73;
   wire n_0_172;
   wire n_0_0_74;
   wire n_0_173;
   wire n_0_0_75;
   wire n_0_174;
   wire n_0_0_76;
   wire n_0_175;
   wire n_0_0_77;
   wire n_0_176;
   wire n_0_0_78;
   wire n_0_177;
   wire n_0_0_79;
   wire n_0_178;
   wire n_0_0_80;
   wire n_0_179;
   wire n_0_0_81;
   wire n_0_180;
   wire n_0_0_82;
   wire n_0_181;
   wire n_0_0_83;
   wire n_0_182;
   wire n_0_0_84;
   wire n_0_183;
   wire n_0_0_85;
   wire n_0_184;
   wire n_0_0_86;
   wire n_0_185;
   wire n_0_0_87;
   wire n_0_186;
   wire n_0_0_88;
   wire n_0_187;
   wire n_0_0_89;
   wire n_0_188;
   wire n_0_0_90;
   wire n_0_189;
   wire n_0_0_91;
   wire n_0_190;
   wire n_0_0_92;
   wire n_0_191;
   wire n_0_0_93;
   wire n_0_192;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_193;
   wire n_0_0_98;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire [1:0]isNeg_in;
   wire n_0_258;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_31;
   wire n_0_0_97;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_108;

   datapath i_0_5 (.p_0({n_0_256, n_0_255, n_0_254, n_0_253, n_0_252, n_0_251, 
      n_0_250, n_0_249, n_0_248, n_0_247, n_0_246, n_0_245, n_0_244, n_0_243, 
      n_0_242, n_0_241, n_0_240, n_0_239, n_0_238, n_0_237, n_0_236, n_0_235, 
      n_0_234, n_0_233, n_0_232, n_0_231, n_0_230, n_0_229, n_0_228, n_0_227, 
      n_0_226, n_0_225}), .accumulator({uc_0, accumulator[30], accumulator[29], 
      accumulator[28], accumulator[27], accumulator[26], accumulator[25], 
      accumulator[24], accumulator[23], accumulator[22], accumulator[21], 
      accumulator[20], accumulator[19], accumulator[18], accumulator[17], 
      accumulator[16], accumulator[15], accumulator[14], accumulator[13], 
      accumulator[12], accumulator[11], accumulator[10], accumulator[9], 
      accumulator[8], accumulator[7], accumulator[6], accumulator[5], 
      accumulator[4], accumulator[3], accumulator[2], accumulator[1], 
      accumulator[0]}), .p_1({n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, 
      n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, 
      n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, 
      n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2}));
   datapath__0_4 i_0_7 (.p_0({n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, 
      n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, 
      n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, 
      n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, uc_1}), .A(A));
   datapath__0_6 i_0_9 (.p_0({n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, 
      n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, 
      n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, 
      n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, uc_2}), .B(B));
   datapath__0_13 i_0_16 (.Res_imm({uc_3, accumulator[30], accumulator[29], 
      accumulator[28], accumulator[27], accumulator[26], accumulator[25], 
      accumulator[24], accumulator[23], accumulator[22], accumulator[21], 
      accumulator[20], accumulator[19], accumulator[18], accumulator[17], 
      accumulator[16], accumulator[15], accumulator[14], accumulator[13], 
      accumulator[12], accumulator[11], accumulator[10], accumulator[9], 
      accumulator[8], accumulator[7], accumulator[6], accumulator[5], 
      accumulator[4], accumulator[3], accumulator[2], accumulator[1], 
      accumulator[0], multiplicand[31], multiplicand[30], multiplicand[29], 
      multiplicand[28], multiplicand[27], multiplicand[26], multiplicand[25], 
      multiplicand[24], multiplicand[23], multiplicand[22], multiplicand[21], 
      multiplicand[20], multiplicand[19], multiplicand[18], multiplicand[17], 
      multiplicand[16], multiplicand[15], multiplicand[14], multiplicand[13], 
      multiplicand[12], multiplicand[11], multiplicand[10], multiplicand[9], 
      multiplicand[8], multiplicand[7], multiplicand[6], multiplicand[5], 
      multiplicand[4], multiplicand[3], multiplicand[2], multiplicand[1], Res[0]}), 
      .p_0({n_0_158, n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, 
      n_0_151, n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, 
      n_0_143, n_0_142, n_0_141, n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, 
      n_0_135, n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, 
      n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, 
      n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, 
      n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, 
      n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, uc_4}));
   DFF_X1 \isNeg_reg[1]  (.D(isNeg_in[1]), .CK(n_0_1), .Q(isNeg[1]), .QN());
   DFF_X1 \isNeg_reg[0]  (.D(isNeg_in[0]), .CK(n_0_1), .Q(isNeg[0]), .QN());
   DFF_X1 \accumulator_reg[30]  (.D(n_0_224), .CK(n_0_0), .Q(accumulator[30]), 
      .QN());
   DFF_X1 \accumulator_reg[29]  (.D(n_0_223), .CK(n_0_0), .Q(accumulator[29]), 
      .QN());
   DFF_X1 \accumulator_reg[28]  (.D(n_0_222), .CK(n_0_0), .Q(accumulator[28]), 
      .QN());
   DFF_X1 \accumulator_reg[27]  (.D(n_0_221), .CK(n_0_0), .Q(accumulator[27]), 
      .QN());
   DFF_X1 \accumulator_reg[26]  (.D(n_0_220), .CK(n_0_0), .Q(accumulator[26]), 
      .QN());
   DFF_X1 \accumulator_reg[25]  (.D(n_0_219), .CK(n_0_0), .Q(accumulator[25]), 
      .QN());
   DFF_X1 \accumulator_reg[24]  (.D(n_0_218), .CK(n_0_0), .Q(accumulator[24]), 
      .QN());
   DFF_X1 \accumulator_reg[23]  (.D(n_0_217), .CK(n_0_0), .Q(accumulator[23]), 
      .QN());
   DFF_X1 \accumulator_reg[22]  (.D(n_0_216), .CK(n_0_0), .Q(accumulator[22]), 
      .QN());
   DFF_X1 \accumulator_reg[21]  (.D(n_0_215), .CK(n_0_0), .Q(accumulator[21]), 
      .QN());
   DFF_X1 \accumulator_reg[20]  (.D(n_0_214), .CK(n_0_0), .Q(accumulator[20]), 
      .QN());
   DFF_X1 \accumulator_reg[19]  (.D(n_0_213), .CK(n_0_0), .Q(accumulator[19]), 
      .QN());
   DFF_X1 \accumulator_reg[18]  (.D(n_0_212), .CK(n_0_0), .Q(accumulator[18]), 
      .QN());
   DFF_X1 \accumulator_reg[17]  (.D(n_0_211), .CK(n_0_0), .Q(accumulator[17]), 
      .QN());
   DFF_X1 \accumulator_reg[16]  (.D(n_0_210), .CK(n_0_0), .Q(accumulator[16]), 
      .QN());
   DFF_X1 \accumulator_reg[15]  (.D(n_0_209), .CK(n_0_0), .Q(accumulator[15]), 
      .QN());
   DFF_X1 \accumulator_reg[14]  (.D(n_0_208), .CK(n_0_0), .Q(accumulator[14]), 
      .QN());
   DFF_X1 \accumulator_reg[13]  (.D(n_0_207), .CK(n_0_0), .Q(accumulator[13]), 
      .QN());
   DFF_X1 \accumulator_reg[12]  (.D(n_0_206), .CK(n_0_0), .Q(accumulator[12]), 
      .QN());
   DFF_X1 \accumulator_reg[11]  (.D(n_0_205), .CK(n_0_0), .Q(accumulator[11]), 
      .QN());
   DFF_X1 \accumulator_reg[10]  (.D(n_0_204), .CK(n_0_0), .Q(accumulator[10]), 
      .QN());
   DFF_X1 \accumulator_reg[9]  (.D(n_0_203), .CK(n_0_0), .Q(accumulator[9]), 
      .QN());
   DFF_X1 \accumulator_reg[8]  (.D(n_0_202), .CK(n_0_0), .Q(accumulator[8]), 
      .QN());
   DFF_X1 \accumulator_reg[7]  (.D(n_0_201), .CK(n_0_0), .Q(accumulator[7]), 
      .QN());
   DFF_X1 \accumulator_reg[6]  (.D(n_0_200), .CK(n_0_0), .Q(accumulator[6]), 
      .QN());
   DFF_X1 \accumulator_reg[5]  (.D(n_0_199), .CK(n_0_0), .Q(accumulator[5]), 
      .QN());
   DFF_X1 \accumulator_reg[4]  (.D(n_0_198), .CK(n_0_0), .Q(accumulator[4]), 
      .QN());
   DFF_X1 \accumulator_reg[3]  (.D(n_0_197), .CK(n_0_0), .Q(accumulator[3]), 
      .QN());
   DFF_X1 \accumulator_reg[2]  (.D(n_0_196), .CK(n_0_0), .Q(accumulator[2]), 
      .QN());
   DFF_X1 \accumulator_reg[1]  (.D(n_0_195), .CK(n_0_0), .Q(accumulator[1]), 
      .QN());
   DFF_X1 \accumulator_reg[0]  (.D(n_0_194), .CK(n_0_0), .Q(accumulator[0]), 
      .QN());
   DFF_X1 \multiplier_reg[31]  (.D(n_0_193), .CK(n_0_1), .Q(multiplier[31]), 
      .QN());
   DFF_X1 \multiplier_reg[30]  (.D(n_0_192), .CK(n_0_1), .Q(multiplier[30]), 
      .QN());
   DFF_X1 \multiplier_reg[29]  (.D(n_0_191), .CK(n_0_1), .Q(multiplier[29]), 
      .QN());
   DFF_X1 \multiplier_reg[28]  (.D(n_0_190), .CK(n_0_1), .Q(multiplier[28]), 
      .QN());
   DFF_X1 \multiplier_reg[27]  (.D(n_0_189), .CK(n_0_1), .Q(multiplier[27]), 
      .QN());
   DFF_X1 \multiplier_reg[26]  (.D(n_0_188), .CK(n_0_1), .Q(multiplier[26]), 
      .QN());
   DFF_X1 \multiplier_reg[25]  (.D(n_0_187), .CK(n_0_1), .Q(multiplier[25]), 
      .QN());
   DFF_X1 \multiplier_reg[24]  (.D(n_0_186), .CK(n_0_1), .Q(multiplier[24]), 
      .QN());
   DFF_X1 \multiplier_reg[23]  (.D(n_0_185), .CK(n_0_1), .Q(multiplier[23]), 
      .QN());
   DFF_X1 \multiplier_reg[22]  (.D(n_0_184), .CK(n_0_1), .Q(multiplier[22]), 
      .QN());
   DFF_X1 \multiplier_reg[21]  (.D(n_0_183), .CK(n_0_1), .Q(multiplier[21]), 
      .QN());
   DFF_X1 \multiplier_reg[20]  (.D(n_0_182), .CK(n_0_1), .Q(multiplier[20]), 
      .QN());
   DFF_X1 \multiplier_reg[19]  (.D(n_0_181), .CK(n_0_1), .Q(multiplier[19]), 
      .QN());
   DFF_X1 \multiplier_reg[18]  (.D(n_0_180), .CK(n_0_1), .Q(multiplier[18]), 
      .QN());
   DFF_X1 \multiplier_reg[17]  (.D(n_0_179), .CK(n_0_1), .Q(multiplier[17]), 
      .QN());
   DFF_X1 \multiplier_reg[16]  (.D(n_0_178), .CK(n_0_1), .Q(multiplier[16]), 
      .QN());
   DFF_X1 \multiplier_reg[15]  (.D(n_0_177), .CK(n_0_1), .Q(multiplier[15]), 
      .QN());
   DFF_X1 \multiplier_reg[14]  (.D(n_0_176), .CK(n_0_1), .Q(multiplier[14]), 
      .QN());
   DFF_X1 \multiplier_reg[13]  (.D(n_0_175), .CK(n_0_1), .Q(multiplier[13]), 
      .QN());
   DFF_X1 \multiplier_reg[12]  (.D(n_0_174), .CK(n_0_1), .Q(multiplier[12]), 
      .QN());
   DFF_X1 \multiplier_reg[11]  (.D(n_0_173), .CK(n_0_1), .Q(multiplier[11]), 
      .QN());
   DFF_X1 \multiplier_reg[10]  (.D(n_0_172), .CK(n_0_1), .Q(multiplier[10]), 
      .QN());
   DFF_X1 \multiplier_reg[9]  (.D(n_0_171), .CK(n_0_1), .Q(multiplier[9]), .QN());
   DFF_X1 \multiplier_reg[8]  (.D(n_0_170), .CK(n_0_1), .Q(multiplier[8]), .QN());
   DFF_X1 \multiplier_reg[7]  (.D(n_0_169), .CK(n_0_1), .Q(multiplier[7]), .QN());
   DFF_X1 \multiplier_reg[6]  (.D(n_0_168), .CK(n_0_1), .Q(multiplier[6]), .QN());
   DFF_X1 \multiplier_reg[5]  (.D(n_0_167), .CK(n_0_1), .Q(multiplier[5]), .QN());
   DFF_X1 \multiplier_reg[4]  (.D(n_0_166), .CK(n_0_1), .Q(multiplier[4]), .QN());
   DFF_X1 \multiplier_reg[3]  (.D(n_0_165), .CK(n_0_1), .Q(multiplier[3]), .QN());
   DFF_X1 \multiplier_reg[2]  (.D(n_0_164), .CK(n_0_1), .Q(multiplier[2]), .QN());
   DFF_X1 \multiplier_reg[1]  (.D(n_0_163), .CK(n_0_1), .Q(multiplier[1]), .QN());
   DFF_X1 \multiplier_reg[0]  (.D(n_0_162), .CK(n_0_1), .Q(multiplier[0]), .QN());
   DFF_X1 \multiplicand_reg[31]  (.D(multiplicand_in[31]), .CK(n_0_0), .Q(
      multiplicand[31]), .QN());
   DFF_X1 \multiplicand_reg[30]  (.D(multiplicand_in[30]), .CK(n_0_0), .Q(
      multiplicand[30]), .QN());
   DFF_X1 \multiplicand_reg[29]  (.D(multiplicand_in[29]), .CK(n_0_0), .Q(
      multiplicand[29]), .QN());
   DFF_X1 \multiplicand_reg[28]  (.D(multiplicand_in[28]), .CK(n_0_0), .Q(
      multiplicand[28]), .QN());
   DFF_X1 \multiplicand_reg[27]  (.D(multiplicand_in[27]), .CK(n_0_0), .Q(
      multiplicand[27]), .QN());
   DFF_X1 \multiplicand_reg[26]  (.D(multiplicand_in[26]), .CK(n_0_0), .Q(
      multiplicand[26]), .QN());
   DFF_X1 \multiplicand_reg[25]  (.D(multiplicand_in[25]), .CK(n_0_0), .Q(
      multiplicand[25]), .QN());
   DFF_X1 \multiplicand_reg[24]  (.D(multiplicand_in[24]), .CK(n_0_0), .Q(
      multiplicand[24]), .QN());
   DFF_X1 \multiplicand_reg[23]  (.D(multiplicand_in[23]), .CK(n_0_0), .Q(
      multiplicand[23]), .QN());
   DFF_X1 \multiplicand_reg[22]  (.D(multiplicand_in[22]), .CK(n_0_0), .Q(
      multiplicand[22]), .QN());
   DFF_X1 \multiplicand_reg[21]  (.D(multiplicand_in[21]), .CK(n_0_0), .Q(
      multiplicand[21]), .QN());
   DFF_X1 \multiplicand_reg[20]  (.D(multiplicand_in[20]), .CK(n_0_0), .Q(
      multiplicand[20]), .QN());
   DFF_X1 \multiplicand_reg[19]  (.D(multiplicand_in[19]), .CK(n_0_0), .Q(
      multiplicand[19]), .QN());
   DFF_X1 \multiplicand_reg[18]  (.D(multiplicand_in[18]), .CK(n_0_0), .Q(
      multiplicand[18]), .QN());
   DFF_X1 \multiplicand_reg[17]  (.D(multiplicand_in[17]), .CK(n_0_0), .Q(
      multiplicand[17]), .QN());
   DFF_X1 \multiplicand_reg[16]  (.D(multiplicand_in[16]), .CK(n_0_0), .Q(
      multiplicand[16]), .QN());
   DFF_X1 \multiplicand_reg[15]  (.D(multiplicand_in[15]), .CK(n_0_0), .Q(
      multiplicand[15]), .QN());
   DFF_X1 \multiplicand_reg[14]  (.D(multiplicand_in[14]), .CK(n_0_0), .Q(
      multiplicand[14]), .QN());
   DFF_X1 \multiplicand_reg[13]  (.D(multiplicand_in[13]), .CK(n_0_0), .Q(
      multiplicand[13]), .QN());
   DFF_X1 \multiplicand_reg[12]  (.D(multiplicand_in[12]), .CK(n_0_0), .Q(
      multiplicand[12]), .QN());
   DFF_X1 \multiplicand_reg[11]  (.D(multiplicand_in[11]), .CK(n_0_0), .Q(
      multiplicand[11]), .QN());
   DFF_X1 \multiplicand_reg[10]  (.D(multiplicand_in[10]), .CK(n_0_0), .Q(
      multiplicand[10]), .QN());
   DFF_X1 \multiplicand_reg[9]  (.D(multiplicand_in[9]), .CK(n_0_0), .Q(
      multiplicand[9]), .QN());
   DFF_X1 \multiplicand_reg[8]  (.D(multiplicand_in[8]), .CK(n_0_0), .Q(
      multiplicand[8]), .QN());
   DFF_X1 \multiplicand_reg[7]  (.D(multiplicand_in[7]), .CK(n_0_0), .Q(
      multiplicand[7]), .QN());
   DFF_X1 \multiplicand_reg[6]  (.D(multiplicand_in[6]), .CK(n_0_0), .Q(
      multiplicand[6]), .QN());
   DFF_X1 \multiplicand_reg[5]  (.D(multiplicand_in[5]), .CK(n_0_0), .Q(
      multiplicand[5]), .QN());
   DFF_X1 \multiplicand_reg[4]  (.D(multiplicand_in[4]), .CK(n_0_0), .Q(
      multiplicand[4]), .QN());
   DFF_X1 \multiplicand_reg[3]  (.D(multiplicand_in[3]), .CK(n_0_0), .Q(
      multiplicand[3]), .QN());
   DFF_X1 \multiplicand_reg[2]  (.D(multiplicand_in[2]), .CK(n_0_0), .Q(
      multiplicand[2]), .QN());
   DFF_X1 \multiplicand_reg[1]  (.D(multiplicand_in[1]), .CK(n_0_0), .Q(
      multiplicand[1]), .QN());
   DFF_X1 \multiplicand_reg[0]  (.D(multiplicand_in[0]), .CK(n_0_0), .Q(Res[0]), 
      .QN());
   DFF_X1 ready_reg (.D(n_0_159), .CK(clk), .Q(ready), .QN());
   MUX2_X1 ready_reg_enable_mux_0 (.A(ready), .B(n_0_160), .S(n_0_161), .Z(
      n_0_159));
   DFF_X1 \counter_reg[4]  (.D(counter_in[4]), .CK(n_0_0), .Q(counter[4]), .QN());
   DFF_X1 \counter_reg[3]  (.D(counter_in[3]), .CK(n_0_0), .Q(counter[3]), .QN());
   DFF_X1 \counter_reg[2]  (.D(counter_in[2]), .CK(n_0_0), .Q(counter[2]), .QN());
   DFF_X1 \counter_reg[1]  (.D(counter_in[1]), .CK(n_0_0), .Q(counter[1]), .QN());
   DFF_X1 \counter_reg[0]  (.D(counter_in[0]), .CK(n_0_0), .Q(counter[0]), .QN());
   CLKGATETST_X1 clk_gate_accumulator_reg (.CK(clk), .E(n_0_257), .SE(1'b0), 
      .GCK(n_0_0));
   CLKGATETST_X1 clk_gate_isNeg_reg (.CK(clk), .E(n_0_258), .SE(1'b0), .GCK(
      n_0_1));
   NOR2_X1 i_0_0_0 (.A1(Res[63]), .A2(n_0_0_101), .ZN(OVF));
   MUX2_X1 i_0_0_1 (.A(n_0_96), .B(multiplicand[1]), .S(n_0_0_0), .Z(Res[1]));
   MUX2_X1 i_0_0_2 (.A(n_0_97), .B(multiplicand[2]), .S(n_0_0_0), .Z(Res[2]));
   MUX2_X1 i_0_0_3 (.A(n_0_98), .B(multiplicand[3]), .S(n_0_0_0), .Z(Res[3]));
   MUX2_X1 i_0_0_4 (.A(n_0_99), .B(multiplicand[4]), .S(n_0_0_0), .Z(Res[4]));
   MUX2_X1 i_0_0_5 (.A(n_0_100), .B(multiplicand[5]), .S(n_0_0_0), .Z(Res[5]));
   MUX2_X1 i_0_0_6 (.A(n_0_101), .B(multiplicand[6]), .S(n_0_0_0), .Z(Res[6]));
   MUX2_X1 i_0_0_7 (.A(n_0_102), .B(multiplicand[7]), .S(n_0_0_0), .Z(Res[7]));
   MUX2_X1 i_0_0_8 (.A(n_0_103), .B(multiplicand[8]), .S(n_0_0_0), .Z(Res[8]));
   MUX2_X1 i_0_0_9 (.A(n_0_104), .B(multiplicand[9]), .S(n_0_0_0), .Z(Res[9]));
   MUX2_X1 i_0_0_10 (.A(n_0_105), .B(multiplicand[10]), .S(n_0_0_0), .Z(Res[10]));
   MUX2_X1 i_0_0_11 (.A(n_0_106), .B(multiplicand[11]), .S(n_0_0_0), .Z(Res[11]));
   MUX2_X1 i_0_0_12 (.A(n_0_107), .B(multiplicand[12]), .S(n_0_0_0), .Z(Res[12]));
   MUX2_X1 i_0_0_13 (.A(n_0_108), .B(multiplicand[13]), .S(n_0_0_0), .Z(Res[13]));
   MUX2_X1 i_0_0_14 (.A(n_0_109), .B(multiplicand[14]), .S(n_0_0_0), .Z(Res[14]));
   MUX2_X1 i_0_0_15 (.A(n_0_110), .B(multiplicand[15]), .S(n_0_0_0), .Z(Res[15]));
   MUX2_X1 i_0_0_16 (.A(n_0_111), .B(multiplicand[16]), .S(n_0_0_0), .Z(Res[16]));
   MUX2_X1 i_0_0_17 (.A(n_0_112), .B(multiplicand[17]), .S(n_0_0_0), .Z(Res[17]));
   MUX2_X1 i_0_0_18 (.A(n_0_113), .B(multiplicand[18]), .S(n_0_0_0), .Z(Res[18]));
   MUX2_X1 i_0_0_19 (.A(n_0_114), .B(multiplicand[19]), .S(n_0_0_0), .Z(Res[19]));
   MUX2_X1 i_0_0_20 (.A(n_0_115), .B(multiplicand[20]), .S(n_0_0_0), .Z(Res[20]));
   MUX2_X1 i_0_0_21 (.A(n_0_116), .B(multiplicand[21]), .S(n_0_0_0), .Z(Res[21]));
   MUX2_X1 i_0_0_22 (.A(n_0_117), .B(multiplicand[22]), .S(n_0_0_0), .Z(Res[22]));
   MUX2_X1 i_0_0_23 (.A(n_0_118), .B(multiplicand[23]), .S(n_0_0_0), .Z(Res[23]));
   MUX2_X1 i_0_0_24 (.A(n_0_119), .B(multiplicand[24]), .S(n_0_0_0), .Z(Res[24]));
   MUX2_X1 i_0_0_25 (.A(n_0_120), .B(multiplicand[25]), .S(n_0_0_0), .Z(Res[25]));
   MUX2_X1 i_0_0_26 (.A(n_0_121), .B(multiplicand[26]), .S(n_0_0_0), .Z(Res[26]));
   MUX2_X1 i_0_0_27 (.A(n_0_122), .B(multiplicand[27]), .S(n_0_0_0), .Z(Res[27]));
   MUX2_X1 i_0_0_28 (.A(n_0_123), .B(multiplicand[28]), .S(n_0_0_0), .Z(Res[28]));
   MUX2_X1 i_0_0_29 (.A(n_0_124), .B(multiplicand[29]), .S(n_0_0_0), .Z(Res[29]));
   MUX2_X1 i_0_0_30 (.A(n_0_125), .B(multiplicand[30]), .S(n_0_0_0), .Z(Res[30]));
   MUX2_X1 i_0_0_31 (.A(n_0_126), .B(multiplicand[31]), .S(n_0_0_0), .Z(Res[31]));
   MUX2_X1 i_0_0_32 (.A(n_0_127), .B(accumulator[0]), .S(n_0_0_0), .Z(Res[32]));
   MUX2_X1 i_0_0_33 (.A(n_0_128), .B(accumulator[1]), .S(n_0_0_0), .Z(Res[33]));
   MUX2_X1 i_0_0_34 (.A(n_0_129), .B(accumulator[2]), .S(n_0_0_0), .Z(Res[34]));
   MUX2_X1 i_0_0_35 (.A(n_0_130), .B(accumulator[3]), .S(n_0_0_0), .Z(Res[35]));
   MUX2_X1 i_0_0_36 (.A(n_0_131), .B(accumulator[4]), .S(n_0_0_0), .Z(Res[36]));
   MUX2_X1 i_0_0_37 (.A(n_0_132), .B(accumulator[5]), .S(n_0_0_0), .Z(Res[37]));
   MUX2_X1 i_0_0_38 (.A(n_0_133), .B(accumulator[6]), .S(n_0_0_0), .Z(Res[38]));
   MUX2_X1 i_0_0_39 (.A(n_0_134), .B(accumulator[7]), .S(n_0_0_0), .Z(Res[39]));
   MUX2_X1 i_0_0_40 (.A(n_0_135), .B(accumulator[8]), .S(n_0_0_0), .Z(Res[40]));
   MUX2_X1 i_0_0_41 (.A(n_0_136), .B(accumulator[9]), .S(n_0_0_0), .Z(Res[41]));
   MUX2_X1 i_0_0_42 (.A(n_0_137), .B(accumulator[10]), .S(n_0_0_0), .Z(Res[42]));
   MUX2_X1 i_0_0_43 (.A(n_0_138), .B(accumulator[11]), .S(n_0_0_0), .Z(Res[43]));
   MUX2_X1 i_0_0_44 (.A(n_0_139), .B(accumulator[12]), .S(n_0_0_0), .Z(Res[44]));
   MUX2_X1 i_0_0_45 (.A(n_0_140), .B(accumulator[13]), .S(n_0_0_0), .Z(Res[45]));
   MUX2_X1 i_0_0_46 (.A(n_0_141), .B(accumulator[14]), .S(n_0_0_0), .Z(Res[46]));
   MUX2_X1 i_0_0_47 (.A(n_0_142), .B(accumulator[15]), .S(n_0_0_0), .Z(Res[47]));
   MUX2_X1 i_0_0_48 (.A(n_0_143), .B(accumulator[16]), .S(n_0_0_0), .Z(Res[48]));
   MUX2_X1 i_0_0_49 (.A(n_0_144), .B(accumulator[17]), .S(n_0_0_0), .Z(Res[49]));
   MUX2_X1 i_0_0_50 (.A(n_0_145), .B(accumulator[18]), .S(n_0_0_0), .Z(Res[50]));
   MUX2_X1 i_0_0_51 (.A(n_0_146), .B(accumulator[19]), .S(n_0_0_0), .Z(Res[51]));
   MUX2_X1 i_0_0_52 (.A(n_0_147), .B(accumulator[20]), .S(n_0_0_0), .Z(Res[52]));
   MUX2_X1 i_0_0_53 (.A(n_0_148), .B(accumulator[21]), .S(n_0_0_0), .Z(Res[53]));
   MUX2_X1 i_0_0_54 (.A(n_0_149), .B(accumulator[22]), .S(n_0_0_0), .Z(Res[54]));
   MUX2_X1 i_0_0_55 (.A(n_0_150), .B(accumulator[23]), .S(n_0_0_0), .Z(Res[55]));
   MUX2_X1 i_0_0_56 (.A(n_0_151), .B(accumulator[24]), .S(n_0_0_0), .Z(Res[56]));
   MUX2_X1 i_0_0_57 (.A(n_0_152), .B(accumulator[25]), .S(n_0_0_0), .Z(Res[57]));
   MUX2_X1 i_0_0_58 (.A(n_0_153), .B(accumulator[26]), .S(n_0_0_0), .Z(Res[58]));
   MUX2_X1 i_0_0_59 (.A(n_0_154), .B(accumulator[27]), .S(n_0_0_0), .Z(Res[59]));
   MUX2_X1 i_0_0_60 (.A(n_0_155), .B(accumulator[28]), .S(n_0_0_0), .Z(Res[60]));
   MUX2_X1 i_0_0_61 (.A(n_0_156), .B(accumulator[29]), .S(n_0_0_0), .Z(Res[61]));
   MUX2_X1 i_0_0_62 (.A(n_0_157), .B(accumulator[30]), .S(n_0_0_0), .Z(Res[62]));
   AND3_X1 i_0_0_63 (.A1(n_0_0_2), .A2(n_0_0_1), .A3(n_0_158), .ZN(Res[63]));
   NAND2_X1 i_0_0_64 (.A1(n_0_0_2), .A2(n_0_0_1), .ZN(n_0_0_0));
   XNOR2_X1 i_0_0_65 (.A(isNeg[1]), .B(n_0_0_101), .ZN(n_0_0_1));
   OR4_X1 i_0_0_66 (.A1(n_0_0_18), .A2(n_0_0_13), .A3(n_0_0_8), .A4(n_0_0_3), 
      .ZN(n_0_0_2));
   NAND4_X1 i_0_0_67 (.A1(n_0_0_7), .A2(n_0_0_6), .A3(n_0_0_5), .A4(n_0_0_4), 
      .ZN(n_0_0_3));
   NOR4_X1 i_0_0_68 (.A1(accumulator[15]), .A2(accumulator[11]), .A3(
      accumulator[10]), .A4(accumulator[9]), .ZN(n_0_0_4));
   NOR4_X1 i_0_0_69 (.A1(accumulator[14]), .A2(accumulator[13]), .A3(
      accumulator[12]), .A4(accumulator[8]), .ZN(n_0_0_5));
   NOR4_X1 i_0_0_70 (.A1(accumulator[3]), .A2(accumulator[2]), .A3(
      accumulator[1]), .A4(accumulator[0]), .ZN(n_0_0_6));
   NOR4_X1 i_0_0_71 (.A1(accumulator[7]), .A2(accumulator[6]), .A3(
      accumulator[5]), .A4(accumulator[4]), .ZN(n_0_0_7));
   NAND4_X1 i_0_0_72 (.A1(n_0_0_12), .A2(n_0_0_11), .A3(n_0_0_10), .A4(n_0_0_9), 
      .ZN(n_0_0_8));
   NOR4_X1 i_0_0_73 (.A1(accumulator[27]), .A2(accumulator[26]), .A3(
      accumulator[25]), .A4(accumulator[16]), .ZN(n_0_0_9));
   NOR4_X1 i_0_0_74 (.A1(accumulator[30]), .A2(accumulator[29]), .A3(
      accumulator[28]), .A4(accumulator[24]), .ZN(n_0_0_10));
   NOR4_X1 i_0_0_75 (.A1(accumulator[19]), .A2(accumulator[18]), .A3(
      accumulator[17]), .A4(Res[0]), .ZN(n_0_0_11));
   NOR4_X1 i_0_0_76 (.A1(accumulator[23]), .A2(accumulator[22]), .A3(
      accumulator[21]), .A4(accumulator[20]), .ZN(n_0_0_12));
   NAND4_X1 i_0_0_77 (.A1(n_0_0_17), .A2(n_0_0_16), .A3(n_0_0_15), .A4(n_0_0_14), 
      .ZN(n_0_0_13));
   NOR3_X1 i_0_0_78 (.A1(multiplicand[19]), .A2(multiplicand[18]), .A3(
      multiplicand[17]), .ZN(n_0_0_14));
   NOR4_X1 i_0_0_79 (.A1(multiplicand[23]), .A2(multiplicand[22]), .A3(
      multiplicand[21]), .A4(multiplicand[20]), .ZN(n_0_0_15));
   NOR4_X1 i_0_0_80 (.A1(multiplicand[27]), .A2(multiplicand[26]), .A3(
      multiplicand[25]), .A4(multiplicand[16]), .ZN(n_0_0_16));
   NOR4_X1 i_0_0_81 (.A1(multiplicand[30]), .A2(multiplicand[29]), .A3(
      multiplicand[28]), .A4(multiplicand[24]), .ZN(n_0_0_17));
   NAND4_X1 i_0_0_82 (.A1(n_0_0_22), .A2(n_0_0_21), .A3(n_0_0_20), .A4(n_0_0_19), 
      .ZN(n_0_0_18));
   NOR4_X1 i_0_0_83 (.A1(multiplicand[15]), .A2(multiplicand[11]), .A3(
      multiplicand[10]), .A4(multiplicand[9]), .ZN(n_0_0_19));
   NOR4_X1 i_0_0_84 (.A1(multiplicand[14]), .A2(multiplicand[13]), .A3(
      multiplicand[12]), .A4(multiplicand[8]), .ZN(n_0_0_20));
   NOR4_X1 i_0_0_85 (.A1(multiplicand[31]), .A2(multiplicand[3]), .A3(
      multiplicand[2]), .A4(multiplicand[1]), .ZN(n_0_0_21));
   NOR4_X1 i_0_0_86 (.A1(multiplicand[7]), .A2(multiplicand[6]), .A3(
      multiplicand[5]), .A4(multiplicand[4]), .ZN(n_0_0_22));
   OAI21_X1 i_0_0_87 (.A(n_0_0_97), .B1(n_0_0_106), .B2(counter[0]), .ZN(
      counter_in[0]));
   OAI21_X1 i_0_0_88 (.A(n_0_0_97), .B1(n_0_0_23), .B2(n_0_0_106), .ZN(
      counter_in[1]));
   XOR2_X1 i_0_0_89 (.A(counter[1]), .B(counter[0]), .Z(n_0_0_23));
   OAI21_X1 i_0_0_90 (.A(n_0_0_97), .B1(n_0_0_24), .B2(n_0_0_106), .ZN(
      counter_in[2]));
   AND2_X1 i_0_0_91 (.A1(n_0_0_30), .A2(n_0_0_25), .ZN(n_0_0_24));
   OAI21_X1 i_0_0_92 (.A(counter[2]), .B1(counter[1]), .B2(counter[0]), .ZN(
      n_0_0_25));
   OAI21_X1 i_0_0_93 (.A(n_0_0_97), .B1(n_0_0_26), .B2(n_0_0_106), .ZN(
      counter_in[3]));
   XOR2_X1 i_0_0_94 (.A(counter[3]), .B(n_0_0_30), .Z(n_0_0_26));
   OAI21_X1 i_0_0_95 (.A(n_0_0_97), .B1(n_0_0_27), .B2(n_0_0_106), .ZN(
      counter_in[4]));
   XOR2_X1 i_0_0_96 (.A(counter[4]), .B(n_0_0_29), .Z(n_0_0_27));
   OR2_X1 i_0_0_97 (.A1(reset), .A2(n_0_0_28), .ZN(n_0_160));
   OR2_X1 i_0_0_98 (.A1(n_0_0_28), .A2(n_0_258), .ZN(n_0_161));
   NOR3_X1 i_0_0_99 (.A1(n_0_0_29), .A2(ready), .A3(counter[4]), .ZN(n_0_0_28));
   OR2_X1 i_0_0_100 (.A1(n_0_0_30), .A2(counter[3]), .ZN(n_0_0_29));
   OR3_X1 i_0_0_101 (.A1(counter[2]), .A2(counter[1]), .A3(counter[0]), .ZN(
      n_0_0_30));
   INV_X1 i_0_0_102 (.A(n_0_0_32), .ZN(multiplicand_in[1]));
   AOI222_X1 i_0_0_103 (.A1(multiplicand[2]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_65), .C1(n_0_0_62), .C2(B[1]), .ZN(n_0_0_32));
   INV_X1 i_0_0_106 (.A(n_0_0_33), .ZN(multiplicand_in[2]));
   AOI222_X1 i_0_0_107 (.A1(multiplicand[3]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_66), .C1(n_0_0_62), .C2(B[2]), .ZN(n_0_0_33));
   INV_X1 i_0_0_108 (.A(n_0_0_34), .ZN(multiplicand_in[3]));
   AOI222_X1 i_0_0_109 (.A1(multiplicand[4]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_67), .C1(n_0_0_62), .C2(B[3]), .ZN(n_0_0_34));
   INV_X1 i_0_0_110 (.A(n_0_0_35), .ZN(multiplicand_in[4]));
   AOI222_X1 i_0_0_111 (.A1(multiplicand[5]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_68), .C1(n_0_0_62), .C2(B[4]), .ZN(n_0_0_35));
   INV_X1 i_0_0_112 (.A(n_0_0_36), .ZN(multiplicand_in[5]));
   AOI222_X1 i_0_0_113 (.A1(multiplicand[6]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_69), .C1(n_0_0_62), .C2(B[5]), .ZN(n_0_0_36));
   INV_X1 i_0_0_114 (.A(n_0_0_37), .ZN(multiplicand_in[6]));
   AOI222_X1 i_0_0_115 (.A1(multiplicand[7]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_70), .C1(n_0_0_62), .C2(B[6]), .ZN(n_0_0_37));
   INV_X1 i_0_0_116 (.A(n_0_0_38), .ZN(multiplicand_in[7]));
   AOI222_X1 i_0_0_117 (.A1(multiplicand[8]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_71), .C1(n_0_0_62), .C2(B[7]), .ZN(n_0_0_38));
   INV_X1 i_0_0_118 (.A(n_0_0_39), .ZN(multiplicand_in[8]));
   AOI222_X1 i_0_0_119 (.A1(multiplicand[9]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_72), .C1(n_0_0_62), .C2(B[8]), .ZN(n_0_0_39));
   INV_X1 i_0_0_120 (.A(n_0_0_40), .ZN(multiplicand_in[9]));
   AOI222_X1 i_0_0_121 (.A1(multiplicand[10]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_73), .C1(n_0_0_62), .C2(B[9]), .ZN(n_0_0_40));
   INV_X1 i_0_0_122 (.A(n_0_0_41), .ZN(multiplicand_in[10]));
   AOI222_X1 i_0_0_123 (.A1(multiplicand[11]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_74), .C1(n_0_0_62), .C2(B[10]), .ZN(n_0_0_41));
   INV_X1 i_0_0_124 (.A(n_0_0_42), .ZN(multiplicand_in[11]));
   AOI222_X1 i_0_0_125 (.A1(multiplicand[12]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_75), .C1(n_0_0_62), .C2(B[11]), .ZN(n_0_0_42));
   INV_X1 i_0_0_126 (.A(n_0_0_43), .ZN(multiplicand_in[12]));
   AOI222_X1 i_0_0_127 (.A1(multiplicand[13]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_76), .C1(n_0_0_62), .C2(B[12]), .ZN(n_0_0_43));
   INV_X1 i_0_0_128 (.A(n_0_0_44), .ZN(multiplicand_in[13]));
   AOI222_X1 i_0_0_129 (.A1(multiplicand[14]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_77), .C1(n_0_0_62), .C2(B[13]), .ZN(n_0_0_44));
   INV_X1 i_0_0_130 (.A(n_0_0_45), .ZN(multiplicand_in[14]));
   AOI222_X1 i_0_0_131 (.A1(multiplicand[15]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_78), .C1(n_0_0_62), .C2(B[14]), .ZN(n_0_0_45));
   INV_X1 i_0_0_132 (.A(n_0_0_46), .ZN(multiplicand_in[15]));
   AOI222_X1 i_0_0_133 (.A1(multiplicand[16]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_79), .C1(n_0_0_62), .C2(B[15]), .ZN(n_0_0_46));
   INV_X1 i_0_0_134 (.A(n_0_0_47), .ZN(multiplicand_in[16]));
   AOI222_X1 i_0_0_135 (.A1(multiplicand[17]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_80), .C1(n_0_0_62), .C2(B[16]), .ZN(n_0_0_47));
   INV_X1 i_0_0_136 (.A(n_0_0_48), .ZN(multiplicand_in[17]));
   AOI222_X1 i_0_0_137 (.A1(multiplicand[18]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_81), .C1(n_0_0_62), .C2(B[17]), .ZN(n_0_0_48));
   INV_X1 i_0_0_138 (.A(n_0_0_49), .ZN(multiplicand_in[18]));
   AOI222_X1 i_0_0_139 (.A1(multiplicand[19]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_82), .C1(n_0_0_62), .C2(B[18]), .ZN(n_0_0_49));
   INV_X1 i_0_0_140 (.A(n_0_0_50), .ZN(multiplicand_in[19]));
   AOI222_X1 i_0_0_141 (.A1(multiplicand[20]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_83), .C1(n_0_0_62), .C2(B[19]), .ZN(n_0_0_50));
   INV_X1 i_0_0_142 (.A(n_0_0_51), .ZN(multiplicand_in[20]));
   AOI222_X1 i_0_0_143 (.A1(multiplicand[21]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_84), .C1(n_0_0_62), .C2(B[20]), .ZN(n_0_0_51));
   INV_X1 i_0_0_144 (.A(n_0_0_52), .ZN(multiplicand_in[21]));
   AOI222_X1 i_0_0_145 (.A1(multiplicand[22]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_85), .C1(n_0_0_62), .C2(B[21]), .ZN(n_0_0_52));
   INV_X1 i_0_0_146 (.A(n_0_0_53), .ZN(multiplicand_in[22]));
   AOI222_X1 i_0_0_147 (.A1(multiplicand[23]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_86), .C1(n_0_0_62), .C2(B[22]), .ZN(n_0_0_53));
   INV_X1 i_0_0_148 (.A(n_0_0_54), .ZN(multiplicand_in[23]));
   AOI222_X1 i_0_0_149 (.A1(multiplicand[24]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_87), .C1(n_0_0_62), .C2(B[23]), .ZN(n_0_0_54));
   INV_X1 i_0_0_150 (.A(n_0_0_55), .ZN(multiplicand_in[24]));
   AOI222_X1 i_0_0_151 (.A1(multiplicand[25]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_88), .C1(n_0_0_62), .C2(B[24]), .ZN(n_0_0_55));
   INV_X1 i_0_0_152 (.A(n_0_0_56), .ZN(multiplicand_in[25]));
   AOI222_X1 i_0_0_153 (.A1(multiplicand[26]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_89), .C1(n_0_0_62), .C2(B[25]), .ZN(n_0_0_56));
   INV_X1 i_0_0_154 (.A(n_0_0_57), .ZN(multiplicand_in[26]));
   AOI222_X1 i_0_0_155 (.A1(multiplicand[27]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_90), .C1(n_0_0_62), .C2(B[26]), .ZN(n_0_0_57));
   INV_X1 i_0_0_156 (.A(n_0_0_58), .ZN(multiplicand_in[27]));
   AOI222_X1 i_0_0_157 (.A1(multiplicand[28]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_91), .C1(n_0_0_62), .C2(B[27]), .ZN(n_0_0_58));
   INV_X1 i_0_0_158 (.A(n_0_0_59), .ZN(multiplicand_in[28]));
   AOI222_X1 i_0_0_159 (.A1(multiplicand[29]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_92), .C1(n_0_0_62), .C2(B[28]), .ZN(n_0_0_59));
   INV_X1 i_0_0_160 (.A(n_0_0_60), .ZN(multiplicand_in[29]));
   AOI222_X1 i_0_0_161 (.A1(multiplicand[30]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_93), .C1(n_0_0_62), .C2(B[29]), .ZN(n_0_0_60));
   INV_X1 i_0_0_162 (.A(n_0_0_61), .ZN(multiplicand_in[30]));
   AOI222_X1 i_0_0_163 (.A1(multiplicand[31]), .A2(n_0_0_108), .B1(n_0_0_64), 
      .B2(n_0_94), .C1(n_0_0_62), .C2(B[30]), .ZN(n_0_0_61));
   NOR2_X1 i_0_0_104 (.A1(n_0_0_97), .A2(B[31]), .ZN(n_0_0_62));
   INV_X1 i_0_0_165 (.A(n_0_0_63), .ZN(multiplicand_in[31]));
   AOI22_X1 i_0_0_166 (.A1(n_0_2), .A2(n_0_0_108), .B1(n_0_0_64), .B2(n_0_95), 
      .ZN(n_0_0_63));
   NOR2_X1 i_0_0_105 (.A1(n_0_0_102), .A2(n_0_0_97), .ZN(n_0_0_64));
   NOR2_X1 i_0_0_168 (.A1(n_0_0_103), .A2(reset), .ZN(n_0_162));
   INV_X1 i_0_0_169 (.A(n_0_0_65), .ZN(n_0_163));
   AOI22_X1 i_0_0_170 (.A1(n_0_34), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[1]), 
      .ZN(n_0_0_65));
   INV_X1 i_0_0_171 (.A(n_0_0_66), .ZN(n_0_164));
   AOI22_X1 i_0_0_172 (.A1(n_0_35), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[2]), 
      .ZN(n_0_0_66));
   INV_X1 i_0_0_173 (.A(n_0_0_67), .ZN(n_0_165));
   AOI22_X1 i_0_0_174 (.A1(n_0_36), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[3]), 
      .ZN(n_0_0_67));
   INV_X1 i_0_0_175 (.A(n_0_0_68), .ZN(n_0_166));
   AOI22_X1 i_0_0_176 (.A1(n_0_37), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[4]), 
      .ZN(n_0_0_68));
   INV_X1 i_0_0_177 (.A(n_0_0_69), .ZN(n_0_167));
   AOI22_X1 i_0_0_178 (.A1(n_0_38), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[5]), 
      .ZN(n_0_0_69));
   INV_X1 i_0_0_179 (.A(n_0_0_70), .ZN(n_0_168));
   AOI22_X1 i_0_0_180 (.A1(n_0_39), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[6]), 
      .ZN(n_0_0_70));
   INV_X1 i_0_0_181 (.A(n_0_0_71), .ZN(n_0_169));
   AOI22_X1 i_0_0_182 (.A1(n_0_40), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[7]), 
      .ZN(n_0_0_71));
   INV_X1 i_0_0_183 (.A(n_0_0_72), .ZN(n_0_170));
   AOI22_X1 i_0_0_184 (.A1(n_0_41), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[8]), 
      .ZN(n_0_0_72));
   INV_X1 i_0_0_185 (.A(n_0_0_73), .ZN(n_0_171));
   AOI22_X1 i_0_0_186 (.A1(n_0_42), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[9]), 
      .ZN(n_0_0_73));
   INV_X1 i_0_0_187 (.A(n_0_0_74), .ZN(n_0_172));
   AOI22_X1 i_0_0_188 (.A1(n_0_43), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[10]), 
      .ZN(n_0_0_74));
   INV_X1 i_0_0_189 (.A(n_0_0_75), .ZN(n_0_173));
   AOI22_X1 i_0_0_190 (.A1(n_0_44), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[11]), 
      .ZN(n_0_0_75));
   INV_X1 i_0_0_191 (.A(n_0_0_76), .ZN(n_0_174));
   AOI22_X1 i_0_0_192 (.A1(n_0_45), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[12]), 
      .ZN(n_0_0_76));
   INV_X1 i_0_0_193 (.A(n_0_0_77), .ZN(n_0_175));
   AOI22_X1 i_0_0_194 (.A1(n_0_46), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[13]), 
      .ZN(n_0_0_77));
   INV_X1 i_0_0_195 (.A(n_0_0_78), .ZN(n_0_176));
   AOI22_X1 i_0_0_196 (.A1(n_0_47), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[14]), 
      .ZN(n_0_0_78));
   INV_X1 i_0_0_164 (.A(n_0_0_79), .ZN(n_0_177));
   AOI22_X1 i_0_0_167 (.A1(n_0_48), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[15]), 
      .ZN(n_0_0_79));
   INV_X1 i_0_0_199 (.A(n_0_0_80), .ZN(n_0_178));
   AOI22_X1 i_0_0_200 (.A1(n_0_49), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[16]), 
      .ZN(n_0_0_80));
   INV_X1 i_0_0_201 (.A(n_0_0_81), .ZN(n_0_179));
   AOI22_X1 i_0_0_202 (.A1(n_0_50), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[17]), 
      .ZN(n_0_0_81));
   INV_X1 i_0_0_203 (.A(n_0_0_82), .ZN(n_0_180));
   AOI22_X1 i_0_0_204 (.A1(n_0_51), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[18]), 
      .ZN(n_0_0_82));
   INV_X1 i_0_0_205 (.A(n_0_0_83), .ZN(n_0_181));
   AOI22_X1 i_0_0_206 (.A1(n_0_52), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[19]), 
      .ZN(n_0_0_83));
   INV_X1 i_0_0_207 (.A(n_0_0_84), .ZN(n_0_182));
   AOI22_X1 i_0_0_208 (.A1(n_0_53), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[20]), 
      .ZN(n_0_0_84));
   INV_X1 i_0_0_209 (.A(n_0_0_85), .ZN(n_0_183));
   AOI22_X1 i_0_0_210 (.A1(n_0_54), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[21]), 
      .ZN(n_0_0_85));
   INV_X1 i_0_0_211 (.A(n_0_0_86), .ZN(n_0_184));
   AOI22_X1 i_0_0_212 (.A1(n_0_55), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[22]), 
      .ZN(n_0_0_86));
   INV_X1 i_0_0_213 (.A(n_0_0_87), .ZN(n_0_185));
   AOI22_X1 i_0_0_214 (.A1(n_0_56), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[23]), 
      .ZN(n_0_0_87));
   INV_X1 i_0_0_215 (.A(n_0_0_88), .ZN(n_0_186));
   AOI22_X1 i_0_0_216 (.A1(n_0_57), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[24]), 
      .ZN(n_0_0_88));
   INV_X1 i_0_0_217 (.A(n_0_0_89), .ZN(n_0_187));
   AOI22_X1 i_0_0_218 (.A1(n_0_58), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[25]), 
      .ZN(n_0_0_89));
   INV_X1 i_0_0_219 (.A(n_0_0_90), .ZN(n_0_188));
   AOI22_X1 i_0_0_220 (.A1(n_0_59), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[26]), 
      .ZN(n_0_0_90));
   INV_X1 i_0_0_221 (.A(n_0_0_91), .ZN(n_0_189));
   AOI22_X1 i_0_0_222 (.A1(n_0_60), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[27]), 
      .ZN(n_0_0_91));
   INV_X1 i_0_0_223 (.A(n_0_0_92), .ZN(n_0_190));
   AOI22_X1 i_0_0_224 (.A1(n_0_61), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[28]), 
      .ZN(n_0_0_92));
   INV_X1 i_0_0_225 (.A(n_0_0_93), .ZN(n_0_191));
   AOI22_X1 i_0_0_226 (.A1(n_0_62), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[29]), 
      .ZN(n_0_0_93));
   INV_X1 i_0_0_227 (.A(n_0_0_94), .ZN(n_0_192));
   AOI22_X1 i_0_0_228 (.A1(n_0_63), .A2(n_0_0_96), .B1(n_0_0_95), .B2(A[30]), 
      .ZN(n_0_0_94));
   AOI21_X1 i_0_0_197 (.A(reset), .B1(A[31]), .B2(n_0_0_107), .ZN(n_0_0_95));
   NOR2_X1 i_0_0_198 (.A1(n_0_0_104), .A2(n_0_0_97), .ZN(n_0_0_96));
   NOR3_X1 i_0_0_232 (.A1(reset), .A2(n_0_0_98), .A3(n_0_0_104), .ZN(n_0_193));
   NOR2_X1 i_0_0_233 (.A1(n_0_0_100), .A2(n_0_64), .ZN(n_0_0_98));
   AND2_X1 i_0_0_234 (.A1(n_0_3), .A2(n_0_0_108), .ZN(n_0_194));
   AND2_X1 i_0_0_235 (.A1(n_0_4), .A2(n_0_0_108), .ZN(n_0_195));
   AND2_X1 i_0_0_236 (.A1(n_0_5), .A2(n_0_0_108), .ZN(n_0_196));
   AND2_X1 i_0_0_237 (.A1(n_0_6), .A2(n_0_0_108), .ZN(n_0_197));
   AND2_X1 i_0_0_238 (.A1(n_0_7), .A2(n_0_0_108), .ZN(n_0_198));
   AND2_X1 i_0_0_239 (.A1(n_0_8), .A2(n_0_0_108), .ZN(n_0_199));
   AND2_X1 i_0_0_240 (.A1(n_0_9), .A2(n_0_0_108), .ZN(n_0_200));
   AND2_X1 i_0_0_241 (.A1(n_0_10), .A2(n_0_0_108), .ZN(n_0_201));
   AND2_X1 i_0_0_242 (.A1(n_0_11), .A2(n_0_0_108), .ZN(n_0_202));
   AND2_X1 i_0_0_243 (.A1(n_0_12), .A2(n_0_0_108), .ZN(n_0_203));
   AND2_X1 i_0_0_244 (.A1(n_0_13), .A2(n_0_0_108), .ZN(n_0_204));
   AND2_X1 i_0_0_245 (.A1(n_0_14), .A2(n_0_0_108), .ZN(n_0_205));
   AND2_X1 i_0_0_246 (.A1(n_0_15), .A2(n_0_0_108), .ZN(n_0_206));
   AND2_X1 i_0_0_247 (.A1(n_0_16), .A2(n_0_0_108), .ZN(n_0_207));
   AND2_X1 i_0_0_248 (.A1(n_0_17), .A2(n_0_0_108), .ZN(n_0_208));
   AND2_X1 i_0_0_249 (.A1(n_0_18), .A2(n_0_0_108), .ZN(n_0_209));
   AND2_X1 i_0_0_250 (.A1(n_0_19), .A2(n_0_0_108), .ZN(n_0_210));
   AND2_X1 i_0_0_251 (.A1(n_0_20), .A2(n_0_0_108), .ZN(n_0_211));
   AND2_X1 i_0_0_252 (.A1(n_0_21), .A2(n_0_0_108), .ZN(n_0_212));
   AND2_X1 i_0_0_253 (.A1(n_0_22), .A2(n_0_0_108), .ZN(n_0_213));
   AND2_X1 i_0_0_254 (.A1(n_0_23), .A2(n_0_0_108), .ZN(n_0_214));
   AND2_X1 i_0_0_255 (.A1(n_0_24), .A2(n_0_0_108), .ZN(n_0_215));
   AND2_X1 i_0_0_256 (.A1(n_0_25), .A2(n_0_0_108), .ZN(n_0_216));
   AND2_X1 i_0_0_257 (.A1(n_0_26), .A2(n_0_0_108), .ZN(n_0_217));
   AND2_X1 i_0_0_258 (.A1(n_0_27), .A2(n_0_0_108), .ZN(n_0_218));
   AND2_X1 i_0_0_259 (.A1(n_0_28), .A2(n_0_0_108), .ZN(n_0_219));
   AND2_X1 i_0_0_260 (.A1(n_0_29), .A2(n_0_0_108), .ZN(n_0_220));
   AND2_X1 i_0_0_261 (.A1(n_0_30), .A2(n_0_0_108), .ZN(n_0_221));
   AND2_X1 i_0_0_262 (.A1(n_0_31), .A2(n_0_0_108), .ZN(n_0_222));
   AND2_X1 i_0_0_263 (.A1(n_0_32), .A2(n_0_0_108), .ZN(n_0_223));
   AND2_X1 i_0_0_264 (.A1(n_0_33), .A2(n_0_0_108), .ZN(n_0_224));
   AND2_X1 i_0_0_266 (.A1(multiplier[0]), .A2(Res[0]), .ZN(n_0_225));
   AND2_X1 i_0_0_267 (.A1(multiplier[1]), .A2(Res[0]), .ZN(n_0_226));
   AND2_X1 i_0_0_268 (.A1(multiplier[2]), .A2(Res[0]), .ZN(n_0_227));
   AND2_X1 i_0_0_269 (.A1(multiplier[3]), .A2(Res[0]), .ZN(n_0_228));
   AND2_X1 i_0_0_270 (.A1(multiplier[4]), .A2(Res[0]), .ZN(n_0_229));
   AND2_X1 i_0_0_271 (.A1(multiplier[5]), .A2(Res[0]), .ZN(n_0_230));
   AND2_X1 i_0_0_272 (.A1(multiplier[6]), .A2(Res[0]), .ZN(n_0_231));
   AND2_X1 i_0_0_273 (.A1(multiplier[7]), .A2(Res[0]), .ZN(n_0_232));
   AND2_X1 i_0_0_274 (.A1(multiplier[8]), .A2(Res[0]), .ZN(n_0_233));
   AND2_X1 i_0_0_275 (.A1(multiplier[9]), .A2(Res[0]), .ZN(n_0_234));
   AND2_X1 i_0_0_276 (.A1(multiplier[10]), .A2(Res[0]), .ZN(n_0_235));
   AND2_X1 i_0_0_277 (.A1(multiplier[11]), .A2(Res[0]), .ZN(n_0_236));
   AND2_X1 i_0_0_278 (.A1(multiplier[12]), .A2(Res[0]), .ZN(n_0_237));
   AND2_X1 i_0_0_279 (.A1(multiplier[13]), .A2(Res[0]), .ZN(n_0_238));
   AND2_X1 i_0_0_280 (.A1(multiplier[14]), .A2(Res[0]), .ZN(n_0_239));
   AND2_X1 i_0_0_281 (.A1(multiplier[15]), .A2(Res[0]), .ZN(n_0_240));
   AND2_X1 i_0_0_282 (.A1(multiplier[16]), .A2(Res[0]), .ZN(n_0_241));
   AND2_X1 i_0_0_283 (.A1(multiplier[17]), .A2(Res[0]), .ZN(n_0_242));
   AND2_X1 i_0_0_284 (.A1(multiplier[18]), .A2(Res[0]), .ZN(n_0_243));
   AND2_X1 i_0_0_285 (.A1(multiplier[19]), .A2(Res[0]), .ZN(n_0_244));
   AND2_X1 i_0_0_286 (.A1(multiplier[20]), .A2(Res[0]), .ZN(n_0_245));
   AND2_X1 i_0_0_287 (.A1(multiplier[21]), .A2(Res[0]), .ZN(n_0_246));
   AND2_X1 i_0_0_288 (.A1(multiplier[22]), .A2(Res[0]), .ZN(n_0_247));
   AND2_X1 i_0_0_289 (.A1(multiplier[23]), .A2(Res[0]), .ZN(n_0_248));
   AND2_X1 i_0_0_290 (.A1(multiplier[24]), .A2(Res[0]), .ZN(n_0_249));
   AND2_X1 i_0_0_291 (.A1(multiplier[25]), .A2(Res[0]), .ZN(n_0_250));
   AND2_X1 i_0_0_292 (.A1(multiplier[26]), .A2(Res[0]), .ZN(n_0_251));
   AND2_X1 i_0_0_293 (.A1(multiplier[27]), .A2(Res[0]), .ZN(n_0_252));
   AND2_X1 i_0_0_294 (.A1(multiplier[28]), .A2(Res[0]), .ZN(n_0_253));
   AND2_X1 i_0_0_295 (.A1(multiplier[29]), .A2(Res[0]), .ZN(n_0_254));
   AND2_X1 i_0_0_296 (.A1(multiplier[30]), .A2(Res[0]), .ZN(n_0_255));
   AND2_X1 i_0_0_297 (.A1(multiplier[31]), .A2(Res[0]), .ZN(n_0_256));
   OR3_X1 i_0_0_229 (.A1(n_0_0_105), .A2(reset), .A3(enable), .ZN(n_0_257));
   NOR2_X1 i_0_0_230 (.A1(n_0_0_102), .A2(reset), .ZN(isNeg_in[0]));
   NOR2_X1 i_0_0_300 (.A1(n_0_0_104), .A2(reset), .ZN(isNeg_in[1]));
   OR2_X1 i_0_0_231 (.A1(reset), .A2(n_0_0_107), .ZN(n_0_258));
   INV_X1 i_0_0_265 (.A(isNeg[0]), .ZN(n_0_0_101));
   INV_X1 i_0_0_298 (.A(B[31]), .ZN(n_0_0_102));
   INV_X1 i_0_0_305 (.A(A[0]), .ZN(n_0_0_103));
   INV_X1 i_0_0_299 (.A(A[31]), .ZN(n_0_0_104));
   INV_X1 i_0_0_301 (.A(ready), .ZN(n_0_0_105));
   INV_X1 i_0_0_302 (.A(n_0_0_108), .ZN(n_0_0_106));
   INV_X1 i_0_0_303 (.A(n_0_0_100), .ZN(n_0_0_107));
   INV_X1 i_0_0_304 (.A(n_0_0_31), .ZN(multiplicand_in[0]));
   AOI22_X1 i_0_0_306 (.A1(multiplicand[1]), .A2(n_0_0_108), .B1(B[0]), .B2(
      n_0_0_99), .ZN(n_0_0_31));
   INV_X1 i_0_0_307 (.A(n_0_0_99), .ZN(n_0_0_97));
   NOR2_X1 i_0_0_308 (.A1(reset), .A2(n_0_0_100), .ZN(n_0_0_99));
   NAND2_X1 i_0_0_309 (.A1(ready), .A2(enable), .ZN(n_0_0_100));
   NOR2_X1 i_0_0_310 (.A1(ready), .A2(reset), .ZN(n_0_0_108));
endmodule
