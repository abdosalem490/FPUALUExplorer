
// 	Thu Dec 22 21:48:58 2022
//	vlsi
//	192.168.126.129

module datapath__0_78 (M_multiplied, p_0, M_resultTruncated);

output [22:0] M_resultTruncated;
input M_multiplied;
input [22:0] p_0;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;


XOR2_X1 i_22 (.Z (M_resultTruncated[22]), .A (p_0[22]), .B (n_21));
HA_X1 i_21 (.CO (n_21), .S (M_resultTruncated[21]), .A (p_0[21]), .B (n_20));
HA_X1 i_20 (.CO (n_20), .S (M_resultTruncated[20]), .A (p_0[20]), .B (n_19));
HA_X1 i_19 (.CO (n_19), .S (M_resultTruncated[19]), .A (p_0[19]), .B (n_18));
HA_X1 i_18 (.CO (n_18), .S (M_resultTruncated[18]), .A (p_0[18]), .B (n_17));
HA_X1 i_17 (.CO (n_17), .S (M_resultTruncated[17]), .A (p_0[17]), .B (n_16));
HA_X1 i_16 (.CO (n_16), .S (M_resultTruncated[16]), .A (p_0[16]), .B (n_15));
HA_X1 i_15 (.CO (n_15), .S (M_resultTruncated[15]), .A (p_0[15]), .B (n_14));
HA_X1 i_14 (.CO (n_14), .S (M_resultTruncated[14]), .A (p_0[14]), .B (n_13));
HA_X1 i_13 (.CO (n_13), .S (M_resultTruncated[13]), .A (p_0[13]), .B (n_12));
HA_X1 i_12 (.CO (n_12), .S (M_resultTruncated[12]), .A (p_0[12]), .B (n_11));
HA_X1 i_11 (.CO (n_11), .S (M_resultTruncated[11]), .A (p_0[11]), .B (n_10));
HA_X1 i_10 (.CO (n_10), .S (M_resultTruncated[10]), .A (p_0[10]), .B (n_9));
HA_X1 i_9 (.CO (n_9), .S (M_resultTruncated[9]), .A (p_0[9]), .B (n_8));
HA_X1 i_8 (.CO (n_8), .S (M_resultTruncated[8]), .A (p_0[8]), .B (n_7));
HA_X1 i_7 (.CO (n_7), .S (M_resultTruncated[7]), .A (p_0[7]), .B (n_6));
HA_X1 i_6 (.CO (n_6), .S (M_resultTruncated[6]), .A (p_0[6]), .B (n_5));
HA_X1 i_5 (.CO (n_5), .S (M_resultTruncated[5]), .A (p_0[5]), .B (n_4));
HA_X1 i_4 (.CO (n_4), .S (M_resultTruncated[4]), .A (p_0[4]), .B (n_3));
HA_X1 i_3 (.CO (n_3), .S (M_resultTruncated[3]), .A (p_0[3]), .B (n_2));
HA_X1 i_2 (.CO (n_2), .S (M_resultTruncated[2]), .A (p_0[2]), .B (n_1));
HA_X1 i_1 (.CO (n_1), .S (M_resultTruncated[1]), .A (p_0[1]), .B (n_0));
HA_X1 i_0 (.CO (n_0), .S (M_resultTruncated[0]), .A (M_multiplied), .B (p_0[0]));

endmodule //datapath__0_78

module datapath__0_67 (p_0, p_1, p_2, p_3, p_4, p_5, p_6, p_7, p_8, p_9, p_10, p_11, 
    p_12, p_13, p_14, p_15, \aggregated_res[14] );

output [63:0] \aggregated_res[14] ;
input [63:0] p_0;
input [63:0] p_10;
input [63:0] p_11;
input [63:0] p_12;
input [63:0] p_13;
input [63:0] p_14;
input [63:0] p_15;
input [63:0] p_1;
input [63:0] p_2;
input [63:0] p_3;
input [63:0] p_4;
input [63:0] p_5;
input [63:0] p_6;
input [63:0] p_7;
input [63:0] p_8;
input [63:0] p_9;
wire n_117;
wire n_116;
wire n_179;
wire n_661;
wire n_665;
wire n_662;
wire n_198;
wire n_201;
wire n_209;
wire n_786;
wire n_203;
wire n_567;
wire n_563;
wire n_489;
wire n_269;
wire n_405;
wire n_570;
wire n_564;
wire n_485;
wire n_566;
wire n_277;
wire n_491;
wire n_281;
wire n_487;
wire n_407;
wire n_409;
wire n_552;
wire n_573;
wire n_545;
wire n_571;
wire n_574;
wire n_568;
wire n_565;
wire n_557;
wire n_581;
wire n_580;
wire n_626;
wire n_627;
wire n_624;
wire n_652;
wire n_621;
wire n_633;
wire n_593;
wire n_582;
wire n_739;
wire n_630;
wire n_660;
wire n_634;
wire n_631;
wire n_685;
wire n_596;
wire n_684;
wire n_594;
wire n_708;
wire n_690;
wire n_689;
wire n_643;
wire n_675;
wire n_732;
wire n_604;
wire n_731;
wire n_602;
wire n_754;
wire n_737;
wire n_736;
wire n_703;
wire n_722;
wire n_781;
wire n_775;
wire n_611;
wire n_610;
wire n_749;
wire n_765;
wire n_777;
wire n_774;
wire n_779;
wire n_205;
wire n_207;
wire n_211;
wire n_131;
wire n_130;
wire n_129;
wire n_128;
wire n_115;
wire n_135;
wire n_134;
wire n_139;
wire n_138;
wire n_102;
wire n_100;
wire n_98;
wire n_107;
wire n_106;
wire n_99;
wire n_105;
wire n_121;
wire n_120;
wire n_91;
wire n_104;
wire n_93;
wire n_109;
wire n_108;
wire n_125;
wire n_124;
wire n_113;
wire n_119;
wire n_132;
wire n_137;
wire n_136;
wire n_114;
wire n_112;
wire n_118;
wire n_123;
wire n_122;
wire n_141;
wire n_140;
wire n_143;
wire n_142;
wire n_145;
wire n_144;
wire n_153;
wire n_152;
wire n_157;
wire n_156;
wire n_150;
wire n_148;
wire n_146;
wire n_155;
wire n_154;
wire n_159;
wire n_158;
wire n_161;
wire n_160;
wire n_163;
wire n_162;
wire n_147;
wire n_151;
wire n_171;
wire n_170;
wire n_175;
wire n_174;
wire n_168;
wire n_166;
wire n_164;
wire n_173;
wire n_172;
wire n_177;
wire n_176;
wire n_213;
wire n_178;
wire n_103;
wire n_101;
wire n_127;
wire n_126;
wire n_75;
wire n_73;
wire n_77;
wire n_90;
wire n_61;
wire n_65;
wire n_76;
wire n_79;
wire n_78;
wire n_74;
wire n_72;
wire n_67;
wire n_81;
wire n_80;
wire n_95;
wire n_94;
wire n_89;
wire n_87;
wire n_85;
wire n_88;
wire n_86;
wire n_84;
wire n_92;
wire n_111;
wire n_110;
wire n_60;
wire n_53;
wire n_52;
wire n_64;
wire n_63;
wire n_62;
wire n_35;
wire n_33;
wire n_45;
wire n_44;
wire n_51;
wire n_50;
wire n_57;
wire n_56;
wire n_69;
wire n_68;
wire n_43;
wire n_41;
wire n_55;
wire n_54;
wire n_66;
wire n_83;
wire n_82;
wire n_97;
wire n_96;
wire n_71;
wire n_70;
wire n_42;
wire n_40;
wire n_34;
wire n_32;
wire n_47;
wire n_46;
wire n_59;
wire n_58;
wire n_27;
wire n_25;
wire n_37;
wire n_36;
wire n_29;
wire n_39;
wire n_38;
wire n_49;
wire n_48;
wire n_24;
wire n_15;
wire n_20;
wire n_18;
wire n_23;
wire n_22;
wire n_31;
wire n_30;
wire n_19;
wire n_21;
wire n_26;
wire n_28;
wire n_13;
wire n_12;
wire n_5;
wire n_7;
wire n_11;
wire n_10;
wire n_9;
wire n_14;
wire n_17;
wire n_16;
wire n_8;
wire n_4;
wire n_3;
wire n_6;
wire n_2;
wire n_1;
wire n_0;
wire n_183;
wire n_182;
wire n_181;
wire n_180;
wire n_133;
wire n_193;
wire n_192;
wire n_149;
wire n_169;
wire n_187;
wire n_186;
wire n_185;
wire n_184;
wire n_191;
wire n_190;
wire n_167;
wire n_165;
wire n_189;
wire n_188;
wire n_195;
wire n_194;
wire n_197;
wire n_196;
wire n_199;
wire n_215;
wire n_217;
wire n_208;
wire n_219;
wire n_214;
wire n_240;
wire n_206;
wire n_241;
wire n_210;
wire n_260;
wire n_204;
wire n_261;
wire n_202;
wire n_263;
wire n_200;
wire n_265;
wire n_212;
wire n_267;
wire n_216;
wire n_218;
wire n_273;
wire n_271;
wire n_275;
wire n_279;
wire n_282;
wire n_369;
wire n_367;
wire n_283;
wire n_323;
wire n_390;
wire n_331;
wire n_327;
wire n_333;
wire n_325;
wire n_329;
wire n_339;
wire n_335;
wire n_362;
wire n_337;
wire n_365;
wire n_361;
wire n_359;
wire n_340;
wire n_341;
wire n_351;
wire n_345;
wire n_353;
wire n_343;
wire n_355;
wire n_347;
wire n_349;
wire n_357;
wire n_358;
wire n_371;
wire n_391;
wire n_375;
wire n_404;
wire n_373;
wire n_226;
wire n_224;
wire n_222;
wire n_233;
wire n_232;
wire n_237;
wire n_236;
wire n_220;
wire n_230;
wire n_228;
wire n_235;
wire n_234;
wire n_239;
wire n_238;
wire n_221;
wire n_231;
wire n_229;
wire n_245;
wire n_244;
wire n_243;
wire n_242;
wire n_561;
wire n_253;
wire n_252;
wire n_247;
wire n_246;
wire n_558;
wire n_251;
wire n_250;
wire n_257;
wire n_256;
wire n_225;
wire n_223;
wire n_249;
wire n_248;
wire n_227;
wire n_255;
wire n_254;
wire n_259;
wire n_258;
wire n_411;
wire n_413;
wire n_268;
wire n_415;
wire n_276;
wire n_417;
wire n_262;
wire n_562;
wire n_418;
wire n_270;
wire n_554;
wire n_419;
wire n_274;
wire n_430;
wire n_266;
wire n_431;
wire n_264;
wire n_556;
wire n_442;
wire n_272;
wire n_445;
wire n_278;
wire n_447;
wire n_280;
wire n_451;
wire n_449;
wire n_462;
wire n_505;
wire n_502;
wire n_453;
wire n_494;
wire n_500;
wire n_455;
wire n_457;
wire n_503;
wire n_501;
wire n_470;
wire n_459;
wire n_461;
wire n_463;
wire n_478;
wire n_499;
wire n_471;
wire n_483;
wire n_481;
wire n_490;
wire n_291;
wire n_290;
wire n_309;
wire n_308;
wire n_553;
wire n_313;
wire n_312;
wire n_297;
wire n_296;
wire n_307;
wire n_306;
wire n_305;
wire n_304;
wire n_549;
wire n_315;
wire n_314;
wire n_319;
wire n_318;
wire n_507;
wire n_324;
wire n_550;
wire n_512;
wire n_330;
wire n_546;
wire n_515;
wire n_334;
wire n_289;
wire n_288;
wire n_287;
wire n_286;
wire n_285;
wire n_284;
wire n_311;
wire n_310;
wire n_517;
wire n_328;
wire n_522;
wire n_326;
wire n_525;
wire n_332;
wire n_551;
wire n_295;
wire n_294;
wire n_293;
wire n_292;
wire n_317;
wire n_316;
wire n_527;
wire n_336;
wire n_532;
wire n_338;
wire n_299;
wire n_298;
wire n_321;
wire n_320;
wire n_537;
wire n_535;
wire n_301;
wire n_300;
wire n_539;
wire n_322;
wire n_303;
wire n_302;
wire n_540;
wire n_583;
wire n_578;
wire n_577;
wire n_579;
wire n_543;
wire n_542;
wire n_569;
wire n_547;
wire n_576;
wire n_560;
wire n_555;
wire n_559;
wire n_572;
wire n_575;
wire n_584;
wire n_346;
wire n_585;
wire n_344;
wire n_586;
wire n_350;
wire n_587;
wire n_342;
wire n_548;
wire n_588;
wire n_348;
wire n_544;
wire n_589;
wire n_352;
wire n_590;
wire n_354;
wire n_591;
wire n_356;
wire n_595;
wire n_592;
wire n_598;
wire n_597;
wire n_601;
wire n_614;
wire n_613;
wire n_603;
wire n_599;
wire n_600;
wire n_607;
wire n_605;
wire n_612;
wire n_606;
wire n_608;
wire n_609;
wire n_615;
wire n_360;
wire n_541;
wire n_616;
wire n_368;
wire n_617;
wire n_364;
wire n_639;
wire n_618;
wire n_366;
wire n_619;
wire n_370;
wire n_620;
wire n_372;
wire n_374;
wire n_622;
wire n_623;
wire n_625;
wire n_628;
wire n_629;
wire n_379;
wire n_377;
wire n_397;
wire n_396;
wire n_378;
wire n_383;
wire n_382;
wire n_536;
wire n_401;
wire n_400;
wire n_376;
wire n_380;
wire n_385;
wire n_384;
wire n_387;
wire n_386;
wire n_389;
wire n_388;
wire n_381;
wire n_394;
wire n_392;
wire n_399;
wire n_398;
wire n_403;
wire n_402;
wire n_632;
wire n_635;
wire n_408;
wire n_636;
wire n_406;
wire n_637;
wire n_412;
wire n_395;
wire n_393;
wire n_538;
wire n_638;
wire n_410;
wire n_363;
wire n_534;
wire n_640;
wire n_414;
wire n_641;
wire n_416;
wire n_642;
wire n_663;
wire n_666;
wire n_646;
wire n_667;
wire n_664;
wire n_647;
wire n_644;
wire n_645;
wire n_653;
wire n_648;
wire n_649;
wire n_654;
wire n_650;
wire n_651;
wire n_656;
wire n_668;
wire n_658;
wire n_655;
wire n_657;
wire n_659;
wire n_425;
wire n_424;
wire n_429;
wire n_428;
wire n_423;
wire n_422;
wire n_421;
wire n_420;
wire n_531;
wire n_427;
wire n_426;
wire n_435;
wire n_434;
wire n_533;
wire n_437;
wire n_436;
wire n_433;
wire n_432;
wire n_529;
wire n_439;
wire n_438;
wire n_441;
wire n_440;
wire n_443;
wire n_669;
wire n_670;
wire n_444;
wire n_526;
wire n_671;
wire n_448;
wire n_530;
wire n_672;
wire n_446;
wire n_673;
wire n_450;
wire n_674;
wire n_452;
wire n_676;
wire n_677;
wire n_696;
wire n_694;
wire n_681;
wire n_678;
wire n_680;
wire n_679;
wire n_695;
wire n_683;
wire n_682;
wire n_692;
wire n_688;
wire n_686;
wire n_687;
wire n_691;
wire n_693;
wire n_697;
wire n_698;
wire n_454;
wire n_524;
wire n_699;
wire n_458;
wire n_528;
wire n_700;
wire n_456;
wire n_701;
wire n_460;
wire n_702;
wire n_704;
wire n_705;
wire n_706;
wire n_707;
wire n_709;
wire n_710;
wire n_711;
wire n_712;
wire n_713;
wire n_714;
wire n_715;
wire n_716;
wire n_717;
wire n_465;
wire n_464;
wire n_467;
wire n_466;
wire n_521;
wire n_469;
wire n_468;
wire n_473;
wire n_472;
wire n_523;
wire n_475;
wire n_474;
wire n_519;
wire n_477;
wire n_476;
wire n_479;
wire n_718;
wire n_719;
wire n_480;
wire n_520;
wire n_516;
wire n_720;
wire n_482;
wire n_721;
wire n_484;
wire n_723;
wire n_724;
wire n_728;
wire n_725;
wire n_727;
wire n_744;
wire n_742;
wire n_726;
wire n_743;
wire n_730;
wire n_729;
wire n_740;
wire n_735;
wire n_733;
wire n_734;
wire n_738;
wire n_741;
wire n_745;
wire n_518;
wire n_746;
wire n_486;
wire n_514;
wire n_747;
wire n_488;
wire n_748;
wire n_750;
wire n_751;
wire n_752;
wire n_753;
wire n_755;
wire n_756;
wire n_757;
wire n_758;
wire n_759;
wire n_760;
wire n_761;
wire n_493;
wire n_492;
wire n_513;
wire n_509;
wire n_497;
wire n_496;
wire n_762;
wire n_498;
wire n_510;
wire n_506;
wire n_764;
wire n_763;
wire n_511;
wire n_495;
wire n_788;
wire n_766;
wire n_769;
wire n_785;
wire n_767;
wire n_789;
wire n_787;
wire n_768;
wire n_772;
wire n_770;
wire n_780;
wire n_771;
wire n_773;
wire n_783;
wire n_776;
wire n_778;
wire n_782;
wire n_784;
wire n_790;
wire n_508;
wire n_504;
wire n_792;
wire n_791;
wire n_793;
wire n_796;
wire n_804;
wire n_795;
wire n_794;
wire n_805;
wire n_803;
wire n_799;
wire n_797;
wire n_802;
wire n_798;
wire n_800;
wire n_801;
wire n_809;
wire n_806;
wire n_807;
wire n_808;
wire n_812;
wire n_810;
wire n_811;


NOR2_X1 i_585 (.ZN (n_812), .A1 (n_791), .A2 (n_764));
NOR2_X1 i_584 (.ZN (n_811), .A1 (n_805), .A2 (n_803));
AOI211_X1 i_583 (.ZN (n_810), .A (n_811), .B (n_799), .C1 (n_758), .C2 (n_797));
NOR2_X1 i_582 (.ZN (n_809), .A1 (n_812), .A2 (n_810));
XOR2_X1 i_581 (.Z (n_808), .A (p_10[47]), .B (p_11[47]));
XOR2_X1 i_580 (.Z (n_807), .A (n_796), .B (n_808));
XOR2_X1 i_579 (.Z (n_806), .A (n_792), .B (n_807));
XOR2_X2 i_578 (.Z (\aggregated_res[14] [47] ), .A (n_809), .B (n_806));
INV_X1 i_577 (.ZN (n_805), .A (n_791));
INV_X1 i_576 (.ZN (n_804), .A (p_10[45]));
INV_X1 i_575 (.ZN (n_803), .A (n_764));
OAI21_X1 i_574 (.ZN (n_802), .A (n_773), .B1 (n_762), .B2 (n_763));
AOI21_X1 i_573 (.ZN (n_801), .A (n_802), .B1 (n_759), .B2 (n_778));
INV_X1 i_572 (.ZN (n_800), .A (n_801));
OAI211_X1 i_571 (.ZN (n_799), .A (n_783), .B (n_800), .C1 (n_780), .C2 (n_784));
NOR2_X1 i_570 (.ZN (n_798), .A1 (n_721), .A2 (n_748));
NOR2_X1 i_569 (.ZN (n_797), .A1 (n_802), .A2 (n_798));
NOR2_X1 i_568 (.ZN (n_796), .A1 (p_10[46]), .A2 (p_11[46]));
AOI21_X1 i_567 (.ZN (n_795), .A (n_799), .B1 (n_758), .B2 (n_797));
OAI22_X1 i_566 (.ZN (n_794), .A1 (n_805), .A2 (n_764), .B1 (n_791), .B2 (n_803));
XNOR2_X1 i_565 (.ZN (\aggregated_res[14] [46] ), .A (n_795), .B (n_794));
OAI222_X1 i_564 (.ZN (n_508), .A1 (p_9[45]), .A2 (n_790), .B1 (n_804), .B2 (p_9[45])
    , .C1 (n_804), .C2 (n_790));
AOI21_X1 i_563 (.ZN (n_793), .A (n_796), .B1 (p_10[46]), .B2 (p_11[46]));
INV_X1 i_562 (.ZN (n_504), .A (n_793));
HA_X1 i_561 (.CO (n_792), .S (n_791), .A (n_508), .B (n_504));
INV_X1 i_560 (.ZN (n_790), .A (p_11[45]));
INV_X1 i_559 (.ZN (n_789), .A (p_10[44]));
INV_X1 i_558 (.ZN (n_788), .A (p_10[43]));
INV_X1 i_557 (.ZN (n_787), .A (p_9[44]));
INV_X1 i_556 (.ZN (n_785), .A (p_9[43]));
NOR2_X1 i_555 (.ZN (n_784), .A1 (n_762), .A2 (n_763));
NAND2_X1 i_554 (.ZN (n_783), .A1 (n_762), .A2 (n_763));
NOR2_X1 i_553 (.ZN (n_782), .A1 (n_721), .A2 (n_748));
AOI21_X1 i_552 (.ZN (n_781), .A (n_782), .B1 (n_761), .B2 (n_759));
NAND2_X1 i_551 (.ZN (n_780), .A1 (n_498), .A2 (n_495));
INV_X1 i_550 (.ZN (n_779), .A (n_780));
NAND2_X1 i_549 (.ZN (n_778), .A1 (n_765), .A2 (n_749));
INV_X1 i_548 (.ZN (n_777), .A (n_778));
NOR2_X1 i_547 (.ZN (n_776), .A1 (n_765), .A2 (n_749));
NOR2_X1 i_546 (.ZN (n_775), .A1 (n_777), .A2 (n_776));
NOR2_X1 i_545 (.ZN (n_774), .A1 (n_498), .A2 (n_495));
NOR2_X1 i_544 (.ZN (n_773), .A1 (n_776), .A2 (n_774));
OAI21_X1 i_543 (.ZN (n_772), .A (n_783), .B1 (n_762), .B2 (n_763));
OAI21_X1 i_542 (.ZN (n_771), .A (n_773), .B1 (n_781), .B2 (n_777));
NAND2_X1 i_541 (.ZN (n_770), .A1 (n_780), .A2 (n_771));
XNOR2_X1 i_540 (.ZN (\aggregated_res[14] [45] ), .A (n_772), .B (n_770));
NOR2_X1 i_539 (.ZN (n_769), .A1 (n_785), .A2 (p_8[45]));
INV_X1 i_538 (.ZN (n_768), .A (n_769));
AOI22_X1 i_537 (.ZN (n_513), .A1 (n_785), .A2 (p_8[45]), .B1 (n_788), .B2 (n_768));
NAND2_X1 i_536 (.ZN (n_510), .A1 (n_789), .A2 (n_787));
OAI21_X1 i_535 (.ZN (n_509), .A (n_510), .B1 (n_789), .B2 (n_787));
XOR2_X1 i_534 (.Z (n_767), .A (p_10[45]), .B (p_9[45]));
XNOR2_X1 i_533 (.ZN (n_506), .A (p_11[45]), .B (n_767));
AOI21_X1 i_532 (.ZN (n_766), .A (n_769), .B1 (n_785), .B2 (p_8[45]));
XNOR2_X1 i_531 (.ZN (n_511), .A (n_788), .B (n_766));
FA_X1 i_530 (.CO (n_495), .S (n_765), .A (n_511), .B (n_492), .CI (n_747));
FA_X1 i_529 (.CO (n_764), .S (n_763), .A (n_510), .B (n_506), .CI (n_497));
HA_X1 i_528 (.CO (n_762), .S (n_498), .A (n_493), .B (n_496));
FA_X1 i_527 (.CO (n_497), .S (n_496), .A (p_11[44]), .B (n_513), .CI (n_509));
FA_X1 i_526 (.CO (n_493), .S (n_492), .A (p_11[43]), .B (n_752), .CI (n_746));
INV_X1 i_525 (.ZN (n_761), .A (n_758));
XNOR2_X1 i_524 (.ZN (\aggregated_res[14] [42] ), .A (n_758), .B (n_760));
OAI21_X1 i_523 (.ZN (n_760), .A (n_759), .B1 (n_748), .B2 (n_721));
NAND2_X1 i_522 (.ZN (n_759), .A1 (n_748), .A2 (n_721));
OAI221_X2 i_521 (.ZN (n_758), .A (n_740), .B1 (n_741), .B2 (n_738), .C1 (n_755), .C2 (n_757));
AND3_X2 i_520 (.ZN (n_757), .A1 (n_756), .A2 (n_735), .A3 (n_716));
OAI22_X1 i_519 (.ZN (n_756), .A1 (n_711), .A2 (n_714), .B1 (n_674), .B2 (n_702));
OR3_X1 i_518 (.ZN (n_755), .A1 (n_754), .A2 (n_736), .A3 (n_741));
NOR2_X1 i_517 (.ZN (n_754), .A1 (n_723), .A2 (n_718));
OAI222_X1 i_516 (.ZN (n_518), .A1 (n_753), .A2 (n_745), .B1 (n_753), .B2 (p_7[45])
    , .C1 (p_7[45]), .C2 (n_745));
INV_X1 i_515 (.ZN (n_753), .A (p_8[41]));
OAI21_X1 i_514 (.ZN (n_514), .A (n_752), .B1 (n_750), .B2 (n_751));
NAND2_X1 i_513 (.ZN (n_752), .A1 (n_750), .A2 (n_751));
INV_X1 i_512 (.ZN (n_751), .A (p_9[42]));
INV_X1 i_511 (.ZN (n_750), .A (p_8[42]));
HA_X1 i_510 (.CO (n_749), .S (n_748), .A (n_720), .B (n_488));
FA_X1 i_509 (.CO (n_747), .S (n_488), .A (n_719), .B (n_486), .CI (n_514));
FA_X1 i_508 (.CO (n_746), .S (n_486), .A (p_10[42]), .B (p_11[42]), .CI (n_518));
INV_X1 i_507 (.ZN (n_745), .A (p_9[41]));
INV_X1 i_506 (.ZN (n_744), .A (p_8[40]));
INV_X1 i_505 (.ZN (n_743), .A (p_6[45]));
INV_X1 i_504 (.ZN (n_742), .A (p_7[40]));
NOR2_X1 i_503 (.ZN (n_741), .A1 (n_479), .A2 (n_484));
NAND2_X1 i_502 (.ZN (n_740), .A1 (n_479), .A2 (n_484));
NAND2_X1 i_501 (.ZN (n_738), .A1 (n_718), .A2 (n_723));
INV_X1 i_500 (.ZN (n_737), .A (n_738));
NOR2_X1 i_499 (.ZN (n_736), .A1 (n_722), .A2 (n_703));
NAND2_X1 i_498 (.ZN (n_735), .A1 (n_722), .A2 (n_703));
NAND2_X1 i_497 (.ZN (n_734), .A1 (n_715), .A2 (n_716));
OAI21_X1 i_496 (.ZN (n_733), .A (n_734), .B1 (n_702), .B2 (n_674));
INV_X1 i_495 (.ZN (n_732), .A (n_733));
AOI21_X1 i_494 (.ZN (n_731), .A (n_736), .B1 (n_735), .B2 (n_733));
OAI21_X1 i_493 (.ZN (n_730), .A (n_740), .B1 (n_479), .B2 (n_484));
OAI22_X1 i_492 (.ZN (n_729), .A1 (n_718), .A2 (n_723), .B1 (n_737), .B2 (n_731));
XOR2_X2 i_491 (.Z (\aggregated_res[14] [41] ), .A (n_730), .B (n_729));
NAND2_X1 i_490 (.ZN (n_728), .A1 (n_743), .A2 (p_7[39]));
OR2_X1 i_489 (.ZN (n_727), .A1 (n_743), .A2 (p_7[39]));
NAND2_X1 i_488 (.ZN (n_726), .A1 (n_728), .A2 (n_727));
XNOR2_X1 i_487 (.ZN (n_521), .A (p_8[39]), .B (n_726));
NAND2_X1 i_486 (.ZN (n_520), .A1 (n_744), .A2 (n_742));
OAI21_X1 i_485 (.ZN (n_519), .A (n_520), .B1 (n_744), .B2 (n_742));
NAND2_X1 i_484 (.ZN (n_725), .A1 (p_8[39]), .A2 (n_727));
NAND2_X1 i_483 (.ZN (n_523), .A1 (n_728), .A2 (n_725));
XOR2_X1 i_482 (.Z (n_724), .A (p_8[41]), .B (p_7[45]));
XNOR2_X1 i_481 (.ZN (n_516), .A (p_9[41]), .B (n_724));
FA_X1 i_480 (.CO (n_723), .S (n_722), .A (n_699), .B (n_468), .CI (n_701));
FA_X1 i_479 (.CO (n_721), .S (n_484), .A (n_475), .B (n_477), .CI (n_482));
FA_X1 i_478 (.CO (n_720), .S (n_482), .A (n_520), .B (n_480), .CI (n_516));
FA_X1 i_477 (.CO (n_719), .S (n_480), .A (p_10[41]), .B (p_11[41]), .CI (n_473));
HA_X1 i_476 (.CO (n_479), .S (n_718), .A (n_469), .B (n_476));
FA_X1 i_475 (.CO (n_477), .S (n_476), .A (n_519), .B (n_467), .CI (n_474));
FA_X1 i_474 (.CO (n_475), .S (n_474), .A (n_465), .B (n_523), .CI (n_472));
FA_X1 i_473 (.CO (n_473), .S (n_472), .A (p_9[40]), .B (p_10[40]), .CI (p_11[40]));
FA_X1 i_472 (.CO (n_469), .S (n_468), .A (n_464), .B (n_521), .CI (n_466));
FA_X1 i_471 (.CO (n_467), .S (n_466), .A (n_698), .B (n_707), .CI (n_700));
FA_X1 i_470 (.CO (n_465), .S (n_464), .A (p_9[39]), .B (p_10[39]), .CI (p_11[39]));
XOR2_X1 i_469 (.Z (\aggregated_res[14] [38] ), .A (n_715), .B (n_717));
OAI21_X1 i_468 (.ZN (n_717), .A (n_716), .B1 (n_702), .B2 (n_674));
NAND2_X1 i_467 (.ZN (n_716), .A1 (n_702), .A2 (n_674));
NOR2_X1 i_466 (.ZN (n_715), .A1 (n_714), .A2 (n_711));
OAI221_X1 i_465 (.ZN (n_714), .A (n_692), .B1 (n_693), .B2 (n_691), .C1 (n_712), .C2 (n_713));
AND2_X1 i_464 (.ZN (n_713), .A1 (n_645), .A2 (n_688));
INV_X1 i_463 (.ZN (n_712), .A (n_709));
AOI21_X2 i_462 (.ZN (n_711), .A (n_710), .B1 (n_653), .B2 (n_648));
OAI21_X1 i_461 (.ZN (n_710), .A (n_709), .B1 (n_632), .B2 (n_642));
NOR3_X1 i_460 (.ZN (n_709), .A1 (n_708), .A2 (n_689), .A3 (n_693));
NOR2_X1 i_459 (.ZN (n_708), .A1 (n_676), .A2 (n_669));
OAI21_X1 i_458 (.ZN (n_524), .A (n_707), .B1 (n_705), .B2 (n_706));
NAND2_X1 i_457 (.ZN (n_707), .A1 (n_705), .A2 (n_706));
INV_X1 i_454 (.ZN (n_706), .A (p_7[38]));
INV_X1 i_453 (.ZN (n_705), .A (p_6[38]));
OAI222_X1 i_452 (.ZN (n_528), .A1 (n_704), .A2 (n_697), .B1 (n_704), .B2 (p_5[43])
    , .C1 (p_5[43]), .C2 (n_697));
INV_X1 i_451 (.ZN (n_704), .A (p_6[37]));
HA_X1 i_450 (.CO (n_703), .S (n_702), .A (n_458), .B (n_460));
FA_X1 i_449 (.CO (n_701), .S (n_460), .A (n_456), .B (n_671), .CI (n_673));
FA_X1 i_448 (.CO (n_700), .S (n_456), .A (p_11[38]), .B (n_670), .CI (n_528));
FA_X1 i_447 (.CO (n_699), .S (n_458), .A (n_672), .B (n_454), .CI (n_524));
FA_X1 i_446 (.CO (n_698), .S (n_454), .A (p_8[38]), .B (p_9[38]), .CI (p_10[38]));
INV_X1 i_445 (.ZN (n_697), .A (p_7[37]));
INV_X1 i_444 (.ZN (n_696), .A (p_6[36]));
INV_X1 i_443 (.ZN (n_695), .A (p_4[42]));
INV_X1 i_442 (.ZN (n_694), .A (p_5[36]));
NOR2_X1 i_441 (.ZN (n_693), .A1 (n_443), .A2 (n_452));
NAND2_X1 i_440 (.ZN (n_692), .A1 (n_443), .A2 (n_452));
NAND2_X1 i_439 (.ZN (n_691), .A1 (n_669), .A2 (n_676));
INV_X1 i_438 (.ZN (n_690), .A (n_691));
NOR2_X1 i_437 (.ZN (n_689), .A1 (n_675), .A2 (n_643));
NAND2_X1 i_436 (.ZN (n_688), .A1 (n_675), .A2 (n_643));
NAND2_X1 i_435 (.ZN (n_687), .A1 (n_647), .A2 (n_645));
OAI21_X1 i_434 (.ZN (n_686), .A (n_687), .B1 (n_632), .B2 (n_642));
INV_X1 i_433 (.ZN (n_685), .A (n_686));
AOI21_X1 i_432 (.ZN (n_684), .A (n_689), .B1 (n_688), .B2 (n_686));
OAI21_X1 i_431 (.ZN (n_683), .A (n_692), .B1 (n_443), .B2 (n_452));
OAI22_X1 i_430 (.ZN (n_682), .A1 (n_669), .A2 (n_676), .B1 (n_690), .B2 (n_684));
XOR2_X2 i_429 (.Z (\aggregated_res[14] [37] ), .A (n_683), .B (n_682));
NAND2_X1 i_428 (.ZN (n_681), .A1 (n_695), .A2 (p_5[35]));
OR2_X1 i_427 (.ZN (n_680), .A1 (n_695), .A2 (p_5[35]));
NAND2_X1 i_426 (.ZN (n_679), .A1 (n_681), .A2 (n_680));
XNOR2_X1 i_425 (.ZN (n_531), .A (p_6[35]), .B (n_679));
NAND2_X1 i_424 (.ZN (n_678), .A1 (p_6[35]), .A2 (n_680));
NAND2_X1 i_423 (.ZN (n_533), .A1 (n_681), .A2 (n_678));
NAND2_X1 i_422 (.ZN (n_530), .A1 (n_696), .A2 (n_694));
OAI21_X1 i_421 (.ZN (n_529), .A (n_530), .B1 (n_696), .B2 (n_694));
XOR2_X1 i_420 (.Z (n_677), .A (p_6[37]), .B (p_5[43]));
XNOR2_X1 i_419 (.ZN (n_526), .A (p_7[37]), .B (n_677));
FA_X1 i_418 (.CO (n_676), .S (n_675), .A (n_426), .B (n_428), .CI (n_641));
FA_X1 i_417 (.CO (n_674), .S (n_452), .A (n_448), .B (n_450), .CI (n_441));
FA_X1 i_416 (.CO (n_673), .S (n_450), .A (n_446), .B (n_437), .CI (n_439));
FA_X1 i_415 (.CO (n_672), .S (n_446), .A (p_11[37]), .B (n_433), .CI (n_530));
FA_X1 i_414 (.CO (n_671), .S (n_448), .A (n_435), .B (n_444), .CI (n_526));
FA_X1 i_413 (.CO (n_670), .S (n_444), .A (p_8[37]), .B (p_9[37]), .CI (p_10[37]));
HA_X1 i_412 (.CO (n_443), .S (n_669), .A (n_429), .B (n_440));
FA_X1 i_411 (.CO (n_441), .S (n_440), .A (n_427), .B (n_436), .CI (n_438));
FA_X1 i_410 (.CO (n_439), .S (n_438), .A (n_432), .B (n_529), .CI (n_425));
FA_X1 i_409 (.CO (n_433), .S (n_432), .A (p_7[36]), .B (p_8[36]), .CI (p_9[36]));
FA_X1 i_408 (.CO (n_437), .S (n_436), .A (n_533), .B (n_423), .CI (n_434));
FA_X1 i_407 (.CO (n_435), .S (n_434), .A (p_10[36]), .B (p_11[36]), .CI (n_421));
FA_X1 i_406 (.CO (n_427), .S (n_426), .A (n_422), .B (n_420), .CI (n_531));
FA_X1 i_405 (.CO (n_421), .S (n_420), .A (p_7[35]), .B (p_8[35]), .CI (p_9[35]));
FA_X1 i_404 (.CO (n_423), .S (n_422), .A (p_10[35]), .B (p_11[35]), .CI (n_635));
FA_X1 i_403 (.CO (n_429), .S (n_428), .A (n_424), .B (n_637), .CI (n_640));
FA_X1 i_402 (.CO (n_425), .S (n_424), .A (n_636), .B (n_646), .CI (n_638));
INV_X1 i_401 (.ZN (n_668), .A (n_605));
INV_X1 i_400 (.ZN (n_667), .A (p_5[34]));
INV_X1 i_399 (.ZN (n_666), .A (p_5[33]));
INV_X1 i_398 (.ZN (n_665), .A (p_3[32]));
INV_X1 i_397 (.ZN (n_664), .A (p_4[34]));
INV_X1 i_396 (.ZN (n_663), .A (p_4[33]));
INV_X1 i_395 (.ZN (n_662), .A (p_4[32]));
NAND2_X1 i_394 (.ZN (n_661), .A1 (n_665), .A2 (n_662));
NOR2_X1 i_393 (.ZN (n_660), .A1 (n_631), .A2 (n_634));
AND3_X1 i_392 (.ZN (n_659), .A1 (n_369), .A2 (n_367), .A3 (n_283));
OAI21_X1 i_391 (.ZN (n_658), .A (n_478), .B1 (n_471), .B2 (n_659));
OAI21_X1 i_390 (.ZN (n_657), .A (n_626), .B1 (n_633), .B2 (n_621));
NOR2_X1 i_389 (.ZN (n_656), .A1 (n_660), .A2 (n_657));
OAI21_X1 i_388 (.ZN (n_655), .A (n_656), .B1 (n_592), .B2 (n_537));
INV_X1 i_387 (.ZN (n_654), .A (n_655));
NAND3_X2 i_386 (.ZN (n_653), .A1 (n_668), .A2 (n_658), .A3 (n_654));
NAND2_X1 i_385 (.ZN (n_652), .A1 (n_633), .A2 (n_621));
OAI21_X1 i_384 (.ZN (n_651), .A (n_656), .B1 (n_622), .B2 (n_627));
NAND2_X1 i_383 (.ZN (n_650), .A1 (n_631), .A2 (n_634));
OAI211_X1 i_382 (.ZN (n_649), .A (n_650), .B (n_651), .C1 (n_660), .C2 (n_652));
AOI21_X2 i_381 (.ZN (n_648), .A (n_649), .B1 (n_606), .B2 (n_654));
AND2_X2 i_380 (.ZN (n_647), .A1 (n_653), .A2 (n_648));
NAND2_X1 i_379 (.ZN (n_646), .A1 (n_667), .A2 (n_664));
NAND2_X1 i_378 (.ZN (n_645), .A1 (n_632), .A2 (n_642));
OAI21_X1 i_377 (.ZN (n_644), .A (n_645), .B1 (n_632), .B2 (n_642));
XOR2_X2 i_376 (.Z (\aggregated_res[14] [34] ), .A (n_647), .B (n_644));
XOR2_X1 i_375 (.Z (n_536), .A (n_179), .B (n_666));
OAI21_X1 i_374 (.ZN (n_534), .A (n_646), .B1 (n_667), .B2 (n_664));
OAI222_X1 i_373 (.ZN (n_538), .A1 (p_3[40]), .A2 (n_663), .B1 (n_666), .B2 (p_3[40])
    , .C1 (n_666), .C2 (n_663));
HA_X1 i_372 (.CO (n_643), .S (n_642), .A (n_403), .B (n_416));
FA_X1 i_371 (.CO (n_641), .S (n_416), .A (n_401), .B (n_412), .CI (n_414));
FA_X1 i_370 (.CO (n_640), .S (n_414), .A (n_534), .B (n_410), .CI (n_399));
FA_X1 i_369 (.CO (n_381), .S (n_380), .A (p_11[32]), .B (n_363), .CI (n_615));
FA_X1 i_368 (.CO (n_363), .S (n_639), .A (p_8[31]), .B (p_9[31]), .CI (p_10[31]));
FA_X1 i_367 (.CO (n_638), .S (n_410), .A (n_395), .B (n_393), .CI (n_538));
FA_X1 i_366 (.CO (n_393), .S (n_392), .A (p_6[33]), .B (p_7[33]), .CI (p_8[33]));
FA_X1 i_365 (.CO (n_395), .S (n_394), .A (p_9[33]), .B (p_10[33]), .CI (p_11[33]));
FA_X1 i_364 (.CO (n_637), .S (n_412), .A (n_397), .B (n_408), .CI (n_406));
FA_X1 i_363 (.CO (n_636), .S (n_406), .A (p_6[34]), .B (p_7[34]), .CI (p_8[34]));
FA_X1 i_362 (.CO (n_635), .S (n_408), .A (p_9[34]), .B (p_10[34]), .CI (p_11[34]));
FA_X1 i_361 (.CO (n_377), .S (n_376), .A (p_5[32]), .B (p_6[32]), .CI (p_7[32]));
FA_X1 i_360 (.CO (n_379), .S (n_378), .A (p_8[32]), .B (p_9[32]), .CI (p_10[32]));
HA_X1 i_359 (.CO (n_634), .S (n_633), .A (n_620), .B (n_388));
FA_X1 i_358 (.CO (n_632), .S (n_631), .A (n_400), .B (n_389), .CI (n_402));
FA_X1 i_357 (.CO (n_403), .S (n_402), .A (n_385), .B (n_398), .CI (n_387));
FA_X1 i_356 (.CO (n_399), .S (n_398), .A (n_381), .B (n_394), .CI (n_392));
FA_X1 i_355 (.CO (n_389), .S (n_388), .A (n_384), .B (n_619), .CI (n_386));
FA_X1 i_354 (.CO (n_387), .S (n_386), .A (n_618), .B (n_616), .CI (n_382));
FA_X1 i_353 (.CO (n_385), .S (n_384), .A (n_376), .B (n_198), .CI (n_380));
FA_X1 i_352 (.CO (n_401), .S (n_400), .A (n_536), .B (n_396), .CI (n_383));
FA_X1 i_351 (.CO (n_383), .S (n_382), .A (n_203), .B (n_617), .CI (n_378));
FA_X1 i_350 (.CO (n_397), .S (n_396), .A (n_379), .B (n_377), .CI (n_661));
OAI21_X1 i_349 (.ZN (\aggregated_res[14] [31] ), .A (n_629), .B1 (n_623), .B2 (n_628));
INV_X1 i_348 (.ZN (n_630), .A (n_629));
NAND2_X1 i_347 (.ZN (n_629), .A1 (n_628), .A2 (n_623));
NOR2_X1 i_346 (.ZN (n_628), .A1 (n_627), .A2 (n_625));
AND2_X1 i_345 (.ZN (n_627), .A1 (n_595), .A2 (n_374));
INV_X1 i_344 (.ZN (n_626), .A (n_625));
NOR2_X1 i_343 (.ZN (n_625), .A1 (n_595), .A2 (n_374));
INV_X1 i_342 (.ZN (n_624), .A (n_623));
OAI22_X1 i_341 (.ZN (n_623), .A1 (n_622), .A2 (n_603), .B1 (n_537), .B2 (n_592));
INV_X1 i_340 (.ZN (n_622), .A (n_600));
XOR2_X1 i_339 (.Z (n_541), .A (n_209), .B (n_201));
FA_X1 i_338 (.CO (n_621), .S (n_374), .A (n_590), .B (n_372), .CI (n_591));
FA_X1 i_337 (.CO (n_620), .S (n_372), .A (n_589), .B (n_368), .CI (n_370));
FA_X1 i_336 (.CO (n_619), .S (n_370), .A (n_364), .B (n_586), .CI (n_366));
FA_X1 i_335 (.CO (n_618), .S (n_366), .A (n_601), .B (n_584), .CI (n_639));
FA_X1 i_334 (.CO (n_617), .S (n_364), .A (p_11[31]), .B (n_585), .CI (n_587));
FA_X1 i_333 (.CO (n_616), .S (n_368), .A (n_360), .B (n_541), .CI (n_588));
FA_X1 i_332 (.CO (n_615), .S (n_360), .A (p_5[31]), .B (p_6[31]), .CI (p_7[31]));
INV_X1 i_331 (.ZN (n_614), .A (p_2[30]));
INV_X1 i_330 (.ZN (n_613), .A (p_3[30]));
NAND3_X1 i_329 (.ZN (n_612), .A1 (n_560), .A2 (n_572), .A3 (n_575));
AOI21_X1 i_328 (.ZN (n_609), .A (n_612), .B1 (n_559), .B2 (n_461));
NOR2_X1 i_327 (.ZN (n_608), .A1 (n_576), .A2 (n_569));
AOI211_X2 i_326 (.ZN (n_607), .A (n_608), .B (n_609), .C1 (n_535), .C2 (n_539));
INV_X1 i_325 (.ZN (n_606), .A (n_607));
OR2_X1 i_324 (.ZN (n_605), .A1 (n_555), .A2 (n_612));
OAI21_X1 i_323 (.ZN (n_603), .A (n_607), .B1 (n_463), .B2 (n_605));
NAND2_X1 i_322 (.ZN (n_601), .A1 (n_614), .A2 (n_613));
NAND2_X1 i_321 (.ZN (n_600), .A1 (n_592), .A2 (n_537));
OAI21_X1 i_320 (.ZN (n_599), .A (n_600), .B1 (n_592), .B2 (n_537));
XNOR2_X1 i_319 (.ZN (\aggregated_res[14] [30] ), .A (n_603), .B (n_599));
OAI21_X1 i_318 (.ZN (n_544), .A (n_601), .B1 (n_614), .B2 (n_613));
NOR2_X1 i_317 (.ZN (n_598), .A1 (p_2[29]), .A2 (p_3[29]));
NAND2_X1 i_316 (.ZN (n_597), .A1 (p_2[29]), .A2 (p_3[29]));
AOI21_X1 i_315 (.ZN (n_548), .A (n_598), .B1 (p_1[36]), .B2 (n_597));
HA_X1 i_314 (.CO (n_595), .S (n_592), .A (n_532), .B (n_356));
FA_X1 i_313 (.CO (n_591), .S (n_356), .A (n_350), .B (n_527), .CI (n_354));
FA_X1 i_312 (.CO (n_590), .S (n_354), .A (n_525), .B (n_515), .CI (n_352));
FA_X1 i_311 (.CO (n_589), .S (n_352), .A (n_342), .B (n_544), .CI (n_348));
FA_X1 i_310 (.CO (n_588), .S (n_348), .A (n_507), .B (n_548), .CI (n_512));
FA_X1 i_309 (.CO (n_587), .S (n_342), .A (p_4[30]), .B (p_5[30]), .CI (p_6[30]));
FA_X1 i_308 (.CO (n_586), .S (n_350), .A (n_517), .B (n_346), .CI (n_344));
FA_X1 i_307 (.CO (n_585), .S (n_344), .A (p_7[30]), .B (p_8[30]), .CI (p_9[30]));
FA_X1 i_306 (.CO (n_584), .S (n_346), .A (p_10[30]), .B (p_11[30]), .CI (n_522));
INV_X1 i_305 (.ZN (n_583), .A (p_2[28]));
INV_X1 i_304 (.ZN (n_579), .A (p_2[27]));
INV_X1 i_303 (.ZN (n_578), .A (p_1[28]));
INV_X1 i_302 (.ZN (n_577), .A (p_1[27]));
NOR2_X1 i_301 (.ZN (n_576), .A1 (n_535), .A2 (n_539));
INV_X1 i_300 (.ZN (n_575), .A (n_576));
NOR2_X1 i_299 (.ZN (n_574), .A1 (n_322), .A2 (n_303));
INV_X1 i_298 (.ZN (n_572), .A (n_574));
NAND2_X1 i_297 (.ZN (n_569), .A1 (n_322), .A2 (n_303));
INV_X1 i_296 (.ZN (n_568), .A (n_569));
NOR2_X2 i_295 (.ZN (n_565), .A1 (n_451), .A2 (n_302));
INV_X1 i_294 (.ZN (n_560), .A (n_565));
NAND2_X1 i_293 (.ZN (n_559), .A1 (n_451), .A2 (n_302));
INV_X1 i_292 (.ZN (n_557), .A (n_559));
NOR2_X1 i_291 (.ZN (n_555), .A1 (n_411), .A2 (n_449));
AOI21_X1 i_289 (.ZN (n_552), .A (n_555), .B1 (n_461), .B2 (n_463));
OAI21_X1 i_288 (.ZN (n_547), .A (n_560), .B1 (n_557), .B2 (n_552));
INV_X1 i_287 (.ZN (n_545), .A (n_547));
AOI21_X1 i_286 (.ZN (n_543), .A (n_576), .B1 (n_535), .B2 (n_539));
AOI21_X1 i_285 (.ZN (n_542), .A (n_574), .B1 (n_569), .B2 (n_547));
XOR2_X2 i_284 (.Z (\aggregated_res[14] [29] ), .A (n_543), .B (n_542));
OAI222_X1 i_283 (.ZN (n_553), .A1 (n_577), .A2 (p_0[34]), .B1 (n_579), .B2 (p_0[34])
    , .C1 (n_579), .C2 (n_577));
NAND2_X1 i_282 (.ZN (n_550), .A1 (n_583), .A2 (n_578));
OAI21_X1 i_281 (.ZN (n_549), .A (n_550), .B1 (n_583), .B2 (n_578));
XOR2_X1 i_280 (.Z (n_540), .A (p_2[29]), .B (p_1[36]));
XNOR2_X1 i_279 (.ZN (n_546), .A (p_3[29]), .B (n_540));
XOR2_X1 i_278 (.Z (n_551), .A (p_2[27]), .B (n_211));
FA_X1 i_277 (.CO (n_303), .S (n_302), .A (n_298), .B (n_300), .CI (n_447));
HA_X1 i_276 (.CO (n_539), .S (n_322), .A (n_301), .B (n_320));
FA_X1 i_275 (.CO (n_301), .S (n_300), .A (n_294), .B (n_296), .CI (n_445));
FA_X1 i_274 (.CO (n_537), .S (n_535), .A (n_319), .B (n_338), .CI (n_321));
FA_X1 i_273 (.CO (n_321), .S (n_320), .A (n_299), .B (n_316), .CI (n_318));
FA_X1 i_272 (.CO (n_299), .S (n_298), .A (n_292), .B (n_415), .CI (n_419));
FA_X1 i_271 (.CO (n_532), .S (n_338), .A (n_334), .B (n_332), .CI (n_336));
FA_X1 i_270 (.CO (n_527), .S (n_336), .A (n_315), .B (n_313), .CI (n_317));
FA_X1 i_269 (.CO (n_317), .S (n_316), .A (n_310), .B (n_295), .CI (n_293));
FA_X1 i_268 (.CO (n_293), .S (n_292), .A (n_462), .B (n_413), .CI (n_288));
FA_X1 i_267 (.CO (n_295), .S (n_294), .A (n_286), .B (n_284), .CI (n_551));
FA_X1 i_266 (.CO (n_525), .S (n_332), .A (n_311), .B (n_328), .CI (n_326));
FA_X1 i_265 (.CO (n_522), .S (n_326), .A (p_7[29]), .B (p_8[29]), .CI (p_9[29]));
FA_X1 i_264 (.CO (n_517), .S (n_328), .A (p_10[29]), .B (p_11[29]), .CI (n_309));
FA_X1 i_263 (.CO (n_311), .S (n_310), .A (n_289), .B (n_287), .CI (n_285));
FA_X1 i_262 (.CO (n_285), .S (n_284), .A (p_3[27]), .B (p_4[27]), .CI (p_5[27]));
FA_X1 i_261 (.CO (n_287), .S (n_286), .A (p_6[27]), .B (p_7[27]), .CI (p_8[27]));
FA_X1 i_260 (.CO (n_289), .S (n_288), .A (p_9[27]), .B (p_10[27]), .CI (p_11[27]));
FA_X1 i_259 (.CO (n_515), .S (n_334), .A (n_324), .B (n_546), .CI (n_330));
FA_X1 i_258 (.CO (n_512), .S (n_330), .A (n_307), .B (n_305), .CI (n_550));
FA_X1 i_257 (.CO (n_507), .S (n_324), .A (p_4[29]), .B (p_5[29]), .CI (p_6[29]));
FA_X1 i_256 (.CO (n_319), .S (n_318), .A (n_312), .B (n_297), .CI (n_314));
FA_X1 i_255 (.CO (n_315), .S (n_314), .A (n_306), .B (n_304), .CI (n_549));
FA_X1 i_254 (.CO (n_305), .S (n_304), .A (p_3[28]), .B (p_4[28]), .CI (p_5[28]));
FA_X1 i_253 (.CO (n_307), .S (n_306), .A (p_6[28]), .B (p_7[28]), .CI (p_8[28]));
FA_X1 i_252 (.CO (n_297), .S (n_296), .A (n_418), .B (n_290), .CI (n_442));
FA_X1 i_251 (.CO (n_313), .S (n_312), .A (n_553), .B (n_291), .CI (n_308));
FA_X1 i_250 (.CO (n_309), .S (n_308), .A (p_9[28]), .B (p_10[28]), .CI (p_11[28]));
FA_X1 i_249 (.CO (n_291), .S (n_290), .A (n_430), .B (n_431), .CI (n_417));
INV_X1 i_248 (.ZN (n_505), .A (p_0[26]));
INV_X1 i_247 (.ZN (n_503), .A (p_0[25]));
INV_X1 i_246 (.ZN (n_502), .A (p_1[26]));
INV_X1 i_245 (.ZN (n_501), .A (p_1[25]));
INV_X1 i_244 (.ZN (n_500), .A (p_11[25]));
INV_X1 i_243 (.ZN (n_499), .A (n_282));
INV_X1 i_242 (.ZN (n_494), .A (n_227));
AOI21_X1 i_241 (.ZN (n_491), .A (n_275), .B1 (n_213), .B2 (n_215));
INV_X1 i_240 (.ZN (n_490), .A (n_491));
NOR2_X1 i_239 (.ZN (n_489), .A1 (n_405), .A2 (n_269));
NOR2_X2 i_238 (.ZN (n_487), .A1 (n_407), .A2 (n_409));
NAND2_X1 i_237 (.ZN (n_485), .A1 (n_405), .A2 (n_269));
NOR3_X2 i_236 (.ZN (n_483), .A1 (n_277), .A2 (n_487), .A3 (n_489));
NOR2_X1 i_235 (.ZN (n_481), .A1 (n_487), .A2 (n_485));
AOI221_X1 i_234 (.ZN (n_478), .A (n_481), .B1 (n_407), .B2 (n_409), .C1 (n_490), .C2 (n_483));
OAI21_X1 i_233 (.ZN (n_471), .A (n_483), .B1 (n_213), .B2 (n_215));
OAI21_X1 i_232 (.ZN (n_470), .A (n_478), .B1 (n_499), .B2 (n_471));
INV_X1 i_231 (.ZN (n_463), .A (n_470));
NAND2_X1 i_230 (.ZN (n_462), .A1 (n_505), .A2 (n_502));
NAND2_X1 i_229 (.ZN (n_461), .A1 (n_411), .A2 (n_449));
OAI21_X1 i_228 (.ZN (n_459), .A (n_461), .B1 (n_411), .B2 (n_449));
XNOR2_X1 i_227 (.ZN (\aggregated_res[14] [26] ), .A (n_470), .B (n_459));
NAND2_X1 i_226 (.ZN (n_562), .A1 (n_503), .A2 (n_501));
OAI21_X1 i_225 (.ZN (n_561), .A (n_562), .B1 (n_503), .B2 (n_501));
NAND2_X1 i_224 (.ZN (n_457), .A1 (p_15[32]), .A2 (n_494));
INV_X1 i_223 (.ZN (n_455), .A (n_457));
OAI21_X1 i_222 (.ZN (n_453), .A (n_457), .B1 (p_15[32]), .B2 (n_494));
OAI22_X1 i_221 (.ZN (n_556), .A1 (p_15[32]), .A2 (n_494), .B1 (n_500), .B2 (n_455));
XNOR2_X1 i_220 (.ZN (n_558), .A (p_11[25]), .B (n_453));
OAI21_X1 i_219 (.ZN (n_554), .A (n_462), .B1 (n_505), .B2 (n_502));
HA_X1 i_218 (.CO (n_451), .S (n_449), .A (n_259), .B (n_280));
FA_X1 i_217 (.CO (n_447), .S (n_280), .A (n_276), .B (n_257), .CI (n_278));
FA_X1 i_216 (.CO (n_445), .S (n_278), .A (n_255), .B (n_274), .CI (n_272));
FA_X1 i_215 (.CO (n_442), .S (n_272), .A (n_556), .B (n_266), .CI (n_264));
FA_X1 i_214 (.CO (n_431), .S (n_264), .A (p_5[26]), .B (p_6[26]), .CI (p_7[26]));
FA_X1 i_213 (.CO (n_430), .S (n_266), .A (p_8[26]), .B (p_9[26]), .CI (p_10[26]));
FA_X1 i_212 (.CO (n_419), .S (n_274), .A (n_262), .B (n_554), .CI (n_270));
FA_X1 i_211 (.CO (n_418), .S (n_270), .A (n_243), .B (n_562), .CI (n_249));
FA_X1 i_210 (.CO (n_417), .S (n_262), .A (p_2[26]), .B (p_3[26]), .CI (p_4[26]));
FA_X1 i_209 (.CO (n_415), .S (n_276), .A (n_268), .B (n_253), .CI (n_251));
FA_X1 i_208 (.CO (n_413), .S (n_268), .A (p_11[26]), .B (n_247), .CI (n_245));
HA_X1 i_207 (.CO (n_411), .S (n_409), .A (n_256), .B (n_258));
FA_X1 i_206 (.CO (n_259), .S (n_258), .A (n_237), .B (n_254), .CI (n_239));
FA_X1 i_205 (.CO (n_255), .S (n_254), .A (n_231), .B (n_248), .CI (n_233));
FA_X1 i_204 (.CO (n_227), .S (n_226), .A (p_9[24]), .B (p_10[24]), .CI (p_11[24]));
FA_X1 i_203 (.CO (n_249), .S (n_248), .A (n_225), .B (n_223), .CI (n_221));
FA_X1 i_202 (.CO (n_223), .S (n_222), .A (p_3[24]), .B (p_4[24]), .CI (p_5[24]));
FA_X1 i_201 (.CO (n_225), .S (n_224), .A (p_6[24]), .B (p_7[24]), .CI (p_8[24]));
FA_X1 i_200 (.CO (n_257), .S (n_256), .A (n_235), .B (n_252), .CI (n_250));
FA_X1 i_199 (.CO (n_251), .S (n_250), .A (n_229), .B (n_558), .CI (n_246));
FA_X1 i_198 (.CO (n_247), .S (n_246), .A (p_8[25]), .B (p_9[25]), .CI (p_10[25]));
FA_X1 i_197 (.CO (n_253), .S (n_252), .A (n_244), .B (n_242), .CI (n_561));
FA_X1 i_196 (.CO (n_243), .S (n_242), .A (p_2[25]), .B (p_3[25]), .CI (p_4[25]));
FA_X1 i_195 (.CO (n_245), .S (n_244), .A (p_5[25]), .B (p_6[25]), .CI (p_7[25]));
FA_X1 i_194 (.CO (n_229), .S (n_228), .A (p_15[24]), .B (n_240), .CI (n_260));
FA_X1 i_193 (.CO (n_231), .S (n_230), .A (n_261), .B (n_263), .CI (n_217));
FA_X1 i_192 (.CO (n_221), .S (n_220), .A (p_0[24]), .B (p_1[24]), .CI (p_2[24]));
HA_X1 i_191 (.CO (n_407), .S (n_405), .A (n_267), .B (n_238));
FA_X1 i_190 (.CO (n_239), .S (n_238), .A (n_232), .B (n_236), .CI (n_234));
FA_X1 i_189 (.CO (n_235), .S (n_234), .A (n_220), .B (n_230), .CI (n_228));
FA_X1 i_188 (.CO (n_237), .S (n_236), .A (n_265), .B (n_241), .CI (n_219));
FA_X1 i_187 (.CO (n_233), .S (n_232), .A (n_226), .B (n_224), .CI (n_222));
INV_X1 i_186 (.ZN (n_404), .A (n_143));
OAI222_X1 i_185 (.ZN (n_391), .A1 (n_143), .A2 (n_160), .B1 (n_161), .B2 (n_178), .C1 (n_142), .C2 (n_127));
INV_X1 i_184 (.ZN (n_390), .A (n_391));
AOI22_X1 i_183 (.ZN (n_375), .A1 (n_126), .A2 (n_111), .B1 (n_142), .B2 (n_127));
OAI21_X1 i_182 (.ZN (n_373), .A (n_160), .B1 (n_161), .B2 (n_178));
OAI22_X1 i_181 (.ZN (n_371), .A1 (n_391), .A2 (n_375), .B1 (n_404), .B2 (n_373));
INV_X1 i_180 (.ZN (n_369), .A (n_371));
NAND2_X1 i_179 (.ZN (n_367), .A1 (n_161), .A2 (n_178));
NOR2_X1 i_178 (.ZN (n_365), .A1 (n_46), .A2 (n_48));
NOR2_X1 i_177 (.ZN (n_362), .A1 (n_58), .A2 (n_49));
OAI22_X1 i_176 (.ZN (n_361), .A1 (n_58), .A2 (n_49), .B1 (n_38), .B2 (n_31));
AOI22_X1 i_175 (.ZN (n_359), .A1 (n_30), .A2 (n_28), .B1 (n_38), .B2 (n_31));
OAI222_X1 i_174 (.ZN (n_358), .A1 (p_0[3]), .A2 (p_15[3]), .B1 (p_15[4]), .B2 (n_0)
    , .C1 (n_207), .C2 (n_205));
INV_X1 i_173 (.ZN (n_357), .A (n_358));
AOI221_X1 i_172 (.ZN (n_355), .A (n_357), .B1 (p_15[4]), .B2 (n_0), .C1 (n_2), .C2 (n_1));
NOR2_X1 i_171 (.ZN (n_353), .A1 (n_22), .A2 (n_17));
OAI222_X1 i_170 (.ZN (n_351), .A1 (n_10), .A2 (n_8), .B1 (n_12), .B2 (n_16), .C1 (n_22), .C2 (n_17));
INV_X1 i_169 (.ZN (n_349), .A (n_351));
OAI221_X1 i_168 (.ZN (n_347), .A (n_349), .B1 (n_4), .B2 (n_6), .C1 (n_2), .C2 (n_1));
AOI22_X1 i_167 (.ZN (n_345), .A1 (n_4), .A2 (n_6), .B1 (n_10), .B2 (n_8));
AOI22_X1 i_166 (.ZN (n_343), .A1 (n_12), .A2 (n_16), .B1 (n_22), .B2 (n_17));
OAI222_X1 i_165 (.ZN (n_341), .A1 (n_351), .A2 (n_345), .B1 (n_353), .B2 (n_343), .C1 (n_355), .C2 (n_347));
OAI21_X1 i_164 (.ZN (n_340), .A (n_341), .B1 (n_30), .B2 (n_28));
AOI211_X2 i_163 (.ZN (n_339), .A (n_365), .B (n_361), .C1 (n_359), .C2 (n_340));
AOI22_X1 i_162 (.ZN (n_337), .A1 (n_58), .A2 (n_49), .B1 (n_46), .B2 (n_48));
NOR2_X1 i_161 (.ZN (n_335), .A1 (n_362), .A2 (n_337));
NOR2_X1 i_160 (.ZN (n_333), .A1 (n_110), .A2 (n_97));
OAI222_X1 i_159 (.ZN (n_331), .A1 (n_83), .A2 (n_96), .B1 (n_110), .B2 (n_97), .C1 (n_82), .C2 (n_71));
OAI22_X1 i_158 (.ZN (n_329), .A1 (n_339), .A2 (n_335), .B1 (n_70), .B2 (n_59));
AOI22_X1 i_157 (.ZN (n_327), .A1 (n_70), .A2 (n_59), .B1 (n_82), .B2 (n_71));
AOI22_X1 i_156 (.ZN (n_325), .A1 (n_110), .A2 (n_97), .B1 (n_83), .B2 (n_96));
OAI222_X2 i_155 (.ZN (n_323), .A1 (n_331), .A2 (n_327), .B1 (n_333), .B2 (n_325), .C1 (n_331), .C2 (n_329));
OAI211_X1 i_154 (.ZN (n_283), .A (n_323), .B (n_390), .C1 (n_126), .C2 (n_111));
NAND3_X1 i_153 (.ZN (n_282), .A1 (n_369), .A2 (n_367), .A3 (n_283));
OAI21_X1 i_152 (.ZN (n_281), .A (n_282), .B1 (n_213), .B2 (n_215));
INV_X1 i_151 (.ZN (n_279), .A (n_281));
NOR2_X1 i_150 (.ZN (n_277), .A1 (n_199), .A2 (n_218));
AND2_X1 i_149 (.ZN (n_275), .A1 (n_199), .A2 (n_218));
AOI21_X1 i_148 (.ZN (n_273), .A (n_279), .B1 (n_213), .B2 (n_215));
NOR2_X1 i_147 (.ZN (n_271), .A1 (n_277), .A2 (n_275));
XNOR2_X1 i_146 (.ZN (\aggregated_res[14] [23] ), .A (n_273), .B (n_271));
FA_X1 i_145 (.CO (n_269), .S (n_218), .A (n_214), .B (n_197), .CI (n_216));
FA_X1 i_144 (.CO (n_267), .S (n_216), .A (n_210), .B (n_212), .CI (n_195));
FA_X1 i_143 (.CO (n_265), .S (n_212), .A (n_204), .B (n_202), .CI (n_200));
FA_X1 i_142 (.CO (n_263), .S (n_200), .A (p_0[23]), .B (p_1[23]), .CI (p_2[23]));
FA_X1 i_141 (.CO (n_261), .S (n_202), .A (p_3[23]), .B (p_4[23]), .CI (p_5[23]));
FA_X1 i_140 (.CO (n_260), .S (n_204), .A (p_6[23]), .B (p_7[23]), .CI (p_8[23]));
FA_X1 i_139 (.CO (n_241), .S (n_210), .A (n_181), .B (n_189), .CI (n_206));
FA_X1 i_138 (.CO (n_240), .S (n_206), .A (p_9[23]), .B (p_10[23]), .CI (p_15[23]));
FA_X1 i_137 (.CO (n_219), .S (n_214), .A (n_208), .B (n_191), .CI (n_193));
FA_X1 i_136 (.CO (n_217), .S (n_208), .A (n_187), .B (n_185), .CI (n_183));
HA_X1 i_135 (.CO (n_199), .S (n_215), .A (n_177), .B (n_196));
FA_X1 i_134 (.CO (n_197), .S (n_196), .A (n_192), .B (n_190), .CI (n_194));
FA_X1 i_133 (.CO (n_195), .S (n_194), .A (n_188), .B (n_173), .CI (n_175));
FA_X1 i_132 (.CO (n_189), .S (n_188), .A (n_167), .B (n_165), .CI (n_163));
FA_X1 i_131 (.CO (n_165), .S (n_164), .A (p_3[21]), .B (p_4[21]), .CI (p_5[21]));
FA_X1 i_130 (.CO (n_167), .S (n_166), .A (p_6[21]), .B (p_7[21]), .CI (p_8[21]));
FA_X1 i_129 (.CO (n_191), .S (n_190), .A (n_169), .B (n_186), .CI (n_184));
FA_X1 i_128 (.CO (n_185), .S (n_184), .A (p_6[22]), .B (p_7[22]), .CI (p_8[22]));
FA_X1 i_127 (.CO (n_187), .S (n_186), .A (p_9[22]), .B (p_10[22]), .CI (p_15[22]));
FA_X1 i_126 (.CO (n_169), .S (n_168), .A (p_9[21]), .B (p_15[21]), .CI (n_149));
FA_X1 i_125 (.CO (n_149), .S (n_148), .A (p_6[20]), .B (p_7[20]), .CI (p_8[20]));
FA_X1 i_124 (.CO (n_193), .S (n_192), .A (n_182), .B (n_180), .CI (n_171));
FA_X1 i_123 (.CO (n_151), .S (n_150), .A (p_9[20]), .B (p_15[20]), .CI (n_133));
FA_X1 i_122 (.CO (n_133), .S (n_132), .A (p_6[19]), .B (p_7[19]), .CI (p_8[19]));
FA_X1 i_121 (.CO (n_147), .S (n_146), .A (p_3[20]), .B (p_4[20]), .CI (p_5[20]));
FA_X1 i_120 (.CO (n_181), .S (n_180), .A (p_0[22]), .B (p_1[22]), .CI (p_2[22]));
FA_X1 i_119 (.CO (n_183), .S (n_182), .A (p_3[22]), .B (p_4[22]), .CI (p_5[22]));
HA_X1 i_118 (.CO (n_1), .S (n_0), .A (p_0[4]), .B (p_1[4]));
FA_X1 i_117 (.CO (n_3), .S (n_2), .A (p_0[5]), .B (p_1[5]), .CI (p_15[5]));
HA_X1 i_116 (.CO (n_7), .S (n_6), .A (p_15[6]), .B (n_3));
FA_X1 i_115 (.CO (n_5), .S (n_4), .A (p_0[6]), .B (p_1[6]), .CI (p_2[6]));
FA_X1 i_114 (.CO (n_9), .S (n_8), .A (p_0[7]), .B (p_1[7]), .CI (p_2[7]));
HA_X1 i_113 (.CO (n_17), .S (n_16), .A (n_11), .B (n_14));
FA_X1 i_112 (.CO (n_15), .S (n_14), .A (p_3[8]), .B (p_15[8]), .CI (n_9));
FA_X1 i_111 (.CO (n_11), .S (n_10), .A (p_15[7]), .B (n_5), .CI (n_7));
FA_X1 i_110 (.CO (n_13), .S (n_12), .A (p_0[8]), .B (p_1[8]), .CI (p_2[8]));
FA_X1 i_109 (.CO (n_27), .S (n_26), .A (p_3[10]), .B (p_4[10]), .CI (p_15[10]));
FA_X1 i_108 (.CO (n_21), .S (n_20), .A (p_3[9]), .B (p_15[9]), .CI (n_13));
FA_X1 i_107 (.CO (n_19), .S (n_18), .A (p_0[9]), .B (p_1[9]), .CI (p_2[9]));
FA_X1 i_106 (.CO (n_29), .S (n_28), .A (n_19), .B (n_21), .CI (n_26));
HA_X1 i_105 (.CO (n_31), .S (n_30), .A (n_24), .B (n_23));
FA_X1 i_104 (.CO (n_23), .S (n_22), .A (n_15), .B (n_20), .CI (n_18));
FA_X1 i_103 (.CO (n_25), .S (n_24), .A (p_0[10]), .B (p_1[10]), .CI (p_2[10]));
HA_X1 i_102 (.CO (n_49), .S (n_48), .A (n_37), .B (n_39));
FA_X1 i_101 (.CO (n_39), .S (n_38), .A (n_32), .B (n_29), .CI (n_36));
FA_X1 i_100 (.CO (n_37), .S (n_36), .A (n_27), .B (n_25), .CI (n_34));
FA_X1 i_99 (.CO (n_59), .S (n_58), .A (n_54), .B (n_47), .CI (n_56));
FA_X1 i_98 (.CO (n_47), .S (n_46), .A (n_42), .B (n_40), .CI (n_44));
FA_X1 i_97 (.CO (n_33), .S (n_32), .A (p_0[11]), .B (p_1[11]), .CI (p_2[11]));
FA_X1 i_96 (.CO (n_35), .S (n_34), .A (p_3[11]), .B (p_4[11]), .CI (p_15[11]));
FA_X1 i_95 (.CO (n_41), .S (n_40), .A (p_0[12]), .B (p_1[12]), .CI (p_2[12]));
FA_X1 i_94 (.CO (n_43), .S (n_42), .A (p_3[12]), .B (p_4[12]), .CI (p_5[12]));
HA_X1 i_93 (.CO (n_71), .S (n_70), .A (n_66), .B (n_68));
HA_X1 i_92 (.CO (n_97), .S (n_96), .A (n_92), .B (n_94));
FA_X1 i_91 (.CO (n_85), .S (n_84), .A (p_0[16]), .B (p_1[16]), .CI (p_2[16]));
FA_X1 i_90 (.CO (n_87), .S (n_86), .A (p_3[16]), .B (p_4[16]), .CI (p_5[16]));
FA_X1 i_89 (.CO (n_89), .S (n_88), .A (p_6[16]), .B (p_7[16]), .CI (p_15[16]));
FA_X1 i_88 (.CO (n_83), .S (n_82), .A (n_78), .B (n_69), .CI (n_80));
FA_X1 i_87 (.CO (n_67), .S (n_66), .A (n_51), .B (n_55), .CI (n_64));
FA_X1 i_86 (.CO (n_55), .S (n_54), .A (p_15[13]), .B (n_43), .CI (n_41));
FA_X1 i_85 (.CO (n_73), .S (n_72), .A (p_0[15]), .B (p_1[15]), .CI (p_2[15]));
FA_X1 i_84 (.CO (n_75), .S (n_74), .A (p_3[15]), .B (p_4[15]), .CI (p_5[15]));
FA_X1 i_83 (.CO (n_69), .S (n_68), .A (n_62), .B (n_60), .CI (n_57));
FA_X1 i_82 (.CO (n_57), .S (n_56), .A (n_45), .B (n_52), .CI (n_50));
FA_X1 i_81 (.CO (n_51), .S (n_50), .A (p_0[13]), .B (p_1[13]), .CI (p_2[13]));
FA_X1 i_80 (.CO (n_45), .S (n_44), .A (p_15[12]), .B (n_35), .CI (n_33));
FA_X1 i_79 (.CO (n_77), .S (n_76), .A (p_6[15]), .B (p_15[15]), .CI (n_63));
FA_X1 i_78 (.CO (n_63), .S (n_62), .A (p_3[14]), .B (p_4[14]), .CI (p_5[14]));
FA_X1 i_77 (.CO (n_65), .S (n_64), .A (p_6[14]), .B (p_15[14]), .CI (n_53));
FA_X1 i_76 (.CO (n_53), .S (n_52), .A (p_3[13]), .B (p_4[13]), .CI (p_5[13]));
FA_X1 i_75 (.CO (n_61), .S (n_60), .A (p_0[14]), .B (p_1[14]), .CI (p_2[14]));
FA_X1 i_74 (.CO (n_111), .S (n_110), .A (n_106), .B (n_95), .CI (n_108));
FA_X1 i_73 (.CO (n_93), .S (n_92), .A (n_88), .B (n_86), .CI (n_84));
FA_X1 i_72 (.CO (n_105), .S (n_104), .A (n_89), .B (n_87), .CI (n_85));
FA_X1 i_71 (.CO (n_95), .S (n_94), .A (n_90), .B (n_79), .CI (n_81));
FA_X1 i_70 (.CO (n_81), .S (n_80), .A (n_74), .B (n_72), .CI (n_67));
FA_X1 i_69 (.CO (n_79), .S (n_78), .A (n_61), .B (n_65), .CI (n_76));
FA_X1 i_68 (.CO (n_91), .S (n_90), .A (n_75), .B (n_73), .CI (n_77));
FA_X1 i_67 (.CO (n_99), .S (n_98), .A (p_0[17]), .B (p_1[17]), .CI (p_2[17]));
FA_X1 i_66 (.CO (n_101), .S (n_100), .A (p_3[17]), .B (p_4[17]), .CI (p_5[17]));
FA_X1 i_65 (.CO (n_103), .S (n_102), .A (p_6[17]), .B (p_7[17]), .CI (p_15[17]));
HA_X1 i_64 (.CO (n_127), .S (n_126), .A (n_122), .B (n_124));
FA_X1 i_63 (.CO (n_119), .S (n_118), .A (p_15[18]), .B (n_103), .CI (n_101));
FA_X1 i_62 (.CO (n_113), .S (n_112), .A (p_0[18]), .B (p_1[18]), .CI (p_2[18]));
FA_X1 i_61 (.CO (n_115), .S (n_114), .A (p_3[18]), .B (p_4[18]), .CI (p_5[18]));
FA_X1 i_60 (.CO (n_213), .S (n_178), .A (n_174), .B (n_159), .CI (n_176));
FA_X1 i_59 (.CO (n_177), .S (n_176), .A (n_155), .B (n_157), .CI (n_172));
FA_X1 i_57 (.CO (n_173), .S (n_172), .A (n_168), .B (n_166), .CI (n_164));
FA_X1 i_56 (.CO (n_175), .S (n_174), .A (n_162), .B (n_153), .CI (n_170));
FA_X1 i_55 (.CO (n_171), .S (n_170), .A (n_147), .B (n_145), .CI (n_151));
FA_X1 i_54 (.CO (n_163), .S (n_162), .A (p_0[21]), .B (p_1[21]), .CI (p_2[21]));
HA_X1 i_53 (.CO (n_161), .S (n_160), .A (n_156), .B (n_158));
FA_X1 i_52 (.CO (n_159), .S (n_158), .A (n_139), .B (n_154), .CI (n_141));
FA_X1 i_51 (.CO (n_155), .S (n_154), .A (n_150), .B (n_148), .CI (n_146));
FA_X1 i_50 (.CO (n_157), .S (n_156), .A (n_144), .B (n_152), .CI (n_137));
FA_X1 i_49 (.CO (n_153), .S (n_152), .A (n_131), .B (n_129), .CI (n_135));
FA_X1 i_48 (.CO (n_145), .S (n_144), .A (p_0[20]), .B (p_1[20]), .CI (p_2[20]));
FA_X1 i_47 (.CO (n_143), .S (n_142), .A (n_138), .B (n_125), .CI (n_140));
FA_X1 i_46 (.CO (n_141), .S (n_140), .A (n_121), .B (n_136), .CI (n_123));
FA_X1 i_45 (.CO (n_123), .S (n_122), .A (n_114), .B (n_112), .CI (n_118));
FA_X1 i_44 (.CO (n_137), .S (n_136), .A (n_113), .B (n_119), .CI (n_132));
FA_X1 i_43 (.CO (n_125), .S (n_124), .A (n_107), .B (n_120), .CI (n_109));
FA_X1 i_42 (.CO (n_109), .S (n_108), .A (n_91), .B (n_104), .CI (n_93));
FA_X1 i_41 (.CO (n_121), .S (n_120), .A (n_99), .B (n_105), .CI (n_116));
FA_X1 i_40 (.CO (n_107), .S (n_106), .A (n_102), .B (n_100), .CI (n_98));
FA_X1 i_39 (.CO (n_139), .S (n_138), .A (n_130), .B (n_128), .CI (n_134));
FA_X1 i_38 (.CO (n_135), .S (n_134), .A (p_15[19]), .B (n_117), .CI (n_115));
FA_X1 i_37 (.CO (n_129), .S (n_128), .A (p_0[19]), .B (p_1[19]), .CI (p_2[19]));
FA_X1 i_36 (.CO (n_131), .S (n_130), .A (p_3[19]), .B (p_4[19]), .CI (p_5[19]));
XNOR2_X1 i_35 (.ZN (n_211), .A (p_1[27]), .B (p_0[34]));
OAI21_X1 i_34 (.ZN (n_739), .A (n_626), .B1 (n_621), .B2 (n_633));
INV_X1 i_33 (.ZN (n_786), .A (p_3[31]));
INV_X1 i_32 (.ZN (n_209), .A (p_4[31]));
AND2_X1 i_456 (.ZN (n_207), .A1 (p_0[2]), .A2 (p_15[2]));
AND2_X1 i_455 (.ZN (n_205), .A1 (p_0[3]), .A2 (p_15[3]));
NOR2_X1 i_31 (.ZN (n_611), .A1 (n_774), .A2 (n_779));
OAI22_X1 i_30 (.ZN (n_610), .A1 (n_749), .A2 (n_765), .B1 (n_777), .B2 (n_781));
XNOR2_X1 i_29 (.ZN (\aggregated_res[14] [44] ), .A (n_611), .B (n_610));
XOR2_X1 i_28 (.Z (\aggregated_res[14] [43] ), .A (n_781), .B (n_775));
AOI21_X1 i_27 (.ZN (n_604), .A (n_736), .B1 (n_703), .B2 (n_722));
NOR2_X1 i_26 (.ZN (n_602), .A1 (n_754), .A2 (n_737));
XOR2_X1 i_25 (.Z (\aggregated_res[14] [40] ), .A (n_731), .B (n_602));
XOR2_X1 i_24 (.Z (\aggregated_res[14] [39] ), .A (n_732), .B (n_604));
AOI21_X1 i_23 (.ZN (n_596), .A (n_689), .B1 (n_643), .B2 (n_675));
NOR2_X1 i_22 (.ZN (n_594), .A1 (n_708), .A2 (n_690));
XOR2_X1 i_21 (.Z (\aggregated_res[14] [36] ), .A (n_684), .B (n_594));
XOR2_X1 i_20 (.Z (\aggregated_res[14] [35] ), .A (n_685), .B (n_596));
AOI21_X1 i_19 (.ZN (n_593), .A (n_660), .B1 (n_634), .B2 (n_631));
OAI21_X1 i_18 (.ZN (n_582), .A (n_652), .B1 (n_739), .B2 (n_630));
XOR2_X2 i_17 (.Z (\aggregated_res[14] [33] ), .A (n_593), .B (n_582));
OAI21_X1 i_16 (.ZN (n_581), .A (n_652), .B1 (n_621), .B2 (n_633));
OAI21_X1 i_15 (.ZN (n_580), .A (n_626), .B1 (n_627), .B2 (n_624));
XOR2_X1 i_14 (.Z (\aggregated_res[14] [32] ), .A (n_581), .B (n_580));
NOR2_X1 i_13 (.ZN (n_573), .A1 (n_565), .A2 (n_557));
NOR2_X1 i_12 (.ZN (n_571), .A1 (n_574), .A2 (n_568));
XOR2_X2 i_11 (.Z (\aggregated_res[14] [28] ), .A (n_545), .B (n_571));
XOR2_X2 i_10 (.Z (\aggregated_res[14] [27] ), .A (n_552), .B (n_573));
AOI21_X1 i_9 (.ZN (n_570), .A (n_487), .B1 (n_407), .B2 (n_409));
AOI21_X1 i_8 (.ZN (n_567), .A (n_277), .B1 (n_491), .B2 (n_281));
INV_X1 i_7 (.ZN (n_566), .A (n_567));
AOI21_X1 i_6 (.ZN (n_564), .A (n_489), .B1 (n_485), .B2 (n_566));
XOR2_X1 i_5 (.Z (\aggregated_res[14] [25] ), .A (n_570), .B (n_564));
AOI21_X1 i_4 (.ZN (n_563), .A (n_489), .B1 (n_269), .B2 (n_405));
XOR2_X1 i_3 (.Z (\aggregated_res[14] [24] ), .A (n_567), .B (n_563));
OAI222_X1 i_2 (.ZN (n_203), .A1 (p_2[38]), .A2 (n_209), .B1 (p_2[38]), .B2 (n_786)
    , .C1 (n_786), .C2 (n_209));
XOR2_X1 i_290 (.Z (n_201), .A (p_2[38]), .B (p_3[31]));
OAI21_X1 i_1 (.ZN (n_198), .A (n_661), .B1 (n_665), .B2 (n_662));
XOR2_X1 i_0 (.Z (n_179), .A (p_3[40]), .B (p_4[33]));
FA_X1 i_58 (.CO (n_117), .S (n_116), .A (p_6[18]), .B (p_7[18]), .CI (p_8[18]));

endmodule //datapath__0_67

module datapath__0_0 (A_imm, A_imm_2s_complement);

output [31:0] A_imm_2s_complement;
input [31:0] A_imm;
wire n_43;
wire n_38;
wire n_5;
wire n_45;
wire n_3;
wire n_4;
wire n_1;
wire n_2;
wire n_40;
wire n_0;
wire n_50;
wire n_9;
wire n_10;
wire n_7;
wire n_8;
wire n_37;
wire n_6;
wire n_47;
wire n_56;
wire n_46;
wire n_17;
wire n_36;
wire n_15;
wire n_16;
wire n_13;
wire n_14;
wire n_34;
wire n_12;
wire n_54;
wire n_23;
wire n_33;
wire n_21;
wire n_22;
wire n_19;
wire n_20;
wire n_31;
wire n_18;
wire n_52;
wire n_25;
wire n_30;
wire n_24;
wire n_26;
wire n_27;
wire n_28;
wire n_32;
wire n_11;
wire n_48;
wire n_29;
wire n_35;
wire n_51;
wire n_53;
wire n_55;
wire n_39;
wire n_41;
wire n_42;
wire n_44;
wire n_49;


OR3_X1 i_80 (.ZN (n_56), .A1 (A_imm[9]), .A2 (A_imm[8]), .A3 (A_imm[10]));
NOR2_X2 i_79 (.ZN (n_55), .A1 (A_imm[11]), .A2 (n_56));
OR3_X1 i_78 (.ZN (n_54), .A1 (A_imm[13]), .A2 (A_imm[12]), .A3 (A_imm[14]));
NOR2_X2 i_77 (.ZN (n_53), .A1 (A_imm[15]), .A2 (n_54));
OR3_X1 i_76 (.ZN (n_52), .A1 (A_imm[17]), .A2 (A_imm[16]), .A3 (A_imm[18]));
NOR2_X1 i_75 (.ZN (n_51), .A1 (A_imm[19]), .A2 (n_52));
OR3_X4 i_74 (.ZN (n_50), .A1 (A_imm[5]), .A2 (A_imm[4]), .A3 (A_imm[6]));
NOR2_X4 i_73 (.ZN (n_49), .A1 (A_imm[7]), .A2 (n_50));
NAND2_X4 i_72 (.ZN (n_47), .A1 (n_44), .A2 (n_49));
NOR2_X1 i_71 (.ZN (n_46), .A1 (A_imm[8]), .A2 (n_47));
AOI21_X2 i_70 (.ZN (A_imm_2s_complement[8]), .A (n_46), .B1 (A_imm[8]), .B2 (n_47));
AOI21_X2 i_69 (.ZN (A_imm_2s_complement[3]), .A (n_44), .B1 (A_imm[3]), .B2 (n_42));
INV_X2 i_68 (.ZN (n_45), .A (n_44));
NOR2_X4 i_67 (.ZN (n_44), .A1 (n_42), .A2 (A_imm[3]));
INV_X1 i_66 (.ZN (n_43), .A (n_42));
NAND2_X2 i_65 (.ZN (n_42), .A1 (n_41), .A2 (n_39));
INV_X1 i_64 (.ZN (n_41), .A (A_imm[2]));
NOR2_X4 i_63 (.ZN (n_39), .A1 (A_imm[1]), .A2 (A_imm[0]));
INV_X1 i_62 (.ZN (n_38), .A (n_39));
AOI21_X1 i_61 (.ZN (A_imm_2s_complement[1]), .A (n_39), .B1 (A_imm[1]), .B2 (A_imm[0]));
INV_X1 i_60 (.ZN (n_35), .A (A_imm[22]));
INV_X1 i_59 (.ZN (n_32), .A (A_imm[21]));
INV_X1 i_58 (.ZN (n_11), .A (A_imm[20]));
INV_X4 i_57 (.ZN (n_40), .A (n_47));
NAND2_X4 i_56 (.ZN (n_36), .A1 (n_40), .A2 (n_55));
INV_X4 i_55 (.ZN (n_37), .A (n_36));
NAND2_X4 i_54 (.ZN (n_33), .A1 (n_37), .A2 (n_53));
INV_X4 i_53 (.ZN (n_34), .A (n_33));
NAND2_X4 i_52 (.ZN (n_30), .A1 (n_34), .A2 (n_51));
INV_X4 i_51 (.ZN (n_31), .A (n_30));
NAND4_X2 i_50 (.ZN (n_48), .A1 (n_31), .A2 (n_35), .A3 (n_32), .A4 (n_11));
OR2_X1 i_49 (.ZN (A_imm_2s_complement[27]), .A1 (n_48), .A2 (A_imm[23]));
XNOR2_X1 i_48 (.ZN (n_29), .A (n_48), .B (A_imm[23]));
INV_X1 i_47 (.ZN (A_imm_2s_complement[23]), .A (n_29));
INV_X2 i_46 (.ZN (n_28), .A (n_48));
NAND3_X4 i_45 (.ZN (n_27), .A1 (n_31), .A2 (n_32), .A3 (n_11));
AOI21_X4 i_44 (.ZN (A_imm_2s_complement[22]), .A (n_28), .B1 (n_27), .B2 (A_imm[22]));
INV_X1 i_43 (.ZN (n_26), .A (n_25));
INV_X2 i_42 (.ZN (n_24), .A (n_27));
AOI21_X4 i_41 (.ZN (A_imm_2s_complement[21]), .A (n_24), .B1 (n_26), .B2 (A_imm[21]));
NOR2_X2 i_40 (.ZN (n_25), .A1 (A_imm[20]), .A2 (n_30));
AOI21_X2 i_39 (.ZN (A_imm_2s_complement[20]), .A (n_25), .B1 (A_imm[20]), .B2 (n_30));
NOR2_X4 i_38 (.ZN (n_23), .A1 (A_imm[16]), .A2 (n_33));
INV_X4 i_37 (.ZN (n_22), .A (n_23));
NOR2_X4 i_36 (.ZN (n_21), .A1 (A_imm[17]), .A2 (n_22));
INV_X1 i_35 (.ZN (n_20), .A (n_21));
NOR2_X2 i_34 (.ZN (n_19), .A1 (n_33), .A2 (n_52));
INV_X1 i_33 (.ZN (n_18), .A (n_19));
AOI21_X2 i_32 (.ZN (A_imm_2s_complement[19]), .A (n_31), .B1 (A_imm[19]), .B2 (n_18));
AOI21_X4 i_31 (.ZN (A_imm_2s_complement[18]), .A (n_19), .B1 (A_imm[18]), .B2 (n_20));
AOI21_X2 i_30 (.ZN (A_imm_2s_complement[17]), .A (n_21), .B1 (A_imm[17]), .B2 (n_22));
AOI21_X2 i_29 (.ZN (A_imm_2s_complement[16]), .A (n_23), .B1 (A_imm[16]), .B2 (n_33));
NOR2_X2 i_28 (.ZN (n_17), .A1 (A_imm[12]), .A2 (n_36));
INV_X1 i_27 (.ZN (n_16), .A (n_17));
NOR2_X2 i_26 (.ZN (n_15), .A1 (A_imm[13]), .A2 (n_16));
INV_X1 i_25 (.ZN (n_14), .A (n_15));
NOR2_X1 i_24 (.ZN (n_13), .A1 (n_36), .A2 (n_54));
INV_X1 i_23 (.ZN (n_12), .A (n_13));
AOI21_X2 i_22 (.ZN (A_imm_2s_complement[15]), .A (n_34), .B1 (A_imm[15]), .B2 (n_12));
AOI21_X4 i_21 (.ZN (A_imm_2s_complement[14]), .A (n_13), .B1 (A_imm[14]), .B2 (n_14));
AOI21_X2 i_20 (.ZN (A_imm_2s_complement[13]), .A (n_15), .B1 (A_imm[13]), .B2 (n_16));
AOI21_X2 i_19 (.ZN (A_imm_2s_complement[12]), .A (n_17), .B1 (A_imm[12]), .B2 (n_36));
INV_X1 i_18 (.ZN (n_10), .A (n_46));
NOR2_X2 i_17 (.ZN (n_9), .A1 (A_imm[9]), .A2 (n_10));
INV_X1 i_16 (.ZN (n_8), .A (n_9));
NOR2_X1 i_15 (.ZN (n_7), .A1 (n_47), .A2 (n_56));
INV_X1 i_14 (.ZN (n_6), .A (n_7));
AOI21_X2 i_13 (.ZN (A_imm_2s_complement[11]), .A (n_37), .B1 (A_imm[11]), .B2 (n_6));
AOI21_X2 i_12 (.ZN (A_imm_2s_complement[10]), .A (n_7), .B1 (A_imm[10]), .B2 (n_8));
AOI21_X2 i_11 (.ZN (A_imm_2s_complement[9]), .A (n_9), .B1 (A_imm[9]), .B2 (n_10));
NOR2_X2 i_10 (.ZN (n_5), .A1 (A_imm[4]), .A2 (n_45));
INV_X1 i_9 (.ZN (n_4), .A (n_5));
NOR2_X2 i_8 (.ZN (n_3), .A1 (A_imm[5]), .A2 (n_4));
INV_X1 i_7 (.ZN (n_2), .A (n_3));
NOR2_X1 i_6 (.ZN (n_1), .A1 (n_45), .A2 (n_50));
INV_X1 i_5 (.ZN (n_0), .A (n_1));
AOI21_X2 i_4 (.ZN (A_imm_2s_complement[7]), .A (n_40), .B1 (A_imm[7]), .B2 (n_0));
AOI21_X2 i_3 (.ZN (A_imm_2s_complement[6]), .A (n_1), .B1 (A_imm[6]), .B2 (n_2));
AOI21_X2 i_2 (.ZN (A_imm_2s_complement[5]), .A (n_3), .B1 (A_imm[5]), .B2 (n_4));
AOI21_X2 i_1 (.ZN (A_imm_2s_complement[4]), .A (n_5), .B1 (A_imm[4]), .B2 (n_45));
AOI21_X2 i_0 (.ZN (A_imm_2s_complement[2]), .A (n_43), .B1 (A_imm[2]), .B2 (n_38));

endmodule //datapath__0_0

module boothAlgoR4 (clk_CTS_1_PP_1, clk_CTS_1_PP_9, Res, OVF, A, B, clk, reset, enable);

output OVF;
output [63:0] Res;
output clk_CTS_1_PP_1;
input [31:0] A;
input [31:0] B;
input clk;
input enable;
input reset;
input clk_CTS_1_PP_9;
wire \A_imm_2s_complement[27] ;
wire \A_imm_2s_complement[23] ;
wire \A_imm_2s_complement[22] ;
wire \A_imm_2s_complement[21] ;
wire \A_imm_2s_complement[20] ;
wire \A_imm_2s_complement[19] ;
wire \A_imm_2s_complement[18] ;
wire \A_imm_2s_complement[17] ;
wire \A_imm_2s_complement[16] ;
wire \A_imm_2s_complement[15] ;
wire \A_imm_2s_complement[14] ;
wire \A_imm_2s_complement[13] ;
wire \A_imm_2s_complement[12] ;
wire \A_imm_2s_complement[11] ;
wire \A_imm_2s_complement[10] ;
wire \A_imm_2s_complement[9] ;
wire \A_imm_2s_complement[8] ;
wire \A_imm_2s_complement[7] ;
wire \A_imm_2s_complement[6] ;
wire \A_imm_2s_complement[5] ;
wire \A_imm_2s_complement[4] ;
wire \A_imm_2s_complement[3] ;
wire \A_imm_2s_complement[2] ;
wire \A_imm_2s_complement[1] ;
wire \aggregated_res[14][47] ;
wire \aggregated_res[14][46] ;
wire \aggregated_res[14][45] ;
wire \aggregated_res[14][44] ;
wire \aggregated_res[14][43] ;
wire \aggregated_res[14][42] ;
wire \aggregated_res[14][41] ;
wire \aggregated_res[14][40] ;
wire \aggregated_res[14][39] ;
wire \aggregated_res[14][38] ;
wire \aggregated_res[14][37] ;
wire \aggregated_res[14][36] ;
wire \aggregated_res[14][35] ;
wire \aggregated_res[14][34] ;
wire \aggregated_res[14][33] ;
wire \aggregated_res[14][32] ;
wire \aggregated_res[14][31] ;
wire \aggregated_res[14][30] ;
wire \aggregated_res[14][29] ;
wire \aggregated_res[14][28] ;
wire \aggregated_res[14][27] ;
wire \aggregated_res[14][26] ;
wire \aggregated_res[14][25] ;
wire \aggregated_res[14][24] ;
wire \aggregated_res[14][23] ;
wire drc_ipo_n30;
wire drc_ipo_n31;
wire drc_ipo_n32;
wire CTS_n_tid1_52;
wire spc__n131;
wire spc__n134;
wire spc__n136;
wire hfn_ipo_n29;
wire hfn_ipo_n28;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_32;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_58;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_89;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_122;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_153;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_169;
wire n_0_170;
wire n_0_171;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_176;
wire n_0_177;
wire n_0_178;
wire n_0_179;
wire n_0_180;
wire n_0_184;
wire n_0_190;
wire n_0_191;
wire n_0_192;
wire n_0_193;
wire n_0_194;
wire n_0_195;
wire n_0_196;
wire n_0_197;
wire n_0_198;
wire n_0_199;
wire n_0_200;
wire n_0_201;
wire n_0_203;
wire n_0_204;
wire n_0_205;
wire n_0_207;
wire n_0_208;
wire n_0_209;
wire n_0_210;
wire n_0_211;
wire n_0_215;
wire n_0_221;
wire n_0_222;
wire n_0_223;
wire n_0_224;
wire n_0_225;
wire n_0_226;
wire n_0_227;
wire n_0_228;
wire n_0_229;
wire n_0_230;
wire n_0_231;
wire n_0_232;
wire n_0_233;
wire n_0_234;
wire n_0_235;
wire n_0_236;
wire n_0_237;
wire n_0_238;
wire n_0_239;
wire n_0_240;
wire n_0_241;
wire n_0_242;
wire n_0_246;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_255;
wire n_0_256;
wire n_0_257;
wire n_0_258;
wire n_0_259;
wire n_0_260;
wire n_0_261;
wire n_0_262;
wire n_0_263;
wire n_0_264;
wire n_0_265;
wire n_0_266;
wire n_0_267;
wire n_0_269;
wire n_0_270;
wire n_0_271;
wire n_0_272;
wire n_0_273;
wire n_0_277;
wire n_0_283;
wire n_0_284;
wire n_0_285;
wire n_0_286;
wire n_0_287;
wire n_0_288;
wire n_0_289;
wire n_0_290;
wire n_0_291;
wire n_0_292;
wire n_0_293;
wire n_0_294;
wire n_0_295;
wire n_0_296;
wire n_0_297;
wire n_0_298;
wire n_0_299;
wire n_0_300;
wire n_0_302;
wire n_0_303;
wire n_0_308;
wire n_0_314;
wire n_0_315;
wire n_0_316;
wire n_0_317;
wire n_0_318;
wire n_0_319;
wire n_0_320;
wire n_0_321;
wire n_0_322;
wire n_0_323;
wire n_0_324;
wire n_0_325;
wire n_0_326;
wire n_0_327;
wire n_0_328;
wire n_0_329;
wire n_0_331;
wire n_0_332;
wire n_0_333;
wire n_0_335;
wire n_0_339;
wire n_0_344;
wire n_0_346;
wire n_0_347;
wire n_0_348;
wire n_0_349;
wire n_0_350;
wire n_0_351;
wire n_0_352;
wire n_0_353;
wire n_0_354;
wire n_0_355;
wire n_0_356;
wire n_0_357;
wire n_0_359;
wire n_0_360;
wire n_0_361;
wire n_0_363;
wire n_0_365;
wire n_0_369;
wire n_0_370;
wire n_0_371;
wire n_0_372;
wire n_0_373;
wire n_0_374;
wire n_0_375;
wire n_0_376;
wire n_0_377;
wire n_0_378;
wire n_0_379;
wire n_0_380;
wire n_0_382;
wire n_0_383;
wire n_0_384;
wire n_0_386;
wire n_0_388;
wire n_0_391;
wire n_0_385;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_33;
wire n_0_34;
wire n_0_57;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_88;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_181;
wire n_0_182;
wire n_0_183;
wire n_0_185;
wire n_0_186;
wire n_0_187;
wire n_0_188;
wire n_0_189;
wire n_0_202;
wire n_0_206;
wire n_0_212;
wire n_0_213;
wire n_0_214;
wire n_0_216;
wire n_0_217;
wire n_0_218;
wire n_0_219;
wire n_0_220;
wire n_0_243;
wire n_0_244;
wire n_0_245;
wire n_0_247;
wire n_0_248;
wire n_0_249;
wire n_0_250;
wire n_0_251;
wire n_0_268;
wire n_0_274;
wire n_0_275;
wire n_0_276;
wire n_0_278;
wire n_0_279;
wire n_0_280;
wire n_0_281;
wire n_0_282;
wire n_0_301;
wire n_0_304;
wire n_0_305;
wire n_0_306;
wire n_0_307;
wire n_0_310;
wire n_0_311;
wire n_0_312;
wire n_0_313;
wire n_0_330;
wire n_0_334;
wire n_0_336;
wire n_0_337;
wire n_0_338;
wire n_0_340;
wire n_0_341;
wire n_0_342;
wire n_0_343;
wire n_0_345;
wire n_0_358;
wire n_0_362;
wire n_0_364;
wire n_0_366;
wire n_0_367;
wire n_0_368;
wire n_0_381;
wire n_0_387;
wire n_0_389;
wire n_0_390;
wire n_0_392;
wire n_0_393;
wire n_0_394;
wire n_0_395;
wire n_0_396;
wire n_0_397;
wire n_0_398;
wire n_0_399;
wire n_0_400;
wire n_0_401;
wire n_0_402;
wire n_0_403;
wire n_0_404;
wire n_0_405;
wire n_0_406;
wire n_0_407;
wire n_0_408;
wire n_0_409;
wire n_0_410;
wire n_0_411;
wire n_0_412;
wire n_0_413;
wire n_0_414;
wire n_0_415;
wire n_0_416;
wire n_0_417;
wire n_0_418;
wire CTS_n39;
wire n_1_0__1;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire n_46;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire uc_28;
wire uc_29;
wire uc_30;
wire uc_31;
wire uc_32;
wire uc_33;
wire uc_34;
wire uc_35;
wire uc_36;
wire uc_37;
wire uc_38;
wire uc_39;
wire uc_40;
wire uc_41;
wire uc_42;
wire uc_43;
wire uc_44;
wire n_361;
wire uc_45;
wire uc_46;
wire uc_47;
wire uc_48;
wire uc_49;
wire uc_50;
wire uc_51;
wire n_360;
wire n_359;
wire n_379;
wire n_358;
wire n_357;
wire n_356;
wire n_378;
wire n_355;
wire n_354;
wire n_353;
wire n_352;
wire n_351;
wire n_350;
wire n_349;
wire n_348;
wire n_347;
wire n_346;
wire n_345;
wire n_344;
wire n_343;
wire n_342;
wire n_341;
wire n_340;
wire n_377;
wire n_339;
wire uc_52;
wire uc_53;
wire uc_54;
wire uc_55;
wire uc_56;
wire uc_57;
wire uc_58;
wire uc_59;
wire uc_60;
wire uc_61;
wire uc_62;
wire uc_63;
wire uc_64;
wire uc_65;
wire uc_66;
wire uc_67;
wire uc_68;
wire uc_69;
wire uc_70;
wire uc_71;
wire uc_72;
wire uc_73;
wire uc_74;
wire uc_75;
wire uc_76;
wire uc_77;
wire uc_78;
wire uc_79;
wire uc_80;
wire n_338;
wire uc_81;
wire uc_82;
wire uc_83;
wire uc_84;
wire uc_85;
wire uc_86;
wire uc_87;
wire n_337;
wire n_376;
wire n_336;
wire n_335;
wire n_375;
wire n_334;
wire n_333;
wire n_332;
wire n_331;
wire n_330;
wire n_329;
wire n_328;
wire n_327;
wire n_326;
wire n_325;
wire n_324;
wire n_323;
wire n_322;
wire n_321;
wire n_320;
wire n_319;
wire n_318;
wire n_317;
wire n_374;
wire n_316;
wire uc_88;
wire uc_89;
wire uc_90;
wire uc_91;
wire uc_92;
wire uc_93;
wire uc_94;
wire uc_95;
wire uc_96;
wire uc_97;
wire uc_98;
wire uc_99;
wire uc_100;
wire uc_101;
wire uc_102;
wire uc_103;
wire uc_104;
wire uc_105;
wire uc_106;
wire uc_107;
wire uc_108;
wire uc_109;
wire uc_110;
wire uc_111;
wire uc_112;
wire uc_113;
wire uc_114;
wire uc_115;
wire uc_116;
wire n_315;
wire uc_117;
wire uc_118;
wire uc_119;
wire uc_120;
wire uc_121;
wire uc_122;
wire uc_123;
wire n_314;
wire n_313;
wire n_312;
wire n_311;
wire n_310;
wire n_309;
wire n_373;
wire n_308;
wire n_307;
wire n_306;
wire n_305;
wire n_304;
wire n_303;
wire n_302;
wire n_301;
wire n_300;
wire n_299;
wire n_298;
wire n_297;
wire n_296;
wire n_295;
wire n_294;
wire n_293;
wire n_372;
wire n_292;
wire uc_124;
wire uc_125;
wire uc_126;
wire uc_127;
wire uc_128;
wire uc_129;
wire uc_130;
wire uc_131;
wire uc_132;
wire uc_133;
wire uc_134;
wire uc_135;
wire uc_136;
wire uc_137;
wire uc_138;
wire uc_139;
wire uc_140;
wire uc_141;
wire uc_142;
wire uc_143;
wire uc_144;
wire uc_145;
wire uc_146;
wire uc_147;
wire uc_148;
wire uc_149;
wire uc_150;
wire uc_151;
wire uc_152;
wire n_291;
wire uc_153;
wire uc_154;
wire uc_155;
wire uc_156;
wire uc_157;
wire uc_158;
wire uc_159;
wire n_290;
wire n_289;
wire n_288;
wire n_287;
wire n_286;
wire n_285;
wire n_284;
wire n_283;
wire n_282;
wire n_281;
wire n_280;
wire n_279;
wire n_278;
wire n_277;
wire n_276;
wire n_275;
wire n_274;
wire n_273;
wire n_272;
wire n_271;
wire n_270;
wire n_269;
wire n_268;
wire n_371;
wire n_267;
wire uc_160;
wire uc_161;
wire uc_162;
wire uc_163;
wire uc_164;
wire uc_165;
wire uc_166;
wire uc_167;
wire uc_168;
wire uc_169;
wire uc_170;
wire uc_171;
wire uc_172;
wire uc_173;
wire uc_174;
wire uc_175;
wire uc_176;
wire uc_177;
wire uc_178;
wire uc_179;
wire uc_180;
wire uc_181;
wire uc_182;
wire uc_183;
wire uc_184;
wire uc_185;
wire uc_186;
wire uc_187;
wire uc_188;
wire n_266;
wire uc_189;
wire uc_190;
wire uc_191;
wire uc_192;
wire uc_193;
wire uc_194;
wire uc_195;
wire n_265;
wire n_264;
wire n_263;
wire n_262;
wire n_261;
wire n_260;
wire n_370;
wire n_259;
wire n_258;
wire n_257;
wire n_369;
wire n_256;
wire n_255;
wire n_254;
wire n_253;
wire n_252;
wire n_251;
wire n_250;
wire n_249;
wire n_248;
wire n_247;
wire n_246;
wire n_245;
wire n_368;
wire n_244;
wire uc_196;
wire uc_197;
wire uc_198;
wire uc_199;
wire uc_200;
wire uc_201;
wire uc_202;
wire uc_203;
wire uc_204;
wire uc_205;
wire uc_206;
wire uc_207;
wire uc_208;
wire uc_209;
wire uc_210;
wire uc_211;
wire uc_212;
wire uc_213;
wire uc_214;
wire uc_215;
wire uc_216;
wire uc_217;
wire uc_218;
wire uc_219;
wire uc_220;
wire uc_221;
wire uc_222;
wire uc_223;
wire uc_224;
wire uc_225;
wire n_243;
wire uc_226;
wire uc_227;
wire uc_228;
wire uc_229;
wire uc_230;
wire uc_231;
wire n_242;
wire n_241;
wire n_240;
wire n_239;
wire n_238;
wire n_237;
wire n_236;
wire n_235;
wire n_234;
wire n_233;
wire n_232;
wire n_231;
wire n_230;
wire n_229;
wire n_228;
wire n_227;
wire n_226;
wire n_225;
wire n_224;
wire n_223;
wire n_222;
wire n_221;
wire n_220;
wire n_367;
wire n_219;
wire uc_232;
wire uc_233;
wire uc_234;
wire uc_235;
wire uc_236;
wire uc_237;
wire uc_238;
wire uc_239;
wire uc_240;
wire uc_241;
wire uc_242;
wire uc_243;
wire uc_244;
wire uc_245;
wire uc_246;
wire uc_247;
wire uc_248;
wire uc_249;
wire uc_250;
wire uc_251;
wire uc_252;
wire uc_253;
wire uc_254;
wire uc_255;
wire uc_256;
wire uc_257;
wire uc_258;
wire uc_259;
wire uc_260;
wire uc_261;
wire n_218;
wire uc_262;
wire uc_263;
wire uc_264;
wire uc_265;
wire uc_266;
wire uc_267;
wire n_217;
wire n_216;
wire n_215;
wire n_214;
wire n_213;
wire n_212;
wire n_211;
wire n_210;
wire n_209;
wire n_208;
wire n_207;
wire n_206;
wire n_205;
wire n_204;
wire n_203;
wire n_202;
wire n_201;
wire n_200;
wire n_199;
wire n_198;
wire n_197;
wire n_196;
wire n_195;
wire n_366;
wire n_194;
wire uc_268;
wire uc_269;
wire uc_270;
wire uc_271;
wire uc_272;
wire uc_273;
wire uc_274;
wire uc_275;
wire uc_276;
wire uc_277;
wire uc_278;
wire uc_279;
wire uc_280;
wire uc_281;
wire uc_282;
wire uc_283;
wire uc_284;
wire uc_285;
wire uc_286;
wire uc_287;
wire uc_288;
wire uc_289;
wire uc_290;
wire uc_291;
wire uc_292;
wire uc_293;
wire uc_294;
wire uc_295;
wire uc_296;
wire uc_297;
wire uc_298;
wire uc_299;
wire n_193;
wire uc_300;
wire uc_301;
wire uc_302;
wire uc_303;
wire n_192;
wire n_191;
wire n_190;
wire n_189;
wire n_188;
wire n_187;
wire n_186;
wire n_185;
wire n_184;
wire n_183;
wire n_182;
wire n_181;
wire n_180;
wire n_179;
wire n_178;
wire n_177;
wire n_176;
wire n_175;
wire n_174;
wire n_173;
wire n_172;
wire n_171;
wire n_170;
wire n_365;
wire n_169;
wire uc_304;
wire uc_305;
wire uc_306;
wire uc_307;
wire uc_308;
wire uc_309;
wire uc_310;
wire uc_311;
wire uc_312;
wire uc_313;
wire uc_314;
wire uc_315;
wire uc_316;
wire uc_317;
wire uc_318;
wire uc_319;
wire uc_320;
wire uc_321;
wire uc_322;
wire uc_323;
wire uc_324;
wire uc_325;
wire uc_326;
wire uc_327;
wire uc_328;
wire uc_329;
wire uc_330;
wire uc_331;
wire uc_332;
wire uc_333;
wire uc_334;
wire uc_335;
wire uc_336;
wire uc_337;
wire n_168;
wire uc_338;
wire uc_339;
wire n_167;
wire n_166;
wire n_165;
wire n_164;
wire n_163;
wire n_162;
wire n_161;
wire n_160;
wire n_159;
wire n_158;
wire n_157;
wire n_156;
wire n_155;
wire n_154;
wire n_153;
wire n_152;
wire n_151;
wire n_150;
wire n_149;
wire n_148;
wire n_147;
wire n_146;
wire n_145;
wire n_364;
wire n_144;
wire uc_340;
wire uc_341;
wire uc_342;
wire uc_343;
wire uc_344;
wire uc_345;
wire uc_346;
wire uc_347;
wire uc_348;
wire uc_349;
wire uc_350;
wire uc_351;
wire uc_352;
wire uc_353;
wire uc_354;
wire uc_355;
wire uc_356;
wire uc_357;
wire uc_358;
wire uc_359;
wire uc_360;
wire uc_361;
wire uc_362;
wire uc_363;
wire uc_364;
wire uc_365;
wire uc_366;
wire uc_367;
wire uc_368;
wire uc_369;
wire uc_370;
wire uc_371;
wire uc_372;
wire uc_373;
wire uc_374;
wire uc_375;
wire n_143;
wire n_142;
wire n_141;
wire n_140;
wire n_139;
wire n_138;
wire n_137;
wire n_136;
wire n_135;
wire n_134;
wire n_133;
wire n_132;
wire n_131;
wire n_130;
wire n_129;
wire n_128;
wire n_127;
wire n_126;
wire n_125;
wire n_124;
wire n_123;
wire n_122;
wire n_121;
wire n_120;
wire n_363;
wire n_119;
wire uc_376;
wire uc_377;
wire uc_378;
wire uc_379;
wire uc_380;
wire uc_381;
wire uc_382;
wire uc_383;
wire uc_384;
wire uc_385;
wire uc_386;
wire uc_387;
wire uc_388;
wire uc_389;
wire uc_390;
wire uc_391;
wire uc_392;
wire uc_393;
wire uc_394;
wire uc_395;
wire uc_396;
wire uc_397;
wire uc_398;
wire uc_399;
wire uc_400;
wire uc_401;
wire uc_402;
wire uc_403;
wire uc_404;
wire uc_405;
wire uc_406;
wire uc_407;
wire uc_408;
wire uc_409;
wire uc_410;
wire uc_411;
wire n_118;
wire n_117;
wire n_362;
wire n_116;
wire n_115;
wire n_114;
wire n_113;
wire n_112;
wire n_111;
wire n_110;
wire n_109;
wire n_108;
wire n_107;
wire n_106;
wire n_105;
wire n_104;
wire n_103;
wire n_102;
wire n_101;
wire n_100;
wire n_99;
wire n_98;
wire n_97;
wire n_96;
wire n_95;
wire n_94;
wire uc_412;
wire uc_413;
wire uc_414;
wire uc_415;
wire uc_416;
wire uc_417;
wire uc_418;
wire uc_419;
wire uc_420;
wire uc_421;
wire uc_422;
wire uc_423;
wire uc_424;
wire uc_425;
wire uc_426;
wire uc_427;
wire uc_428;
wire uc_429;
wire uc_430;
wire uc_431;
wire uc_432;
wire uc_433;
wire uc_434;
wire uc_435;
wire uc_436;
wire uc_437;
wire uc_438;
wire uc_439;
wire uc_440;
wire uc_441;
wire uc_442;
wire uc_443;
wire uc_444;
wire uc_445;
wire uc_446;
wire uc_447;
wire uc_448;
wire uc_449;
wire n_93;
wire n_92;
wire n_91;
wire n_90;
wire n_89;
wire n_88;
wire n_87;
wire n_86;
wire n_85;
wire n_84;
wire n_83;
wire n_82;
wire n_81;
wire n_80;
wire n_79;
wire n_78;
wire n_77;
wire n_76;
wire n_75;
wire n_74;
wire n_73;
wire n_72;
wire n_71;
wire uc_450;
wire uc_451;
wire uc_452;
wire uc_453;
wire uc_454;
wire uc_455;
wire uc_456;
wire uc_457;
wire uc_458;
wire uc_459;
wire uc_460;
wire uc_461;
wire uc_462;
wire uc_463;
wire uc_464;
wire uc_465;
wire uc_466;
wire uc_467;
wire uc_468;
wire uc_469;
wire uc_470;
wire uc_471;
wire uc_472;
wire uc_473;
wire uc_474;
wire uc_475;
wire uc_476;
wire uc_477;
wire uc_478;
wire uc_479;
wire uc_480;
wire uc_481;
wire uc_482;
wire uc_483;
wire uc_484;
wire uc_485;
wire uc_486;
wire uc_487;
wire uc_488;
wire uc_489;
wire uc_490;
wire uc_491;
wire uc_492;
wire uc_493;
wire uc_494;
wire uc_495;
wire uc_496;
wire uc_497;
wire uc_498;
wire uc_499;
wire uc_500;
wire uc_501;
wire uc_502;
wire uc_503;
wire uc_504;
wire n_70;
wire uc_505;
wire uc_506;
wire uc_507;
wire uc_508;
wire uc_509;
wire uc_510;
wire uc_511;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire uc_512;
wire uc_513;
wire uc_514;
wire uc_515;
wire uc_516;
wire uc_517;
wire uc_518;
wire uc_519;
wire uc_520;
wire uc_521;
wire uc_522;
wire uc_523;
wire uc_524;
wire uc_525;
wire uc_526;
wire uc_527;
wire uc_528;
wire uc_529;
wire uc_530;
wire uc_531;
wire uc_532;
wire uc_533;
wire uc_534;
wire uc_535;
wire uc_536;
wire uc_537;
wire uc_538;
wire uc_539;
wire uc_540;
wire uc_541;
wire uc_542;
wire uc_543;
wire uc_544;
wire uc_545;
wire uc_546;
wire uc_547;
wire uc_548;
wire uc_549;
wire uc_550;
wire uc_551;
wire uc_552;
wire n_404;
wire n_452;
wire n_403;
wire n_402;
wire n_401;
wire n_400;
wire n_399;
wire n_398;
wire n_397;
wire n_396;
wire n_395;
wire n_394;
wire n_393;
wire n_392;
wire n_391;
wire n_390;
wire n_389;
wire n_388;
wire n_387;
wire n_386;
wire n_385;
wire n_384;
wire n_383;
wire n_382;
wire n_381;
wire n_380;
wire n_451;
wire CTS_n38;
wire n_450;
wire n_449;
wire n_448;
wire n_447;
wire n_446;
wire n_445;
wire n_444;
wire n_443;
wire n_442;
wire n_441;
wire n_440;
wire n_439;
wire n_438;
wire n_437;
wire n_436;
wire n_435;
wire n_434;
wire n_433;
wire n_432;
wire n_431;
wire n_430;
wire n_429;
wire n_427;
wire n_23;
wire n_426;
wire n_24;
wire n_425;
wire n_25;
wire n_424;
wire n_26;
wire n_423;
wire n_27;
wire n_422;
wire n_28;
wire n_421;
wire n_29;
wire n_420;
wire n_30;
wire n_419;
wire n_31;
wire n_418;
wire n_32;
wire n_417;
wire n_33;
wire n_416;
wire n_34;
wire n_415;
wire n_35;
wire n_414;
wire n_36;
wire n_413;
wire n_37;
wire n_412;
wire n_38;
wire n_411;
wire n_39;
wire n_410;
wire n_40;
wire n_409;
wire n_41;
wire n_408;
wire n_42;
wire n_407;
wire n_43;
wire n_406;
wire n_44;
wire n_405;
wire n_45;


INV_X1 i_1_74 (.ZN (n_1_0__1), .A (reset));
NAND2_X2 i_1_73 (.ZN (n_452), .A1 (hfn_ipo_n28), .A2 (CTS_n_tid1_52));
AND2_X1 i_1_72 (.ZN (n_451), .A1 (hfn_ipo_n28), .A2 (A[22]));
AND2_X1 i_1_71 (.ZN (n_450), .A1 (hfn_ipo_n28), .A2 (A[21]));
AND2_X1 i_1_70 (.ZN (n_449), .A1 (hfn_ipo_n28), .A2 (A[20]));
AND2_X1 i_1_69 (.ZN (n_448), .A1 (hfn_ipo_n28), .A2 (A[19]));
AND2_X1 i_1_68 (.ZN (n_447), .A1 (hfn_ipo_n28), .A2 (A[18]));
AND2_X1 i_1_67 (.ZN (n_446), .A1 (hfn_ipo_n28), .A2 (A[17]));
AND2_X1 i_1_66 (.ZN (n_445), .A1 (hfn_ipo_n28), .A2 (A[16]));
AND2_X1 i_1_65 (.ZN (n_444), .A1 (hfn_ipo_n28), .A2 (A[15]));
AND2_X1 i_1_64 (.ZN (n_443), .A1 (hfn_ipo_n28), .A2 (A[14]));
AND2_X1 i_1_63 (.ZN (n_442), .A1 (hfn_ipo_n28), .A2 (A[13]));
AND2_X1 i_1_62 (.ZN (n_441), .A1 (hfn_ipo_n28), .A2 (A[12]));
AND2_X1 i_1_61 (.ZN (n_440), .A1 (hfn_ipo_n28), .A2 (A[11]));
AND2_X1 i_1_60 (.ZN (n_439), .A1 (hfn_ipo_n28), .A2 (A[10]));
AND2_X1 i_1_59 (.ZN (n_438), .A1 (hfn_ipo_n28), .A2 (A[9]));
AND2_X1 i_1_58 (.ZN (n_437), .A1 (hfn_ipo_n28), .A2 (A[8]));
AND2_X1 i_1_57 (.ZN (n_436), .A1 (hfn_ipo_n28), .A2 (A[7]));
AND2_X1 i_1_56 (.ZN (n_435), .A1 (hfn_ipo_n28), .A2 (A[6]));
AND2_X1 i_1_55 (.ZN (n_434), .A1 (hfn_ipo_n28), .A2 (A[5]));
AND2_X1 i_1_54 (.ZN (n_433), .A1 (hfn_ipo_n28), .A2 (A[4]));
AND2_X1 i_1_53 (.ZN (n_432), .A1 (hfn_ipo_n28), .A2 (A[3]));
AND2_X1 i_1_52 (.ZN (n_431), .A1 (hfn_ipo_n28), .A2 (A[2]));
AND2_X1 i_1_51 (.ZN (n_430), .A1 (hfn_ipo_n28), .A2 (A[1]));
AND2_X1 i_1_50 (.ZN (n_429), .A1 (hfn_ipo_n28), .A2 (A[0]));
AOI21_X1 i_1_49 (.ZN (CTS_n39), .A (reset), .B1 (clk_CTS_1_PP_1), .B2 (enable));
INV_X4 CTS_L3_remove_c41 (.ZN (CTS_n38), .A (CTS_n39));
AND2_X1 i_1_47 (.ZN (n_427), .A1 (hfn_ipo_n29), .A2 (B[22]));
AND2_X1 i_1_46 (.ZN (n_426), .A1 (hfn_ipo_n29), .A2 (B[21]));
AND2_X1 i_1_45 (.ZN (n_425), .A1 (hfn_ipo_n29), .A2 (B[20]));
AND2_X1 i_1_44 (.ZN (n_424), .A1 (hfn_ipo_n29), .A2 (B[19]));
AND2_X1 i_1_43 (.ZN (n_423), .A1 (hfn_ipo_n29), .A2 (B[18]));
AND2_X1 i_1_42 (.ZN (n_422), .A1 (hfn_ipo_n29), .A2 (B[17]));
AND2_X1 i_1_41 (.ZN (n_421), .A1 (hfn_ipo_n29), .A2 (B[16]));
AND2_X1 i_1_40 (.ZN (n_420), .A1 (hfn_ipo_n29), .A2 (B[15]));
AND2_X1 i_1_39 (.ZN (n_419), .A1 (hfn_ipo_n29), .A2 (B[14]));
AND2_X1 i_1_38 (.ZN (n_418), .A1 (hfn_ipo_n29), .A2 (B[13]));
AND2_X1 i_1_37 (.ZN (n_417), .A1 (hfn_ipo_n29), .A2 (B[12]));
AND2_X1 i_1_36 (.ZN (n_416), .A1 (hfn_ipo_n29), .A2 (B[11]));
AND2_X1 i_1_35 (.ZN (n_415), .A1 (hfn_ipo_n29), .A2 (B[10]));
AND2_X1 i_1_34 (.ZN (n_414), .A1 (hfn_ipo_n29), .A2 (B[9]));
AND2_X1 i_1_33 (.ZN (n_413), .A1 (hfn_ipo_n29), .A2 (B[8]));
AND2_X1 i_1_32 (.ZN (n_412), .A1 (hfn_ipo_n29), .A2 (B[7]));
AND2_X1 i_1_31 (.ZN (n_411), .A1 (hfn_ipo_n29), .A2 (B[6]));
AND2_X1 i_1_30 (.ZN (n_410), .A1 (hfn_ipo_n29), .A2 (B[5]));
AND2_X1 i_1_29 (.ZN (n_409), .A1 (hfn_ipo_n29), .A2 (B[4]));
AND2_X1 i_1_28 (.ZN (n_408), .A1 (hfn_ipo_n29), .A2 (B[3]));
AND2_X1 i_1_27 (.ZN (n_407), .A1 (hfn_ipo_n29), .A2 (B[2]));
AND2_X1 i_1_26 (.ZN (n_406), .A1 (hfn_ipo_n29), .A2 (B[1]));
AND2_X1 i_1_25 (.ZN (n_405), .A1 (hfn_ipo_n29), .A2 (B[0]));
AND2_X1 i_1_24 (.ZN (n_404), .A1 (hfn_ipo_n29), .A2 (\aggregated_res[14][47] ));
AND2_X1 i_1_23 (.ZN (n_403), .A1 (hfn_ipo_n29), .A2 (\aggregated_res[14][46] ));
AND2_X1 i_1_22 (.ZN (n_402), .A1 (hfn_ipo_n29), .A2 (\aggregated_res[14][45] ));
AND2_X1 i_1_21 (.ZN (n_401), .A1 (hfn_ipo_n29), .A2 (\aggregated_res[14][44] ));
AND2_X1 i_1_20 (.ZN (n_400), .A1 (hfn_ipo_n29), .A2 (\aggregated_res[14][43] ));
AND2_X1 i_1_19 (.ZN (n_399), .A1 (hfn_ipo_n29), .A2 (\aggregated_res[14][42] ));
AND2_X1 i_1_18 (.ZN (n_398), .A1 (hfn_ipo_n29), .A2 (\aggregated_res[14][41] ));
AND2_X1 i_1_17 (.ZN (n_397), .A1 (hfn_ipo_n29), .A2 (\aggregated_res[14][40] ));
AND2_X1 i_1_16 (.ZN (n_396), .A1 (hfn_ipo_n29), .A2 (\aggregated_res[14][39] ));
AND2_X1 i_1_15 (.ZN (n_395), .A1 (hfn_ipo_n29), .A2 (\aggregated_res[14][38] ));
AND2_X1 i_1_14 (.ZN (n_394), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][37] ));
AND2_X1 i_1_13 (.ZN (n_393), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][36] ));
AND2_X1 i_1_12 (.ZN (n_392), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][35] ));
AND2_X1 i_1_11 (.ZN (n_391), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][34] ));
AND2_X1 i_1_10 (.ZN (n_390), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][33] ));
AND2_X1 i_1_9 (.ZN (n_389), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][32] ));
AND2_X1 i_1_8 (.ZN (n_388), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][31] ));
AND2_X1 i_1_7 (.ZN (n_387), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][30] ));
AND2_X1 i_1_6 (.ZN (n_386), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][29] ));
AND2_X1 i_1_5 (.ZN (n_385), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][28] ));
AND2_X1 i_1_4 (.ZN (n_384), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][27] ));
AND2_X1 i_1_3 (.ZN (n_383), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][26] ));
AND2_X1 i_1_2 (.ZN (n_382), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][25] ));
AND2_X1 i_1_1 (.ZN (n_381), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][24] ));
AND2_X1 i_1_0 (.ZN (n_380), .A1 (hfn_ipo_n28), .A2 (\aggregated_res[14][23] ));
AOI22_X1 i_0_751 (.ZN (n_0_418), .A1 (\A_imm_2s_complement[21] ), .A2 (n_0_406), .B1 (n_0_411), .B2 (n_1));
OAI221_X1 i_0_750 (.ZN (n_379), .A (n_0_418), .B1 (n_0_27), .B2 (n_0_414), .C1 (n_0_415), .C2 (n_0_31));
AOI22_X1 i_0_749 (.ZN (n_0_417), .A1 (\A_imm_2s_complement[18] ), .A2 (n_0_413), .B1 (\A_imm_2s_complement[17] ), .B2 (n_0_406));
OAI221_X1 i_0_748 (.ZN (n_378), .A (n_0_417), .B1 (n_0_415), .B2 (n_0_310), .C1 (n_0_410), .C2 (n_0_361));
OAI221_X1 i_0_747 (.ZN (n_377), .A (n_0_416), .B1 (n_0_415), .B2 (n_0_95), .C1 (n_0_414), .C2 (n_0_92));
OAI21_X1 i_0_746 (.ZN (n_0_416), .A (n_22), .B1 (n_0_411), .B2 (n_0_406));
OR2_X2 i_0_745 (.ZN (n_0_415), .A1 (n_0_412), .A2 (n_42));
INV_X2 i_0_744 (.ZN (n_0_414), .A (n_0_413));
NOR2_X1 i_0_743 (.ZN (n_0_413), .A1 (n_0_412), .A2 (n_0_392));
OAI21_X1 i_0_742 (.ZN (n_0_412), .A (n_0_408), .B1 (n_43), .B2 (n_44));
INV_X1 i_0_741 (.ZN (n_0_411), .A (n_0_410));
NAND2_X1 i_0_740 (.ZN (n_0_410), .A1 (n_0_409), .A2 (n_0_392));
INV_X1 i_0_739 (.ZN (n_0_409), .A (n_0_408));
NAND2_X1 i_0_738 (.ZN (n_0_408), .A1 (n_43), .A2 (n_44));
INV_X1 i_0_737 (.ZN (n_0_407), .A (n_44));
NOR3_X4 i_0_736 (.ZN (n_0_406), .A1 (n_43), .A2 (n_44), .A3 (n_0_392));
AOI22_X1 i_0_735 (.ZN (n_0_405), .A1 (\A_imm_2s_complement[23] ), .A2 (n_0_398), .B1 (\A_imm_2s_complement[22] ), .B2 (n_0_390));
OAI221_X1 i_0_734 (.ZN (n_376), .A (n_0_405), .B1 (n_0_400), .B2 (n_0_28), .C1 (n_0_395), .C2 (n_0_31));
INV_X1 i_0_733 (.ZN (n_0_404), .A (n_2));
INV_X4 i_0_732 (.ZN (n_0_403), .A (\A_imm_2s_complement[20] ));
AOI22_X1 i_0_731 (.ZN (n_0_402), .A1 (\A_imm_2s_complement[19] ), .A2 (n_0_390), .B1 (n_0_396), .B2 (n_3));
OAI221_X1 i_0_730 (.ZN (n_375), .A (n_0_402), .B1 (n_0_403), .B2 (n_0_399), .C1 (n_0_404), .C2 (n_0_400));
OAI221_X1 i_0_729 (.ZN (n_374), .A (n_0_401), .B1 (n_0_400), .B2 (n_0_95), .C1 (n_0_399), .C2 (n_0_92));
OAI21_X1 i_0_728 (.ZN (n_0_401), .A (n_22), .B1 (n_0_396), .B2 (n_0_390));
OR2_X2 i_0_727 (.ZN (n_0_400), .A1 (n_0_397), .A2 (n_40));
INV_X2 i_0_726 (.ZN (n_0_399), .A (n_0_398));
NOR2_X1 i_0_725 (.ZN (n_0_398), .A1 (n_0_397), .A2 (n_0_343));
OAI21_X1 i_0_724 (.ZN (n_0_397), .A (n_0_393), .B1 (n_41), .B2 (n_42));
INV_X2 i_0_723 (.ZN (n_0_396), .A (n_0_395));
NAND2_X1 i_0_722 (.ZN (n_0_395), .A1 (n_0_394), .A2 (n_0_343));
INV_X1 i_0_720 (.ZN (n_0_394), .A (n_0_393));
NAND2_X1 i_0_718 (.ZN (n_0_393), .A1 (n_41), .A2 (n_42));
INV_X1 i_0_714 (.ZN (n_0_392), .A (n_42));
NOR3_X4 i_0_702 (.ZN (n_0_390), .A1 (n_41), .A2 (n_42), .A3 (n_0_343));
AOI22_X1 i_0_701 (.ZN (n_0_389), .A1 (\A_imm_2s_complement[18] ), .A2 (n_0_367), .B1 (\A_imm_2s_complement[17] ), .B2 (n_0_342));
OAI221_X1 i_0_700 (.ZN (n_373), .A (n_0_389), .B1 (n_0_381), .B2 (n_0_310), .C1 (n_0_362), .C2 (n_0_361));
OAI221_X1 i_0_699 (.ZN (n_372), .A (n_0_387), .B1 (n_0_381), .B2 (n_0_95), .C1 (n_0_368), .C2 (n_0_92));
OAI21_X1 i_0_697 (.ZN (n_0_387), .A (n_22), .B1 (n_0_364), .B2 (n_0_342));
OR2_X2 i_0_695 (.ZN (n_0_381), .A1 (n_0_366), .A2 (n_38));
INV_X2 i_0_691 (.ZN (n_0_368), .A (n_0_367));
NOR2_X1 i_0_679 (.ZN (n_0_367), .A1 (n_0_366), .A2 (n_0_312));
OAI21_X1 i_0_678 (.ZN (n_0_366), .A (n_0_345), .B1 (n_39), .B2 (n_40));
INV_X2 i_0_677 (.ZN (n_0_364), .A (n_0_362));
NAND2_X1 i_0_676 (.ZN (n_0_362), .A1 (n_0_358), .A2 (n_0_312));
INV_X1 i_0_674 (.ZN (n_0_358), .A (n_0_345));
NAND2_X1 i_0_673 (.ZN (n_0_345), .A1 (n_39), .A2 (n_40));
INV_X1 i_0_672 (.ZN (n_0_343), .A (n_40));
NOR3_X4 i_0_670 (.ZN (n_0_342), .A1 (n_39), .A2 (n_40), .A3 (n_0_312));
OAI221_X1 i_0_669 (.ZN (n_371), .A (n_0_341), .B1 (n_0_338), .B2 (n_0_95), .C1 (n_0_340), .C2 (n_0_92));
OAI21_X1 i_0_667 (.ZN (n_0_341), .A (n_22), .B1 (n_0_336), .B2 (drc_ipo_n32));
OR2_X2 i_0_664 (.ZN (n_0_340), .A1 (n_0_337), .A2 (n_0_268));
OR2_X2 i_0_663 (.ZN (n_0_338), .A1 (n_0_337), .A2 (n_36));
OAI21_X1 i_0_656 (.ZN (n_0_337), .A (n_0_313), .B1 (n_37), .B2 (n_38));
INV_X2 i_0_655 (.ZN (n_0_336), .A (n_0_334));
NAND2_X1 i_0_622 (.ZN (n_0_334), .A1 (n_0_330), .A2 (n_0_268));
INV_X1 i_0_621 (.ZN (n_0_330), .A (n_0_313));
NAND2_X1 i_0_619 (.ZN (n_0_313), .A1 (n_37), .A2 (n_38));
INV_X1 i_0_617 (.ZN (n_0_312), .A (n_38));
NOR3_X1 i_0_616 (.ZN (n_0_311), .A1 (n_37), .A2 (n_38), .A3 (n_0_268));
INV_X1 i_0_615 (.ZN (n_0_310), .A (n_4));
AOI22_X1 i_0_612 (.ZN (n_0_307), .A1 (\A_imm_2s_complement[18] ), .A2 (n_0_280), .B1 (\A_imm_2s_complement[17] ), .B2 (spc__n131));
OAI221_X1 i_0_610 (.ZN (n_370), .A (n_0_307), .B1 (n_0_310), .B2 (n_0_282), .C1 (n_0_361), .C2 (n_0_276));
INV_X1 i_0_609 (.ZN (n_0_306), .A (n_8));
INV_X2 i_0_608 (.ZN (n_0_305), .A (\A_imm_2s_complement[14] ));
AOI22_X1 i_0_603 (.ZN (n_0_304), .A1 (\A_imm_2s_complement[13] ), .A2 (spc__n131)
    , .B1 (n_0_278), .B2 (n_9));
OAI221_X1 i_0_602 (.ZN (n_369), .A (n_0_304), .B1 (n_0_305), .B2 (n_0_281), .C1 (n_0_306), .C2 (n_0_282));
OAI221_X1 i_0_565 (.ZN (n_368), .A (n_0_301), .B1 (n_0_282), .B2 (n_0_95), .C1 (n_0_281), .C2 (n_0_92));
OAI21_X1 i_0_564 (.ZN (n_0_301), .A (n_22), .B1 (n_0_278), .B2 (spc__n131));
OR2_X2 i_0_562 (.ZN (n_0_282), .A1 (n_0_279), .A2 (n_34));
INV_X2 i_0_560 (.ZN (n_0_281), .A (n_0_280));
NOR2_X1 i_0_559 (.ZN (n_0_280), .A1 (n_0_279), .A2 (n_0_219));
OAI21_X1 i_0_558 (.ZN (n_0_279), .A (n_0_274), .B1 (n_35), .B2 (n_36));
INV_X1 i_0_556 (.ZN (n_0_278), .A (n_0_276));
NAND2_X1 i_0_555 (.ZN (n_0_276), .A1 (n_0_275), .A2 (n_0_219));
INV_X1 i_0_553 (.ZN (n_0_275), .A (n_0_274));
NAND2_X1 i_0_542 (.ZN (n_0_274), .A1 (n_35), .A2 (n_36));
INV_X1 i_0_541 (.ZN (n_0_268), .A (n_36));
NOR3_X1 i_0_508 (.ZN (n_0_251), .A1 (n_35), .A2 (n_36), .A3 (n_0_219));
OAI221_X1 i_0_507 (.ZN (n_367), .A (n_0_250), .B1 (n_0_248), .B2 (n_0_95), .C1 (n_0_249), .C2 (n_0_92));
OAI21_X1 i_0_505 (.ZN (n_0_250), .A (n_22), .B1 (n_0_245), .B2 (spc__n134));
OR2_X2 i_0_503 (.ZN (n_0_249), .A1 (n_0_247), .A2 (n_0_188));
OR2_X2 i_0_502 (.ZN (n_0_248), .A1 (n_0_247), .A2 (n_32));
OAI21_X1 i_0_501 (.ZN (n_0_247), .A (n_0_220), .B1 (n_33), .B2 (n_34));
INV_X2 i_0_499 (.ZN (n_0_245), .A (n_0_244));
NAND2_X1 i_0_498 (.ZN (n_0_244), .A1 (n_0_243), .A2 (n_0_188));
INV_X1 i_0_496 (.ZN (n_0_243), .A (n_0_220));
NAND2_X1 i_0_485 (.ZN (n_0_220), .A1 (n_33), .A2 (n_34));
INV_X1 i_0_484 (.ZN (n_0_219), .A (n_34));
NOR3_X4 i_0_451 (.ZN (n_0_218), .A1 (n_33), .A2 (n_34), .A3 (n_0_188));
OAI221_X1 i_0_450 (.ZN (n_366), .A (n_0_217), .B1 (n_0_214), .B2 (n_0_95), .C1 (n_0_216), .C2 (n_0_92));
OAI21_X1 i_0_448 (.ZN (n_0_217), .A (n_22), .B1 (n_0_212), .B2 (drc_ipo_n30));
OR2_X2 i_0_446 (.ZN (n_0_216), .A1 (n_0_213), .A2 (n_0_155));
OR2_X2 i_0_445 (.ZN (n_0_214), .A1 (n_0_213), .A2 (n_30));
OAI21_X1 i_0_444 (.ZN (n_0_213), .A (n_0_189), .B1 (n_31), .B2 (n_32));
INV_X2 i_0_442 (.ZN (n_0_212), .A (n_0_206));
NAND2_X1 i_0_441 (.ZN (n_0_206), .A1 (n_0_202), .A2 (n_0_155));
INV_X1 i_0_439 (.ZN (n_0_202), .A (n_0_189));
NAND2_X1 i_0_428 (.ZN (n_0_189), .A1 (n_31), .A2 (n_32));
INV_X1 i_0_427 (.ZN (n_0_188), .A (n_32));
NOR3_X1 i_0_420 (.ZN (n_0_187), .A1 (n_31), .A2 (n_32), .A3 (n_0_155));
OAI221_X1 i_0_419 (.ZN (n_365), .A (n_0_186), .B1 (n_0_183), .B2 (n_0_95), .C1 (n_0_185), .C2 (n_0_92));
OAI21_X1 i_0_394 (.ZN (n_0_186), .A (n_22), .B1 (n_0_181), .B2 (drc_ipo_n31));
OR2_X2 i_0_393 (.ZN (n_0_185), .A1 (n_0_182), .A2 (n_0_120));
OR2_X2 i_0_391 (.ZN (n_0_183), .A1 (n_0_182), .A2 (n_28));
OAI21_X1 i_0_389 (.ZN (n_0_182), .A (n_0_156), .B1 (n_29), .B2 (n_30));
INV_X2 i_0_388 (.ZN (n_0_181), .A (n_0_158));
NAND2_X1 i_0_387 (.ZN (n_0_158), .A1 (n_0_157), .A2 (n_0_120));
INV_X1 i_0_385 (.ZN (n_0_157), .A (n_0_156));
NAND2_X1 i_0_384 (.ZN (n_0_156), .A1 (n_29), .A2 (n_30));
INV_X1 i_0_382 (.ZN (n_0_155), .A (n_30));
NOR3_X1 i_0_337 (.ZN (n_0_154), .A1 (n_29), .A2 (n_30), .A3 (n_0_120));
OAI221_X1 i_0_336 (.ZN (n_364), .A (n_0_152), .B1 (n_0_151), .B2 (n_0_95), .C1 (n_0_150), .C2 (n_0_92));
OAI21_X1 i_0_334 (.ZN (n_0_152), .A (n_22), .B1 (n_0_125), .B2 (n_0_126));
OR2_X1 i_0_332 (.ZN (n_0_151), .A1 (n_0_127), .A2 (n_26));
OR2_X2 i_0_331 (.ZN (n_0_150), .A1 (n_0_127), .A2 (n_0_63));
OAI21_X1 i_0_330 (.ZN (n_0_127), .A (n_0_121), .B1 (n_27), .B2 (n_28));
NOR3_X4 i_0_328 (.ZN (n_0_126), .A1 (n_27), .A2 (n_28), .A3 (n_0_63));
INV_X2 i_0_327 (.ZN (n_0_125), .A (n_0_124));
NAND2_X1 i_0_325 (.ZN (n_0_124), .A1 (n_0_123), .A2 (n_0_63));
INV_X1 i_0_280 (.ZN (n_0_123), .A (n_0_121));
NAND2_X1 i_0_279 (.ZN (n_0_121), .A1 (n_27), .A2 (n_28));
INV_X1 i_0_277 (.ZN (n_0_120), .A (n_28));
OAI221_X1 i_0_275 (.ZN (n_363), .A (n_0_119), .B1 (n_0_96), .B2 (n_0_95), .C1 (n_0_94), .C2 (n_0_92));
OAI21_X1 i_0_274 (.ZN (n_0_119), .A (n_22), .B1 (n_0_90), .B2 (spc__n136));
OR2_X1 i_0_273 (.ZN (n_0_96), .A1 (n_0_93), .A2 (n_24));
INV_X1 i_0_272 (.ZN (n_0_95), .A (n_21));
OR2_X2 i_0_271 (.ZN (n_0_94), .A1 (n_0_93), .A2 (n_0_33));
OAI21_X1 i_0_270 (.ZN (n_0_93), .A (n_0_64), .B1 (n_25), .B2 (n_26));
INV_X1 i_0_269 (.ZN (n_0_92), .A (\A_imm_2s_complement[1] ));
NOR3_X4 i_0_268 (.ZN (n_0_91), .A1 (n_25), .A2 (n_26), .A3 (n_0_33));
INV_X1 i_0_223 (.ZN (n_0_90), .A (n_0_88));
NAND2_X1 i_0_222 (.ZN (n_0_88), .A1 (n_0_65), .A2 (n_0_33));
INV_X1 i_0_220 (.ZN (n_0_65), .A (n_0_64));
NAND2_X1 i_0_218 (.ZN (n_0_64), .A1 (n_25), .A2 (n_26));
INV_X1 i_0_217 (.ZN (n_0_63), .A (n_26));
OAI222_X1 i_0_216 (.ZN (n_362), .A1 (n_0_62), .A2 (n_0_60), .B1 (n_0_30), .B2 (n_0_27)
    , .C1 (n_0_59), .C2 (n_0_31));
OR2_X1 i_0_215 (.ZN (n_0_62), .A1 (n_0_61), .A2 (n_0_28));
OAI21_X1 i_0_214 (.ZN (n_0_61), .A (n_0_34), .B1 (n_23), .B2 (n_24));
INV_X2 i_0_211 (.ZN (n_0_60), .A (\A_imm_2s_complement[23] ));
NAND2_X1 i_0_166 (.ZN (n_0_59), .A1 (n_0_57), .A2 (n_0_28));
INV_X1 i_0_165 (.ZN (n_0_57), .A (n_0_34));
NAND2_X1 i_0_163 (.ZN (n_0_34), .A1 (n_23), .A2 (n_24));
INV_X1 i_0_162 (.ZN (n_0_33), .A (n_24));
INV_X2 i_0_161 (.ZN (n_0_31), .A (n_0));
INV_X1 i_0_160 (.ZN (n_0_30), .A (n_0_29));
NOR3_X4 i_0_159 (.ZN (n_0_29), .A1 (n_0_28), .A2 (n_23), .A3 (n_24));
INV_X4 i_0_158 (.ZN (n_0_28), .A (n_46));
INV_X8 i_0_157 (.ZN (n_0_27), .A (\A_imm_2s_complement[22] ));
INV_X2 i_0_156 (.ZN (n_0_385), .A (\A_imm_2s_complement[18] ));
INV_X2 i_0_155 (.ZN (n_0_391), .A (\A_imm_2s_complement[27] ));
INV_X2 i_0_721 (.ZN (n_0_388), .A (\A_imm_2s_complement[21] ));
INV_X4 i_0_719 (.ZN (n_0_386), .A (\A_imm_2s_complement[19] ));
INV_X2 i_0_717 (.ZN (n_0_384), .A (\A_imm_2s_complement[17] ));
INV_X2 i_0_716 (.ZN (n_0_383), .A (\A_imm_2s_complement[16] ));
INV_X2 i_0_715 (.ZN (n_0_382), .A (\A_imm_2s_complement[15] ));
INV_X2 i_0_713 (.ZN (n_0_380), .A (\A_imm_2s_complement[13] ));
INV_X1 i_0_712 (.ZN (n_0_379), .A (\A_imm_2s_complement[12] ));
INV_X1 i_0_711 (.ZN (n_0_378), .A (\A_imm_2s_complement[11] ));
INV_X2 i_0_710 (.ZN (n_0_377), .A (\A_imm_2s_complement[10] ));
INV_X2 i_0_709 (.ZN (n_0_376), .A (\A_imm_2s_complement[9] ));
INV_X1 i_0_708 (.ZN (n_0_375), .A (\A_imm_2s_complement[8] ));
INV_X1 i_0_707 (.ZN (n_0_374), .A (\A_imm_2s_complement[7] ));
INV_X2 i_0_706 (.ZN (n_0_373), .A (\A_imm_2s_complement[6] ));
INV_X2 i_0_705 (.ZN (n_0_372), .A (\A_imm_2s_complement[5] ));
INV_X1 i_0_704 (.ZN (n_0_371), .A (\A_imm_2s_complement[4] ));
INV_X1 i_0_703 (.ZN (n_0_370), .A (\A_imm_2s_complement[3] ));
INV_X1 i_0_154 (.ZN (n_0_369), .A (\A_imm_2s_complement[2] ));
INV_X1 i_0_698 (.ZN (n_0_365), .A (n_1));
INV_X1 i_0_696 (.ZN (n_0_363), .A (n_3));
INV_X2 i_0_694 (.ZN (n_0_361), .A (n_5));
INV_X1 i_0_693 (.ZN (n_0_360), .A (n_6));
INV_X1 i_0_692 (.ZN (n_0_359), .A (n_7));
INV_X1 i_0_690 (.ZN (n_0_357), .A (n_9));
INV_X1 i_0_689 (.ZN (n_0_356), .A (n_10));
INV_X1 i_0_688 (.ZN (n_0_355), .A (n_11));
INV_X1 i_0_687 (.ZN (n_0_354), .A (n_12));
INV_X1 i_0_686 (.ZN (n_0_353), .A (n_13));
INV_X1 i_0_685 (.ZN (n_0_352), .A (n_14));
INV_X1 i_0_684 (.ZN (n_0_351), .A (n_15));
INV_X1 i_0_683 (.ZN (n_0_350), .A (n_16));
INV_X1 i_0_682 (.ZN (n_0_349), .A (n_17));
INV_X1 i_0_681 (.ZN (n_0_348), .A (n_18));
INV_X1 i_0_680 (.ZN (n_0_347), .A (n_19));
INV_X1 i_0_151 (.ZN (n_0_346), .A (n_20));
INV_X1 i_0_150 (.ZN (n_0_344), .A (n_22));
NOR3_X1 i_0_675 (.ZN (n_361), .A1 (n_0_392), .A2 (n_0_391), .A3 (n_0_409));
INV_X1 i_0_671 (.ZN (n_0_339), .A (n_0_406));
OAI222_X1 i_0_668 (.ZN (n_360), .A1 (n_0_60), .A2 (n_0_339), .B1 (n_0_28), .B2 (n_0_410)
    , .C1 (n_0_391), .C2 (n_0_414));
AOI22_X1 i_0_666 (.ZN (n_0_335), .A1 (n_0), .A2 (n_0_411), .B1 (\A_imm_2s_complement[22] ), .B2 (n_0_406));
OAI221_X1 i_0_665 (.ZN (n_359), .A (n_0_335), .B1 (n_0_28), .B2 (n_0_415), .C1 (n_0_60), .C2 (n_0_414));
AOI22_X1 i_0_662 (.ZN (n_0_333), .A1 (n_2), .A2 (n_0_411), .B1 (\A_imm_2s_complement[20] ), .B2 (n_0_406));
OAI221_X1 i_0_661 (.ZN (n_358), .A (n_0_333), .B1 (n_0_365), .B2 (n_0_415), .C1 (n_0_388), .C2 (n_0_414));
AOI22_X1 i_0_660 (.ZN (n_0_332), .A1 (n_3), .A2 (n_0_411), .B1 (\A_imm_2s_complement[19] ), .B2 (n_0_406));
OAI221_X1 i_0_659 (.ZN (n_357), .A (n_0_332), .B1 (n_0_404), .B2 (n_0_415), .C1 (n_0_403), .C2 (n_0_414));
AOI22_X1 i_0_658 (.ZN (n_0_331), .A1 (n_4), .A2 (n_0_411), .B1 (\A_imm_2s_complement[18] ), .B2 (n_0_406));
OAI221_X1 i_0_657 (.ZN (n_356), .A (n_0_331), .B1 (n_0_363), .B2 (n_0_415), .C1 (n_0_386), .C2 (n_0_414));
AOI22_X1 i_0_654 (.ZN (n_0_329), .A1 (n_6), .A2 (n_0_411), .B1 (\A_imm_2s_complement[16] ), .B2 (n_0_406));
OAI221_X1 i_0_653 (.ZN (n_355), .A (n_0_329), .B1 (n_0_361), .B2 (n_0_415), .C1 (n_0_384), .C2 (n_0_414));
AOI22_X1 i_0_652 (.ZN (n_0_328), .A1 (n_7), .A2 (n_0_411), .B1 (\A_imm_2s_complement[15] ), .B2 (n_0_406));
OAI221_X1 i_0_651 (.ZN (n_354), .A (n_0_328), .B1 (n_0_360), .B2 (n_0_415), .C1 (n_0_383), .C2 (n_0_414));
AOI22_X1 i_0_650 (.ZN (n_0_327), .A1 (n_8), .A2 (n_0_411), .B1 (\A_imm_2s_complement[14] ), .B2 (n_0_406));
OAI221_X1 i_0_649 (.ZN (n_353), .A (n_0_327), .B1 (n_0_359), .B2 (n_0_415), .C1 (n_0_382), .C2 (n_0_414));
AOI22_X1 i_0_648 (.ZN (n_0_326), .A1 (n_9), .A2 (n_0_411), .B1 (\A_imm_2s_complement[13] ), .B2 (n_0_406));
OAI221_X1 i_0_647 (.ZN (n_352), .A (n_0_326), .B1 (n_0_306), .B2 (n_0_415), .C1 (n_0_305), .C2 (n_0_414));
AOI22_X1 i_0_646 (.ZN (n_0_325), .A1 (n_10), .A2 (n_0_411), .B1 (\A_imm_2s_complement[12] ), .B2 (n_0_406));
OAI221_X1 i_0_645 (.ZN (n_351), .A (n_0_325), .B1 (n_0_357), .B2 (n_0_415), .C1 (n_0_380), .C2 (n_0_414));
AOI22_X1 i_0_644 (.ZN (n_0_324), .A1 (n_11), .A2 (n_0_411), .B1 (\A_imm_2s_complement[11] ), .B2 (n_0_406));
OAI221_X1 i_0_643 (.ZN (n_350), .A (n_0_324), .B1 (n_0_356), .B2 (n_0_415), .C1 (n_0_379), .C2 (n_0_414));
AOI22_X1 i_0_642 (.ZN (n_0_323), .A1 (n_12), .A2 (n_0_411), .B1 (\A_imm_2s_complement[10] ), .B2 (n_0_406));
OAI221_X1 i_0_641 (.ZN (n_349), .A (n_0_323), .B1 (n_0_355), .B2 (n_0_415), .C1 (n_0_378), .C2 (n_0_414));
AOI22_X1 i_0_640 (.ZN (n_0_322), .A1 (n_13), .A2 (n_0_411), .B1 (\A_imm_2s_complement[9] ), .B2 (n_0_406));
OAI221_X1 i_0_639 (.ZN (n_348), .A (n_0_322), .B1 (n_0_354), .B2 (n_0_415), .C1 (n_0_377), .C2 (n_0_414));
AOI22_X1 i_0_638 (.ZN (n_0_321), .A1 (n_14), .A2 (n_0_411), .B1 (\A_imm_2s_complement[8] ), .B2 (n_0_406));
OAI221_X1 i_0_637 (.ZN (n_347), .A (n_0_321), .B1 (n_0_353), .B2 (n_0_415), .C1 (n_0_376), .C2 (n_0_414));
AOI22_X1 i_0_636 (.ZN (n_0_320), .A1 (n_15), .A2 (n_0_411), .B1 (\A_imm_2s_complement[7] ), .B2 (n_0_406));
OAI221_X1 i_0_635 (.ZN (n_346), .A (n_0_320), .B1 (n_0_352), .B2 (n_0_415), .C1 (n_0_375), .C2 (n_0_414));
AOI22_X1 i_0_634 (.ZN (n_0_319), .A1 (n_16), .A2 (n_0_411), .B1 (\A_imm_2s_complement[6] ), .B2 (n_0_406));
OAI221_X1 i_0_633 (.ZN (n_345), .A (n_0_319), .B1 (n_0_351), .B2 (n_0_415), .C1 (n_0_374), .C2 (n_0_414));
AOI22_X1 i_0_632 (.ZN (n_0_318), .A1 (n_17), .A2 (n_0_411), .B1 (\A_imm_2s_complement[5] ), .B2 (n_0_406));
OAI221_X1 i_0_631 (.ZN (n_344), .A (n_0_318), .B1 (n_0_350), .B2 (n_0_415), .C1 (n_0_373), .C2 (n_0_414));
AOI22_X1 i_0_630 (.ZN (n_0_317), .A1 (n_18), .A2 (n_0_411), .B1 (\A_imm_2s_complement[4] ), .B2 (n_0_406));
OAI221_X1 i_0_629 (.ZN (n_343), .A (n_0_317), .B1 (n_0_349), .B2 (n_0_415), .C1 (n_0_372), .C2 (n_0_414));
AOI22_X1 i_0_628 (.ZN (n_0_316), .A1 (n_19), .A2 (n_0_411), .B1 (\A_imm_2s_complement[3] ), .B2 (n_0_406));
OAI221_X1 i_0_627 (.ZN (n_342), .A (n_0_316), .B1 (n_0_348), .B2 (n_0_415), .C1 (n_0_371), .C2 (n_0_414));
AOI22_X1 i_0_626 (.ZN (n_0_315), .A1 (n_20), .A2 (n_0_411), .B1 (\A_imm_2s_complement[2] ), .B2 (n_0_406));
OAI221_X1 i_0_625 (.ZN (n_341), .A (n_0_315), .B1 (n_0_347), .B2 (n_0_415), .C1 (n_0_370), .C2 (n_0_414));
AOI22_X1 i_0_624 (.ZN (n_0_314), .A1 (n_21), .A2 (n_0_411), .B1 (\A_imm_2s_complement[1] ), .B2 (n_0_406));
OAI221_X1 i_0_623 (.ZN (n_340), .A (n_0_314), .B1 (n_0_346), .B2 (n_0_415), .C1 (n_0_369), .C2 (n_0_414));
NOR2_X1 i_0_620 (.ZN (n_339), .A1 (n_0_344), .A2 (n_0_412));
NOR3_X1 i_0_618 (.ZN (n_338), .A1 (n_0_343), .A2 (n_0_391), .A3 (n_0_394));
INV_X1 i_0_614 (.ZN (n_0_308), .A (n_0_390));
OAI222_X1 i_0_611 (.ZN (n_337), .A1 (n_0_60), .A2 (n_0_308), .B1 (n_0_28), .B2 (n_0_395)
    , .C1 (n_0_391), .C2 (n_0_399));
AOI22_X1 i_0_607 (.ZN (n_0_303), .A1 (n_1), .A2 (n_0_396), .B1 (\A_imm_2s_complement[21] ), .B2 (n_0_390));
OAI221_X1 i_0_606 (.ZN (n_336), .A (n_0_303), .B1 (n_0_31), .B2 (n_0_400), .C1 (n_0_27), .C2 (n_0_399));
AOI22_X1 i_0_605 (.ZN (n_0_302), .A1 (n_2), .A2 (n_0_396), .B1 (\A_imm_2s_complement[20] ), .B2 (n_0_390));
OAI221_X1 i_0_604 (.ZN (n_335), .A (n_0_302), .B1 (n_0_365), .B2 (n_0_400), .C1 (n_0_388), .C2 (n_0_399));
AOI22_X1 i_0_601 (.ZN (n_0_300), .A1 (n_4), .A2 (n_0_396), .B1 (\A_imm_2s_complement[18] ), .B2 (n_0_390));
OAI221_X1 i_0_600 (.ZN (n_334), .A (n_0_300), .B1 (n_0_363), .B2 (n_0_400), .C1 (n_0_386), .C2 (n_0_399));
AOI22_X1 i_0_599 (.ZN (n_0_299), .A1 (n_5), .A2 (n_0_396), .B1 (\A_imm_2s_complement[17] ), .B2 (n_0_390));
OAI221_X1 i_0_598 (.ZN (n_333), .A (n_0_299), .B1 (n_0_310), .B2 (n_0_400), .C1 (n_0_385), .C2 (n_0_399));
AOI22_X1 i_0_597 (.ZN (n_0_298), .A1 (n_6), .A2 (n_0_396), .B1 (\A_imm_2s_complement[16] ), .B2 (n_0_390));
OAI221_X1 i_0_596 (.ZN (n_332), .A (n_0_298), .B1 (n_0_361), .B2 (n_0_400), .C1 (n_0_384), .C2 (n_0_399));
AOI22_X1 i_0_595 (.ZN (n_0_297), .A1 (n_7), .A2 (n_0_396), .B1 (\A_imm_2s_complement[15] ), .B2 (n_0_390));
OAI221_X1 i_0_594 (.ZN (n_331), .A (n_0_297), .B1 (n_0_360), .B2 (n_0_400), .C1 (n_0_383), .C2 (n_0_399));
AOI22_X1 i_0_593 (.ZN (n_0_296), .A1 (n_8), .A2 (n_0_396), .B1 (\A_imm_2s_complement[14] ), .B2 (n_0_390));
OAI221_X1 i_0_592 (.ZN (n_330), .A (n_0_296), .B1 (n_0_359), .B2 (n_0_400), .C1 (n_0_382), .C2 (n_0_399));
AOI22_X1 i_0_591 (.ZN (n_0_295), .A1 (n_9), .A2 (n_0_396), .B1 (\A_imm_2s_complement[13] ), .B2 (n_0_390));
OAI221_X1 i_0_590 (.ZN (n_329), .A (n_0_295), .B1 (n_0_306), .B2 (n_0_400), .C1 (n_0_305), .C2 (n_0_399));
AOI22_X1 i_0_589 (.ZN (n_0_294), .A1 (n_10), .A2 (n_0_396), .B1 (\A_imm_2s_complement[12] ), .B2 (n_0_390));
OAI221_X1 i_0_588 (.ZN (n_328), .A (n_0_294), .B1 (n_0_357), .B2 (n_0_400), .C1 (n_0_380), .C2 (n_0_399));
AOI22_X1 i_0_587 (.ZN (n_0_293), .A1 (n_11), .A2 (n_0_396), .B1 (\A_imm_2s_complement[11] ), .B2 (n_0_390));
OAI221_X1 i_0_586 (.ZN (n_327), .A (n_0_293), .B1 (n_0_356), .B2 (n_0_400), .C1 (n_0_379), .C2 (n_0_399));
AOI22_X1 i_0_585 (.ZN (n_0_292), .A1 (n_12), .A2 (n_0_396), .B1 (\A_imm_2s_complement[10] ), .B2 (n_0_390));
OAI221_X1 i_0_584 (.ZN (n_326), .A (n_0_292), .B1 (n_0_355), .B2 (n_0_400), .C1 (n_0_378), .C2 (n_0_399));
AOI22_X1 i_0_583 (.ZN (n_0_291), .A1 (n_13), .A2 (n_0_396), .B1 (\A_imm_2s_complement[9] ), .B2 (n_0_390));
OAI221_X1 i_0_582 (.ZN (n_325), .A (n_0_291), .B1 (n_0_354), .B2 (n_0_400), .C1 (n_0_377), .C2 (n_0_399));
AOI22_X1 i_0_581 (.ZN (n_0_290), .A1 (n_14), .A2 (n_0_396), .B1 (\A_imm_2s_complement[8] ), .B2 (n_0_390));
OAI221_X1 i_0_580 (.ZN (n_324), .A (n_0_290), .B1 (n_0_353), .B2 (n_0_400), .C1 (n_0_376), .C2 (n_0_399));
AOI22_X1 i_0_579 (.ZN (n_0_289), .A1 (n_15), .A2 (n_0_396), .B1 (\A_imm_2s_complement[7] ), .B2 (n_0_390));
OAI221_X1 i_0_578 (.ZN (n_323), .A (n_0_289), .B1 (n_0_352), .B2 (n_0_400), .C1 (n_0_375), .C2 (n_0_399));
AOI22_X1 i_0_577 (.ZN (n_0_288), .A1 (n_16), .A2 (n_0_396), .B1 (\A_imm_2s_complement[6] ), .B2 (n_0_390));
OAI221_X1 i_0_576 (.ZN (n_322), .A (n_0_288), .B1 (n_0_351), .B2 (n_0_400), .C1 (n_0_374), .C2 (n_0_399));
AOI22_X1 i_0_575 (.ZN (n_0_287), .A1 (n_17), .A2 (n_0_396), .B1 (\A_imm_2s_complement[5] ), .B2 (n_0_390));
OAI221_X1 i_0_574 (.ZN (n_321), .A (n_0_287), .B1 (n_0_350), .B2 (n_0_400), .C1 (n_0_373), .C2 (n_0_399));
AOI22_X1 i_0_573 (.ZN (n_0_286), .A1 (n_18), .A2 (n_0_396), .B1 (\A_imm_2s_complement[4] ), .B2 (n_0_390));
OAI221_X1 i_0_572 (.ZN (n_320), .A (n_0_286), .B1 (n_0_349), .B2 (n_0_400), .C1 (n_0_372), .C2 (n_0_399));
AOI22_X1 i_0_571 (.ZN (n_0_285), .A1 (n_19), .A2 (n_0_396), .B1 (\A_imm_2s_complement[3] ), .B2 (n_0_390));
OAI221_X1 i_0_570 (.ZN (n_319), .A (n_0_285), .B1 (n_0_348), .B2 (n_0_400), .C1 (n_0_371), .C2 (n_0_399));
AOI22_X1 i_0_569 (.ZN (n_0_284), .A1 (n_20), .A2 (n_0_396), .B1 (\A_imm_2s_complement[2] ), .B2 (n_0_390));
OAI221_X1 i_0_568 (.ZN (n_318), .A (n_0_284), .B1 (n_0_347), .B2 (n_0_400), .C1 (n_0_370), .C2 (n_0_399));
AOI22_X1 i_0_567 (.ZN (n_0_283), .A1 (n_21), .A2 (n_0_396), .B1 (\A_imm_2s_complement[1] ), .B2 (n_0_390));
OAI221_X1 i_0_566 (.ZN (n_317), .A (n_0_283), .B1 (n_0_346), .B2 (n_0_400), .C1 (n_0_369), .C2 (n_0_399));
NOR2_X1 i_0_563 (.ZN (n_316), .A1 (n_0_344), .A2 (n_0_397));
NOR3_X1 i_0_561 (.ZN (n_315), .A1 (n_0_312), .A2 (n_0_391), .A3 (n_0_358));
INV_X1 i_0_557 (.ZN (n_0_277), .A (n_0_342));
OAI222_X1 i_0_554 (.ZN (n_314), .A1 (n_0_60), .A2 (n_0_277), .B1 (n_0_28), .B2 (n_0_362)
    , .C1 (n_0_391), .C2 (n_0_368));
AOI22_X1 i_0_552 (.ZN (n_0_273), .A1 (n_0), .A2 (n_0_364), .B1 (\A_imm_2s_complement[22] ), .B2 (n_0_342));
OAI221_X1 i_0_551 (.ZN (n_313), .A (n_0_273), .B1 (n_0_28), .B2 (n_0_381), .C1 (n_0_60), .C2 (n_0_368));
AOI22_X1 i_0_550 (.ZN (n_0_272), .A1 (n_1), .A2 (n_0_364), .B1 (\A_imm_2s_complement[21] ), .B2 (n_0_342));
OAI221_X1 i_0_549 (.ZN (n_312), .A (n_0_272), .B1 (n_0_31), .B2 (n_0_381), .C1 (n_0_27), .C2 (n_0_368));
AOI22_X1 i_0_548 (.ZN (n_0_271), .A1 (n_2), .A2 (n_0_364), .B1 (\A_imm_2s_complement[20] ), .B2 (n_0_342));
OAI221_X1 i_0_547 (.ZN (n_311), .A (n_0_271), .B1 (n_0_365), .B2 (n_0_381), .C1 (n_0_388), .C2 (n_0_368));
AOI22_X1 i_0_546 (.ZN (n_0_270), .A1 (n_3), .A2 (n_0_364), .B1 (\A_imm_2s_complement[19] ), .B2 (n_0_342));
OAI221_X1 i_0_545 (.ZN (n_310), .A (n_0_270), .B1 (n_0_404), .B2 (n_0_381), .C1 (n_0_403), .C2 (n_0_368));
AOI22_X1 i_0_544 (.ZN (n_0_269), .A1 (n_4), .A2 (n_0_364), .B1 (\A_imm_2s_complement[18] ), .B2 (n_0_342));
OAI221_X1 i_0_543 (.ZN (n_309), .A (n_0_269), .B1 (n_0_363), .B2 (n_0_381), .C1 (n_0_386), .C2 (n_0_368));
AOI22_X1 i_0_540 (.ZN (n_0_267), .A1 (n_6), .A2 (n_0_364), .B1 (\A_imm_2s_complement[16] ), .B2 (n_0_342));
OAI221_X1 i_0_539 (.ZN (n_308), .A (n_0_267), .B1 (n_0_361), .B2 (n_0_381), .C1 (n_0_384), .C2 (n_0_368));
AOI22_X1 i_0_538 (.ZN (n_0_266), .A1 (n_7), .A2 (n_0_364), .B1 (\A_imm_2s_complement[15] ), .B2 (n_0_342));
OAI221_X1 i_0_537 (.ZN (n_307), .A (n_0_266), .B1 (n_0_360), .B2 (n_0_381), .C1 (n_0_383), .C2 (n_0_368));
AOI22_X1 i_0_536 (.ZN (n_0_265), .A1 (n_8), .A2 (n_0_364), .B1 (\A_imm_2s_complement[14] ), .B2 (n_0_342));
OAI221_X1 i_0_535 (.ZN (n_306), .A (n_0_265), .B1 (n_0_359), .B2 (n_0_381), .C1 (n_0_382), .C2 (n_0_368));
AOI22_X1 i_0_534 (.ZN (n_0_264), .A1 (n_9), .A2 (n_0_364), .B1 (\A_imm_2s_complement[13] ), .B2 (n_0_342));
OAI221_X1 i_0_533 (.ZN (n_305), .A (n_0_264), .B1 (n_0_306), .B2 (n_0_381), .C1 (n_0_305), .C2 (n_0_368));
AOI22_X1 i_0_532 (.ZN (n_0_263), .A1 (n_10), .A2 (n_0_364), .B1 (\A_imm_2s_complement[12] ), .B2 (n_0_342));
OAI221_X1 i_0_531 (.ZN (n_304), .A (n_0_263), .B1 (n_0_357), .B2 (n_0_381), .C1 (n_0_380), .C2 (n_0_368));
AOI22_X1 i_0_530 (.ZN (n_0_262), .A1 (n_11), .A2 (n_0_364), .B1 (\A_imm_2s_complement[11] ), .B2 (n_0_342));
OAI221_X1 i_0_529 (.ZN (n_303), .A (n_0_262), .B1 (n_0_356), .B2 (n_0_381), .C1 (n_0_379), .C2 (n_0_368));
AOI22_X1 i_0_528 (.ZN (n_0_261), .A1 (n_12), .A2 (n_0_364), .B1 (\A_imm_2s_complement[10] ), .B2 (n_0_342));
OAI221_X1 i_0_527 (.ZN (n_302), .A (n_0_261), .B1 (n_0_355), .B2 (n_0_381), .C1 (n_0_378), .C2 (n_0_368));
AOI22_X1 i_0_526 (.ZN (n_0_260), .A1 (n_13), .A2 (n_0_364), .B1 (\A_imm_2s_complement[9] ), .B2 (n_0_342));
OAI221_X1 i_0_525 (.ZN (n_301), .A (n_0_260), .B1 (n_0_354), .B2 (n_0_381), .C1 (n_0_377), .C2 (n_0_368));
AOI22_X1 i_0_524 (.ZN (n_0_259), .A1 (n_14), .A2 (n_0_364), .B1 (\A_imm_2s_complement[8] ), .B2 (n_0_342));
OAI221_X1 i_0_523 (.ZN (n_300), .A (n_0_259), .B1 (n_0_353), .B2 (n_0_381), .C1 (n_0_376), .C2 (n_0_368));
AOI22_X1 i_0_522 (.ZN (n_0_258), .A1 (n_15), .A2 (n_0_364), .B1 (\A_imm_2s_complement[7] ), .B2 (n_0_342));
OAI221_X1 i_0_521 (.ZN (n_299), .A (n_0_258), .B1 (n_0_352), .B2 (n_0_381), .C1 (n_0_375), .C2 (n_0_368));
AOI22_X1 i_0_520 (.ZN (n_0_257), .A1 (n_16), .A2 (n_0_364), .B1 (\A_imm_2s_complement[6] ), .B2 (n_0_342));
OAI221_X1 i_0_519 (.ZN (n_298), .A (n_0_257), .B1 (n_0_351), .B2 (n_0_381), .C1 (n_0_374), .C2 (n_0_368));
AOI22_X1 i_0_518 (.ZN (n_0_256), .A1 (n_17), .A2 (n_0_364), .B1 (\A_imm_2s_complement[5] ), .B2 (n_0_342));
OAI221_X1 i_0_517 (.ZN (n_297), .A (n_0_256), .B1 (n_0_350), .B2 (n_0_381), .C1 (n_0_373), .C2 (n_0_368));
AOI22_X1 i_0_516 (.ZN (n_0_255), .A1 (n_18), .A2 (n_0_364), .B1 (\A_imm_2s_complement[4] ), .B2 (n_0_342));
OAI221_X1 i_0_515 (.ZN (n_296), .A (n_0_255), .B1 (n_0_349), .B2 (n_0_381), .C1 (n_0_372), .C2 (n_0_368));
AOI22_X1 i_0_514 (.ZN (n_0_254), .A1 (n_19), .A2 (n_0_364), .B1 (\A_imm_2s_complement[3] ), .B2 (n_0_342));
OAI221_X1 i_0_513 (.ZN (n_295), .A (n_0_254), .B1 (n_0_348), .B2 (n_0_381), .C1 (n_0_371), .C2 (n_0_368));
AOI22_X1 i_0_512 (.ZN (n_0_253), .A1 (n_20), .A2 (n_0_364), .B1 (\A_imm_2s_complement[2] ), .B2 (n_0_342));
OAI221_X1 i_0_511 (.ZN (n_294), .A (n_0_253), .B1 (n_0_347), .B2 (n_0_381), .C1 (n_0_370), .C2 (n_0_368));
AOI22_X1 i_0_510 (.ZN (n_0_252), .A1 (n_21), .A2 (n_0_364), .B1 (\A_imm_2s_complement[1] ), .B2 (n_0_342));
OAI221_X1 i_0_509 (.ZN (n_293), .A (n_0_252), .B1 (n_0_346), .B2 (n_0_381), .C1 (n_0_369), .C2 (n_0_368));
NOR2_X1 i_0_506 (.ZN (n_292), .A1 (n_0_344), .A2 (n_0_366));
NOR3_X1 i_0_504 (.ZN (n_291), .A1 (n_0_268), .A2 (n_0_391), .A3 (n_0_330));
INV_X1 i_0_500 (.ZN (n_0_246), .A (drc_ipo_n32));
OAI222_X1 i_0_497 (.ZN (n_290), .A1 (n_0_60), .A2 (n_0_246), .B1 (n_0_28), .B2 (n_0_334)
    , .C1 (n_0_391), .C2 (n_0_340));
AOI22_X1 i_0_495 (.ZN (n_0_242), .A1 (n_0), .A2 (n_0_336), .B1 (\A_imm_2s_complement[22] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_494 (.ZN (n_289), .A (n_0_242), .B1 (n_0_28), .B2 (n_0_338), .C1 (n_0_60), .C2 (n_0_340));
AOI22_X1 i_0_493 (.ZN (n_0_241), .A1 (n_1), .A2 (n_0_336), .B1 (\A_imm_2s_complement[21] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_492 (.ZN (n_288), .A (n_0_241), .B1 (n_0_31), .B2 (n_0_338), .C1 (n_0_27), .C2 (n_0_340));
AOI22_X1 i_0_491 (.ZN (n_0_240), .A1 (n_2), .A2 (n_0_336), .B1 (\A_imm_2s_complement[20] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_490 (.ZN (n_287), .A (n_0_240), .B1 (n_0_365), .B2 (n_0_338), .C1 (n_0_388), .C2 (n_0_340));
AOI22_X1 i_0_489 (.ZN (n_0_239), .A1 (n_3), .A2 (n_0_336), .B1 (\A_imm_2s_complement[19] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_488 (.ZN (n_286), .A (n_0_239), .B1 (n_0_404), .B2 (n_0_338), .C1 (n_0_403), .C2 (n_0_340));
AOI22_X1 i_0_487 (.ZN (n_0_238), .A1 (n_4), .A2 (n_0_336), .B1 (\A_imm_2s_complement[18] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_486 (.ZN (n_285), .A (n_0_238), .B1 (n_0_363), .B2 (n_0_338), .C1 (n_0_386), .C2 (n_0_340));
AOI22_X1 i_0_111 (.ZN (n_0_237), .A1 (n_5), .A2 (n_0_336), .B1 (\A_imm_2s_complement[17] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_110 (.ZN (n_284), .A (n_0_237), .B1 (n_0_310), .B2 (n_0_338), .C1 (n_0_385), .C2 (n_0_340));
AOI22_X1 i_0_483 (.ZN (n_0_236), .A1 (n_6), .A2 (n_0_336), .B1 (\A_imm_2s_complement[16] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_482 (.ZN (n_283), .A (n_0_236), .B1 (n_0_361), .B2 (n_0_338), .C1 (n_0_384), .C2 (n_0_340));
AOI22_X1 i_0_481 (.ZN (n_0_235), .A1 (n_7), .A2 (n_0_336), .B1 (\A_imm_2s_complement[15] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_480 (.ZN (n_282), .A (n_0_235), .B1 (n_0_360), .B2 (n_0_338), .C1 (n_0_383), .C2 (n_0_340));
AOI22_X1 i_0_479 (.ZN (n_0_234), .A1 (n_8), .A2 (n_0_336), .B1 (\A_imm_2s_complement[14] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_478 (.ZN (n_281), .A (n_0_234), .B1 (n_0_359), .B2 (n_0_338), .C1 (n_0_382), .C2 (n_0_340));
AOI22_X1 i_0_477 (.ZN (n_0_233), .A1 (n_9), .A2 (n_0_336), .B1 (\A_imm_2s_complement[13] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_476 (.ZN (n_280), .A (n_0_233), .B1 (n_0_306), .B2 (n_0_338), .C1 (n_0_305), .C2 (n_0_340));
AOI22_X1 i_0_475 (.ZN (n_0_232), .A1 (n_10), .A2 (n_0_336), .B1 (\A_imm_2s_complement[12] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_474 (.ZN (n_279), .A (n_0_232), .B1 (n_0_357), .B2 (n_0_338), .C1 (n_0_380), .C2 (n_0_340));
AOI22_X1 i_0_473 (.ZN (n_0_231), .A1 (n_11), .A2 (n_0_336), .B1 (\A_imm_2s_complement[11] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_472 (.ZN (n_278), .A (n_0_231), .B1 (n_0_356), .B2 (n_0_338), .C1 (n_0_379), .C2 (n_0_340));
AOI22_X1 i_0_471 (.ZN (n_0_230), .A1 (n_12), .A2 (n_0_336), .B1 (\A_imm_2s_complement[10] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_470 (.ZN (n_277), .A (n_0_230), .B1 (n_0_355), .B2 (n_0_338), .C1 (n_0_378), .C2 (n_0_340));
AOI22_X1 i_0_469 (.ZN (n_0_229), .A1 (n_13), .A2 (n_0_336), .B1 (\A_imm_2s_complement[9] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_468 (.ZN (n_276), .A (n_0_229), .B1 (n_0_354), .B2 (n_0_338), .C1 (n_0_377), .C2 (n_0_340));
AOI22_X1 i_0_467 (.ZN (n_0_228), .A1 (n_14), .A2 (n_0_336), .B1 (\A_imm_2s_complement[8] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_466 (.ZN (n_275), .A (n_0_228), .B1 (n_0_353), .B2 (n_0_338), .C1 (n_0_376), .C2 (n_0_340));
AOI22_X1 i_0_465 (.ZN (n_0_227), .A1 (n_15), .A2 (n_0_336), .B1 (\A_imm_2s_complement[7] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_464 (.ZN (n_274), .A (n_0_227), .B1 (n_0_352), .B2 (n_0_338), .C1 (n_0_375), .C2 (n_0_340));
AOI22_X1 i_0_463 (.ZN (n_0_226), .A1 (n_16), .A2 (n_0_336), .B1 (\A_imm_2s_complement[6] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_462 (.ZN (n_273), .A (n_0_226), .B1 (n_0_351), .B2 (n_0_338), .C1 (n_0_374), .C2 (n_0_340));
AOI22_X1 i_0_461 (.ZN (n_0_225), .A1 (n_17), .A2 (n_0_336), .B1 (\A_imm_2s_complement[5] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_460 (.ZN (n_272), .A (n_0_225), .B1 (n_0_350), .B2 (n_0_338), .C1 (n_0_373), .C2 (n_0_340));
AOI22_X1 i_0_459 (.ZN (n_0_224), .A1 (n_18), .A2 (n_0_336), .B1 (\A_imm_2s_complement[4] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_458 (.ZN (n_271), .A (n_0_224), .B1 (n_0_349), .B2 (n_0_338), .C1 (n_0_372), .C2 (n_0_340));
AOI22_X1 i_0_457 (.ZN (n_0_223), .A1 (n_19), .A2 (n_0_336), .B1 (\A_imm_2s_complement[3] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_456 (.ZN (n_270), .A (n_0_223), .B1 (n_0_348), .B2 (n_0_338), .C1 (n_0_371), .C2 (n_0_340));
AOI22_X1 i_0_455 (.ZN (n_0_222), .A1 (n_20), .A2 (n_0_336), .B1 (\A_imm_2s_complement[2] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_454 (.ZN (n_269), .A (n_0_222), .B1 (n_0_347), .B2 (n_0_338), .C1 (n_0_370), .C2 (n_0_340));
AOI22_X1 i_0_453 (.ZN (n_0_221), .A1 (n_21), .A2 (n_0_336), .B1 (\A_imm_2s_complement[1] ), .B2 (drc_ipo_n32));
OAI221_X1 i_0_452 (.ZN (n_268), .A (n_0_221), .B1 (n_0_346), .B2 (n_0_338), .C1 (n_0_369), .C2 (n_0_340));
NOR2_X1 i_0_449 (.ZN (n_267), .A1 (n_0_344), .A2 (n_0_337));
NOR3_X1 i_0_447 (.ZN (n_266), .A1 (n_0_219), .A2 (n_0_391), .A3 (n_0_275));
INV_X1 i_0_443 (.ZN (n_0_215), .A (spc__n131));
OAI222_X1 i_0_440 (.ZN (n_265), .A1 (n_0_60), .A2 (n_0_215), .B1 (n_0_28), .B2 (n_0_276)
    , .C1 (n_0_391), .C2 (n_0_281));
AOI22_X1 i_0_438 (.ZN (n_0_211), .A1 (n_0), .A2 (n_0_278), .B1 (\A_imm_2s_complement[22] ), .B2 (spc__n131));
OAI221_X1 i_0_437 (.ZN (n_264), .A (n_0_211), .B1 (n_0_28), .B2 (n_0_282), .C1 (n_0_60), .C2 (n_0_281));
AOI22_X1 i_0_436 (.ZN (n_0_210), .A1 (n_1), .A2 (n_0_278), .B1 (\A_imm_2s_complement[21] ), .B2 (spc__n131));
OAI221_X1 i_0_435 (.ZN (n_263), .A (n_0_210), .B1 (n_0_31), .B2 (n_0_282), .C1 (n_0_27), .C2 (n_0_281));
AOI22_X1 i_0_434 (.ZN (n_0_209), .A1 (n_2), .A2 (n_0_278), .B1 (\A_imm_2s_complement[20] ), .B2 (spc__n131));
OAI221_X1 i_0_433 (.ZN (n_262), .A (n_0_209), .B1 (n_0_365), .B2 (n_0_282), .C1 (n_0_388), .C2 (n_0_281));
AOI22_X1 i_0_432 (.ZN (n_0_208), .A1 (n_3), .A2 (n_0_278), .B1 (\A_imm_2s_complement[19] ), .B2 (spc__n131));
OAI221_X1 i_0_431 (.ZN (n_261), .A (n_0_208), .B1 (n_0_404), .B2 (n_0_282), .C1 (n_0_403), .C2 (n_0_281));
AOI22_X1 i_0_430 (.ZN (n_0_207), .A1 (n_4), .A2 (n_0_278), .B1 (\A_imm_2s_complement[18] ), .B2 (spc__n131));
OAI221_X1 i_0_429 (.ZN (n_260), .A (n_0_207), .B1 (n_0_363), .B2 (n_0_282), .C1 (n_0_386), .C2 (n_0_281));
AOI22_X1 i_0_426 (.ZN (n_0_205), .A1 (n_6), .A2 (n_0_278), .B1 (\A_imm_2s_complement[16] ), .B2 (spc__n131));
OAI221_X1 i_0_425 (.ZN (n_259), .A (n_0_205), .B1 (n_0_361), .B2 (n_0_282), .C1 (n_0_384), .C2 (n_0_281));
AOI22_X1 i_0_424 (.ZN (n_0_204), .A1 (n_7), .A2 (n_0_278), .B1 (\A_imm_2s_complement[15] ), .B2 (spc__n131));
OAI221_X1 i_0_423 (.ZN (n_258), .A (n_0_204), .B1 (n_0_360), .B2 (n_0_282), .C1 (n_0_383), .C2 (n_0_281));
AOI22_X1 i_0_422 (.ZN (n_0_203), .A1 (n_8), .A2 (n_0_278), .B1 (\A_imm_2s_complement[14] ), .B2 (spc__n131));
OAI221_X1 i_0_421 (.ZN (n_257), .A (n_0_203), .B1 (n_0_359), .B2 (n_0_282), .C1 (n_0_382), .C2 (n_0_281));
AOI22_X1 i_0_418 (.ZN (n_0_201), .A1 (n_10), .A2 (n_0_278), .B1 (\A_imm_2s_complement[12] ), .B2 (spc__n131));
OAI221_X1 i_0_417 (.ZN (n_256), .A (n_0_201), .B1 (n_0_357), .B2 (n_0_282), .C1 (n_0_380), .C2 (n_0_281));
AOI22_X1 i_0_416 (.ZN (n_0_200), .A1 (n_11), .A2 (n_0_278), .B1 (\A_imm_2s_complement[11] ), .B2 (spc__n131));
OAI221_X1 i_0_415 (.ZN (n_255), .A (n_0_200), .B1 (n_0_356), .B2 (n_0_282), .C1 (n_0_379), .C2 (n_0_281));
AOI22_X1 i_0_414 (.ZN (n_0_199), .A1 (n_12), .A2 (n_0_278), .B1 (\A_imm_2s_complement[10] ), .B2 (spc__n131));
OAI221_X1 i_0_413 (.ZN (n_254), .A (n_0_199), .B1 (n_0_355), .B2 (n_0_282), .C1 (n_0_378), .C2 (n_0_281));
AOI22_X1 i_0_412 (.ZN (n_0_198), .A1 (n_13), .A2 (n_0_278), .B1 (\A_imm_2s_complement[9] ), .B2 (spc__n131));
OAI221_X1 i_0_411 (.ZN (n_253), .A (n_0_198), .B1 (n_0_354), .B2 (n_0_282), .C1 (n_0_377), .C2 (n_0_281));
AOI22_X1 i_0_410 (.ZN (n_0_197), .A1 (n_14), .A2 (n_0_278), .B1 (\A_imm_2s_complement[8] ), .B2 (spc__n131));
OAI221_X1 i_0_409 (.ZN (n_252), .A (n_0_197), .B1 (n_0_353), .B2 (n_0_282), .C1 (n_0_376), .C2 (n_0_281));
AOI22_X1 i_0_408 (.ZN (n_0_196), .A1 (n_15), .A2 (n_0_278), .B1 (\A_imm_2s_complement[7] ), .B2 (spc__n131));
OAI221_X1 i_0_407 (.ZN (n_251), .A (n_0_196), .B1 (n_0_352), .B2 (n_0_282), .C1 (n_0_375), .C2 (n_0_281));
AOI22_X1 i_0_406 (.ZN (n_0_195), .A1 (n_16), .A2 (n_0_278), .B1 (\A_imm_2s_complement[6] ), .B2 (spc__n131));
OAI221_X1 i_0_405 (.ZN (n_250), .A (n_0_195), .B1 (n_0_351), .B2 (n_0_282), .C1 (n_0_374), .C2 (n_0_281));
AOI22_X1 i_0_404 (.ZN (n_0_194), .A1 (n_17), .A2 (n_0_278), .B1 (\A_imm_2s_complement[5] ), .B2 (spc__n131));
OAI221_X1 i_0_403 (.ZN (n_249), .A (n_0_194), .B1 (n_0_350), .B2 (n_0_282), .C1 (n_0_373), .C2 (n_0_281));
AOI22_X1 i_0_402 (.ZN (n_0_193), .A1 (n_18), .A2 (n_0_278), .B1 (\A_imm_2s_complement[4] ), .B2 (spc__n131));
OAI221_X1 i_0_401 (.ZN (n_248), .A (n_0_193), .B1 (n_0_349), .B2 (n_0_282), .C1 (n_0_372), .C2 (n_0_281));
AOI22_X1 i_0_400 (.ZN (n_0_192), .A1 (n_19), .A2 (n_0_278), .B1 (\A_imm_2s_complement[3] ), .B2 (spc__n131));
OAI221_X1 i_0_399 (.ZN (n_247), .A (n_0_192), .B1 (n_0_348), .B2 (n_0_282), .C1 (n_0_371), .C2 (n_0_281));
AOI22_X1 i_0_398 (.ZN (n_0_191), .A1 (n_20), .A2 (n_0_278), .B1 (\A_imm_2s_complement[2] ), .B2 (spc__n131));
OAI221_X1 i_0_397 (.ZN (n_246), .A (n_0_191), .B1 (n_0_347), .B2 (n_0_282), .C1 (n_0_370), .C2 (n_0_281));
AOI22_X1 i_0_396 (.ZN (n_0_190), .A1 (n_21), .A2 (n_0_278), .B1 (\A_imm_2s_complement[1] ), .B2 (spc__n131));
OAI221_X1 i_0_395 (.ZN (n_245), .A (n_0_190), .B1 (n_0_346), .B2 (n_0_282), .C1 (n_0_369), .C2 (n_0_281));
NOR2_X1 i_0_392 (.ZN (n_244), .A1 (n_0_344), .A2 (n_0_279));
NOR3_X1 i_0_390 (.ZN (n_243), .A1 (n_0_188), .A2 (n_0_391), .A3 (n_0_243));
INV_X1 i_0_386 (.ZN (n_0_184), .A (spc__n134));
OAI222_X1 i_0_383 (.ZN (n_242), .A1 (n_0_60), .A2 (n_0_184), .B1 (n_0_28), .B2 (n_0_244)
    , .C1 (n_0_391), .C2 (n_0_249));
AOI22_X1 i_0_381 (.ZN (n_0_180), .A1 (n_0), .A2 (n_0_245), .B1 (\A_imm_2s_complement[22] ), .B2 (spc__n134));
OAI221_X1 i_0_380 (.ZN (n_241), .A (n_0_180), .B1 (n_0_28), .B2 (n_0_248), .C1 (n_0_60), .C2 (n_0_249));
AOI22_X1 i_0_379 (.ZN (n_0_179), .A1 (n_1), .A2 (n_0_245), .B1 (\A_imm_2s_complement[21] ), .B2 (spc__n134));
OAI221_X1 i_0_378 (.ZN (n_240), .A (n_0_179), .B1 (n_0_31), .B2 (n_0_248), .C1 (n_0_27), .C2 (n_0_249));
AOI22_X1 i_0_377 (.ZN (n_0_178), .A1 (n_2), .A2 (n_0_245), .B1 (\A_imm_2s_complement[20] ), .B2 (spc__n134));
OAI221_X1 i_0_376 (.ZN (n_239), .A (n_0_178), .B1 (n_0_365), .B2 (n_0_248), .C1 (n_0_388), .C2 (n_0_249));
AOI22_X1 i_0_375 (.ZN (n_0_177), .A1 (n_3), .A2 (n_0_245), .B1 (\A_imm_2s_complement[19] ), .B2 (spc__n134));
OAI221_X1 i_0_374 (.ZN (n_238), .A (n_0_177), .B1 (n_0_404), .B2 (n_0_248), .C1 (n_0_403), .C2 (n_0_249));
AOI22_X1 i_0_373 (.ZN (n_0_176), .A1 (n_4), .A2 (n_0_245), .B1 (\A_imm_2s_complement[18] ), .B2 (spc__n134));
OAI221_X1 i_0_372 (.ZN (n_237), .A (n_0_176), .B1 (n_0_363), .B2 (n_0_248), .C1 (n_0_386), .C2 (n_0_249));
AOI22_X1 i_0_371 (.ZN (n_0_175), .A1 (n_5), .A2 (n_0_245), .B1 (\A_imm_2s_complement[17] ), .B2 (spc__n134));
OAI221_X1 i_0_370 (.ZN (n_236), .A (n_0_175), .B1 (n_0_310), .B2 (n_0_248), .C1 (n_0_385), .C2 (n_0_249));
AOI22_X1 i_0_369 (.ZN (n_0_174), .A1 (n_6), .A2 (n_0_245), .B1 (\A_imm_2s_complement[16] ), .B2 (spc__n134));
OAI221_X1 i_0_368 (.ZN (n_235), .A (n_0_174), .B1 (n_0_361), .B2 (n_0_248), .C1 (n_0_384), .C2 (n_0_249));
AOI22_X1 i_0_367 (.ZN (n_0_173), .A1 (n_7), .A2 (n_0_245), .B1 (\A_imm_2s_complement[15] ), .B2 (spc__n134));
OAI221_X1 i_0_366 (.ZN (n_234), .A (n_0_173), .B1 (n_0_360), .B2 (n_0_248), .C1 (n_0_383), .C2 (n_0_249));
AOI22_X1 i_0_365 (.ZN (n_0_172), .A1 (n_8), .A2 (n_0_245), .B1 (\A_imm_2s_complement[14] ), .B2 (spc__n134));
OAI221_X1 i_0_364 (.ZN (n_233), .A (n_0_172), .B1 (n_0_359), .B2 (n_0_248), .C1 (n_0_382), .C2 (n_0_249));
AOI22_X1 i_0_363 (.ZN (n_0_171), .A1 (n_9), .A2 (n_0_245), .B1 (\A_imm_2s_complement[13] ), .B2 (spc__n134));
OAI221_X1 i_0_362 (.ZN (n_232), .A (n_0_171), .B1 (n_0_306), .B2 (n_0_248), .C1 (n_0_305), .C2 (n_0_249));
AOI22_X1 i_0_361 (.ZN (n_0_170), .A1 (n_10), .A2 (n_0_245), .B1 (\A_imm_2s_complement[12] ), .B2 (spc__n134));
OAI221_X1 i_0_360 (.ZN (n_231), .A (n_0_170), .B1 (n_0_357), .B2 (n_0_248), .C1 (n_0_380), .C2 (n_0_249));
AOI22_X1 i_0_359 (.ZN (n_0_169), .A1 (n_11), .A2 (n_0_245), .B1 (\A_imm_2s_complement[11] ), .B2 (spc__n134));
OAI221_X1 i_0_358 (.ZN (n_230), .A (n_0_169), .B1 (n_0_356), .B2 (n_0_248), .C1 (n_0_379), .C2 (n_0_249));
AOI22_X1 i_0_357 (.ZN (n_0_168), .A1 (n_12), .A2 (n_0_245), .B1 (\A_imm_2s_complement[10] ), .B2 (spc__n134));
OAI221_X1 i_0_356 (.ZN (n_229), .A (n_0_168), .B1 (n_0_355), .B2 (n_0_248), .C1 (n_0_378), .C2 (n_0_249));
AOI22_X1 i_0_355 (.ZN (n_0_167), .A1 (n_13), .A2 (n_0_245), .B1 (\A_imm_2s_complement[9] ), .B2 (spc__n134));
OAI221_X1 i_0_354 (.ZN (n_228), .A (n_0_167), .B1 (n_0_354), .B2 (n_0_248), .C1 (n_0_377), .C2 (n_0_249));
AOI22_X1 i_0_353 (.ZN (n_0_166), .A1 (n_14), .A2 (n_0_245), .B1 (\A_imm_2s_complement[8] ), .B2 (spc__n134));
OAI221_X1 i_0_352 (.ZN (n_227), .A (n_0_166), .B1 (n_0_353), .B2 (n_0_248), .C1 (n_0_376), .C2 (n_0_249));
AOI22_X1 i_0_351 (.ZN (n_0_165), .A1 (n_15), .A2 (n_0_245), .B1 (\A_imm_2s_complement[7] ), .B2 (spc__n134));
OAI221_X1 i_0_350 (.ZN (n_226), .A (n_0_165), .B1 (n_0_352), .B2 (n_0_248), .C1 (n_0_375), .C2 (n_0_249));
AOI22_X1 i_0_349 (.ZN (n_0_164), .A1 (n_16), .A2 (n_0_245), .B1 (\A_imm_2s_complement[6] ), .B2 (spc__n134));
OAI221_X1 i_0_348 (.ZN (n_225), .A (n_0_164), .B1 (n_0_351), .B2 (n_0_248), .C1 (n_0_374), .C2 (n_0_249));
AOI22_X1 i_0_347 (.ZN (n_0_163), .A1 (n_17), .A2 (n_0_245), .B1 (\A_imm_2s_complement[5] ), .B2 (spc__n134));
OAI221_X1 i_0_346 (.ZN (n_224), .A (n_0_163), .B1 (n_0_350), .B2 (n_0_248), .C1 (n_0_373), .C2 (n_0_249));
AOI22_X1 i_0_345 (.ZN (n_0_162), .A1 (n_18), .A2 (n_0_245), .B1 (\A_imm_2s_complement[4] ), .B2 (spc__n134));
OAI221_X1 i_0_344 (.ZN (n_223), .A (n_0_162), .B1 (n_0_349), .B2 (n_0_248), .C1 (n_0_372), .C2 (n_0_249));
AOI22_X1 i_0_343 (.ZN (n_0_161), .A1 (n_19), .A2 (n_0_245), .B1 (\A_imm_2s_complement[3] ), .B2 (spc__n134));
OAI221_X1 i_0_342 (.ZN (n_222), .A (n_0_161), .B1 (n_0_348), .B2 (n_0_248), .C1 (n_0_371), .C2 (n_0_249));
AOI22_X1 i_0_341 (.ZN (n_0_160), .A1 (n_20), .A2 (n_0_245), .B1 (\A_imm_2s_complement[2] ), .B2 (spc__n134));
OAI221_X1 i_0_340 (.ZN (n_221), .A (n_0_160), .B1 (n_0_347), .B2 (n_0_248), .C1 (n_0_370), .C2 (n_0_249));
AOI22_X1 i_0_339 (.ZN (n_0_159), .A1 (n_21), .A2 (n_0_245), .B1 (\A_imm_2s_complement[1] ), .B2 (spc__n134));
OAI221_X1 i_0_338 (.ZN (n_220), .A (n_0_159), .B1 (n_0_346), .B2 (n_0_248), .C1 (n_0_369), .C2 (n_0_249));
NOR2_X1 i_0_335 (.ZN (n_219), .A1 (n_0_344), .A2 (n_0_247));
NOR3_X1 i_0_333 (.ZN (n_218), .A1 (n_0_155), .A2 (n_0_391), .A3 (n_0_202));
INV_X1 i_0_329 (.ZN (n_0_153), .A (drc_ipo_n30));
OAI222_X1 i_0_326 (.ZN (n_217), .A1 (n_0_60), .A2 (n_0_153), .B1 (n_0_28), .B2 (n_0_206)
    , .C1 (n_0_391), .C2 (n_0_216));
AOI22_X1 i_0_324 (.ZN (n_0_149), .A1 (n_0), .A2 (n_0_212), .B1 (\A_imm_2s_complement[22] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_323 (.ZN (n_216), .A (n_0_149), .B1 (n_0_28), .B2 (n_0_214), .C1 (n_0_60), .C2 (n_0_216));
AOI22_X1 i_0_322 (.ZN (n_0_148), .A1 (n_1), .A2 (n_0_212), .B1 (\A_imm_2s_complement[21] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_321 (.ZN (n_215), .A (n_0_148), .B1 (n_0_31), .B2 (n_0_214), .C1 (n_0_27), .C2 (n_0_216));
AOI22_X1 i_0_320 (.ZN (n_0_147), .A1 (n_2), .A2 (n_0_212), .B1 (\A_imm_2s_complement[20] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_319 (.ZN (n_214), .A (n_0_147), .B1 (n_0_365), .B2 (n_0_214), .C1 (n_0_388), .C2 (n_0_216));
AOI22_X1 i_0_318 (.ZN (n_0_146), .A1 (n_3), .A2 (n_0_212), .B1 (\A_imm_2s_complement[19] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_317 (.ZN (n_213), .A (n_0_146), .B1 (n_0_404), .B2 (n_0_214), .C1 (n_0_403), .C2 (n_0_216));
AOI22_X1 i_0_316 (.ZN (n_0_145), .A1 (n_4), .A2 (n_0_212), .B1 (\A_imm_2s_complement[18] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_315 (.ZN (n_212), .A (n_0_145), .B1 (n_0_363), .B2 (n_0_214), .C1 (n_0_386), .C2 (n_0_216));
AOI22_X1 i_0_314 (.ZN (n_0_144), .A1 (n_5), .A2 (n_0_212), .B1 (\A_imm_2s_complement[17] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_313 (.ZN (n_211), .A (n_0_144), .B1 (n_0_310), .B2 (n_0_214), .C1 (n_0_385), .C2 (n_0_216));
AOI22_X1 i_0_312 (.ZN (n_0_143), .A1 (n_6), .A2 (n_0_212), .B1 (\A_imm_2s_complement[16] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_311 (.ZN (n_210), .A (n_0_143), .B1 (n_0_361), .B2 (n_0_214), .C1 (n_0_384), .C2 (n_0_216));
AOI22_X1 i_0_310 (.ZN (n_0_142), .A1 (n_7), .A2 (n_0_212), .B1 (\A_imm_2s_complement[15] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_309 (.ZN (n_209), .A (n_0_142), .B1 (n_0_360), .B2 (n_0_214), .C1 (n_0_383), .C2 (n_0_216));
AOI22_X1 i_0_308 (.ZN (n_0_141), .A1 (n_8), .A2 (n_0_212), .B1 (\A_imm_2s_complement[14] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_307 (.ZN (n_208), .A (n_0_141), .B1 (n_0_359), .B2 (n_0_214), .C1 (n_0_382), .C2 (n_0_216));
AOI22_X1 i_0_306 (.ZN (n_0_140), .A1 (n_9), .A2 (n_0_212), .B1 (\A_imm_2s_complement[13] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_305 (.ZN (n_207), .A (n_0_140), .B1 (n_0_306), .B2 (n_0_214), .C1 (n_0_305), .C2 (n_0_216));
AOI22_X1 i_0_304 (.ZN (n_0_139), .A1 (n_10), .A2 (n_0_212), .B1 (\A_imm_2s_complement[12] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_303 (.ZN (n_206), .A (n_0_139), .B1 (n_0_357), .B2 (n_0_214), .C1 (n_0_380), .C2 (n_0_216));
AOI22_X1 i_0_302 (.ZN (n_0_138), .A1 (n_11), .A2 (n_0_212), .B1 (\A_imm_2s_complement[11] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_301 (.ZN (n_205), .A (n_0_138), .B1 (n_0_356), .B2 (n_0_214), .C1 (n_0_379), .C2 (n_0_216));
AOI22_X1 i_0_300 (.ZN (n_0_137), .A1 (n_12), .A2 (n_0_212), .B1 (\A_imm_2s_complement[10] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_299 (.ZN (n_204), .A (n_0_137), .B1 (n_0_355), .B2 (n_0_214), .C1 (n_0_378), .C2 (n_0_216));
AOI22_X1 i_0_298 (.ZN (n_0_136), .A1 (n_13), .A2 (n_0_212), .B1 (\A_imm_2s_complement[9] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_297 (.ZN (n_203), .A (n_0_136), .B1 (n_0_354), .B2 (n_0_214), .C1 (n_0_377), .C2 (n_0_216));
AOI22_X1 i_0_296 (.ZN (n_0_135), .A1 (n_14), .A2 (n_0_212), .B1 (\A_imm_2s_complement[8] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_295 (.ZN (n_202), .A (n_0_135), .B1 (n_0_353), .B2 (n_0_214), .C1 (n_0_376), .C2 (n_0_216));
AOI22_X1 i_0_294 (.ZN (n_0_134), .A1 (n_15), .A2 (n_0_212), .B1 (\A_imm_2s_complement[7] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_293 (.ZN (n_201), .A (n_0_134), .B1 (n_0_352), .B2 (n_0_214), .C1 (n_0_375), .C2 (n_0_216));
AOI22_X1 i_0_292 (.ZN (n_0_133), .A1 (n_16), .A2 (n_0_212), .B1 (\A_imm_2s_complement[6] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_291 (.ZN (n_200), .A (n_0_133), .B1 (n_0_351), .B2 (n_0_214), .C1 (n_0_374), .C2 (n_0_216));
AOI22_X1 i_0_290 (.ZN (n_0_132), .A1 (n_17), .A2 (n_0_212), .B1 (\A_imm_2s_complement[5] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_289 (.ZN (n_199), .A (n_0_132), .B1 (n_0_350), .B2 (n_0_214), .C1 (n_0_373), .C2 (n_0_216));
AOI22_X1 i_0_288 (.ZN (n_0_131), .A1 (n_18), .A2 (n_0_212), .B1 (\A_imm_2s_complement[4] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_287 (.ZN (n_198), .A (n_0_131), .B1 (n_0_349), .B2 (n_0_214), .C1 (n_0_372), .C2 (n_0_216));
AOI22_X1 i_0_286 (.ZN (n_0_130), .A1 (n_19), .A2 (n_0_212), .B1 (\A_imm_2s_complement[3] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_285 (.ZN (n_197), .A (n_0_130), .B1 (n_0_348), .B2 (n_0_214), .C1 (n_0_371), .C2 (n_0_216));
AOI22_X1 i_0_284 (.ZN (n_0_129), .A1 (n_20), .A2 (n_0_212), .B1 (\A_imm_2s_complement[2] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_283 (.ZN (n_196), .A (n_0_129), .B1 (n_0_347), .B2 (n_0_214), .C1 (n_0_370), .C2 (n_0_216));
AOI22_X1 i_0_282 (.ZN (n_0_128), .A1 (n_21), .A2 (n_0_212), .B1 (\A_imm_2s_complement[1] ), .B2 (drc_ipo_n30));
OAI221_X1 i_0_281 (.ZN (n_195), .A (n_0_128), .B1 (n_0_346), .B2 (n_0_214), .C1 (n_0_369), .C2 (n_0_216));
NOR2_X1 i_0_278 (.ZN (n_194), .A1 (n_0_344), .A2 (n_0_213));
NOR3_X1 i_0_276 (.ZN (n_193), .A1 (n_0_120), .A2 (n_0_391), .A3 (n_0_157));
INV_X1 i_0_109 (.ZN (n_0_122), .A (drc_ipo_n31));
OAI222_X1 i_0_108 (.ZN (n_192), .A1 (n_0_60), .A2 (n_0_122), .B1 (n_0_28), .B2 (n_0_158)
    , .C1 (n_0_391), .C2 (n_0_185));
AOI22_X1 i_0_267 (.ZN (n_0_118), .A1 (n_0), .A2 (n_0_181), .B1 (\A_imm_2s_complement[22] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_266 (.ZN (n_191), .A (n_0_118), .B1 (n_0_28), .B2 (n_0_183), .C1 (n_0_60), .C2 (n_0_185));
AOI22_X1 i_0_265 (.ZN (n_0_117), .A1 (n_1), .A2 (n_0_181), .B1 (\A_imm_2s_complement[21] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_264 (.ZN (n_190), .A (n_0_117), .B1 (n_0_31), .B2 (n_0_183), .C1 (n_0_27), .C2 (n_0_185));
AOI22_X1 i_0_263 (.ZN (n_0_116), .A1 (n_2), .A2 (n_0_181), .B1 (\A_imm_2s_complement[20] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_262 (.ZN (n_189), .A (n_0_116), .B1 (n_0_365), .B2 (n_0_183), .C1 (n_0_388), .C2 (n_0_185));
AOI22_X1 i_0_261 (.ZN (n_0_115), .A1 (n_3), .A2 (n_0_181), .B1 (\A_imm_2s_complement[19] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_260 (.ZN (n_188), .A (n_0_115), .B1 (n_0_404), .B2 (n_0_183), .C1 (n_0_403), .C2 (n_0_185));
AOI22_X1 i_0_259 (.ZN (n_0_114), .A1 (n_4), .A2 (n_0_181), .B1 (\A_imm_2s_complement[18] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_258 (.ZN (n_187), .A (n_0_114), .B1 (n_0_363), .B2 (n_0_183), .C1 (n_0_386), .C2 (n_0_185));
AOI22_X1 i_0_257 (.ZN (n_0_113), .A1 (n_5), .A2 (n_0_181), .B1 (\A_imm_2s_complement[17] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_256 (.ZN (n_186), .A (n_0_113), .B1 (n_0_310), .B2 (n_0_183), .C1 (n_0_385), .C2 (n_0_185));
AOI22_X1 i_0_255 (.ZN (n_0_112), .A1 (n_6), .A2 (n_0_181), .B1 (\A_imm_2s_complement[16] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_254 (.ZN (n_185), .A (n_0_112), .B1 (n_0_361), .B2 (n_0_183), .C1 (n_0_384), .C2 (n_0_185));
AOI22_X1 i_0_253 (.ZN (n_0_111), .A1 (n_7), .A2 (n_0_181), .B1 (\A_imm_2s_complement[15] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_252 (.ZN (n_184), .A (n_0_111), .B1 (n_0_360), .B2 (n_0_183), .C1 (n_0_383), .C2 (n_0_185));
AOI22_X1 i_0_251 (.ZN (n_0_110), .A1 (n_8), .A2 (n_0_181), .B1 (\A_imm_2s_complement[14] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_250 (.ZN (n_183), .A (n_0_110), .B1 (n_0_359), .B2 (n_0_183), .C1 (n_0_382), .C2 (n_0_185));
AOI22_X1 i_0_249 (.ZN (n_0_109), .A1 (n_9), .A2 (n_0_181), .B1 (\A_imm_2s_complement[13] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_248 (.ZN (n_182), .A (n_0_109), .B1 (n_0_306), .B2 (n_0_183), .C1 (n_0_305), .C2 (n_0_185));
AOI22_X1 i_0_247 (.ZN (n_0_108), .A1 (n_10), .A2 (n_0_181), .B1 (\A_imm_2s_complement[12] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_246 (.ZN (n_181), .A (n_0_108), .B1 (n_0_357), .B2 (n_0_183), .C1 (n_0_380), .C2 (n_0_185));
AOI22_X1 i_0_245 (.ZN (n_0_107), .A1 (n_11), .A2 (n_0_181), .B1 (\A_imm_2s_complement[11] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_244 (.ZN (n_180), .A (n_0_107), .B1 (n_0_356), .B2 (n_0_183), .C1 (n_0_379), .C2 (n_0_185));
AOI22_X1 i_0_243 (.ZN (n_0_106), .A1 (n_12), .A2 (n_0_181), .B1 (\A_imm_2s_complement[10] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_242 (.ZN (n_179), .A (n_0_106), .B1 (n_0_355), .B2 (n_0_183), .C1 (n_0_378), .C2 (n_0_185));
AOI22_X1 i_0_241 (.ZN (n_0_105), .A1 (n_13), .A2 (n_0_181), .B1 (\A_imm_2s_complement[9] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_240 (.ZN (n_178), .A (n_0_105), .B1 (n_0_354), .B2 (n_0_183), .C1 (n_0_377), .C2 (n_0_185));
AOI22_X1 i_0_239 (.ZN (n_0_104), .A1 (n_14), .A2 (n_0_181), .B1 (\A_imm_2s_complement[8] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_238 (.ZN (n_177), .A (n_0_104), .B1 (n_0_353), .B2 (n_0_183), .C1 (n_0_376), .C2 (n_0_185));
AOI22_X1 i_0_237 (.ZN (n_0_103), .A1 (n_15), .A2 (n_0_181), .B1 (\A_imm_2s_complement[7] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_236 (.ZN (n_176), .A (n_0_103), .B1 (n_0_352), .B2 (n_0_183), .C1 (n_0_375), .C2 (n_0_185));
AOI22_X1 i_0_235 (.ZN (n_0_102), .A1 (n_16), .A2 (n_0_181), .B1 (\A_imm_2s_complement[6] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_234 (.ZN (n_175), .A (n_0_102), .B1 (n_0_351), .B2 (n_0_183), .C1 (n_0_374), .C2 (n_0_185));
AOI22_X1 i_0_233 (.ZN (n_0_101), .A1 (n_17), .A2 (n_0_181), .B1 (\A_imm_2s_complement[5] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_232 (.ZN (n_174), .A (n_0_101), .B1 (n_0_350), .B2 (n_0_183), .C1 (n_0_373), .C2 (n_0_185));
AOI22_X1 i_0_231 (.ZN (n_0_100), .A1 (n_18), .A2 (n_0_181), .B1 (\A_imm_2s_complement[4] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_230 (.ZN (n_173), .A (n_0_100), .B1 (n_0_349), .B2 (n_0_183), .C1 (n_0_372), .C2 (n_0_185));
AOI22_X1 i_0_229 (.ZN (n_0_99), .A1 (n_19), .A2 (n_0_181), .B1 (\A_imm_2s_complement[3] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_228 (.ZN (n_172), .A (n_0_99), .B1 (n_0_348), .B2 (n_0_183), .C1 (n_0_371), .C2 (n_0_185));
AOI22_X1 i_0_227 (.ZN (n_0_98), .A1 (n_20), .A2 (n_0_181), .B1 (\A_imm_2s_complement[2] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_226 (.ZN (n_171), .A (n_0_98), .B1 (n_0_347), .B2 (n_0_183), .C1 (n_0_370), .C2 (n_0_185));
AOI22_X1 i_0_225 (.ZN (n_0_97), .A1 (n_21), .A2 (n_0_181), .B1 (\A_imm_2s_complement[1] ), .B2 (drc_ipo_n31));
OAI221_X1 i_0_224 (.ZN (n_170), .A (n_0_97), .B1 (n_0_346), .B2 (n_0_183), .C1 (n_0_369), .C2 (n_0_185));
NOR2_X1 i_0_221 (.ZN (n_169), .A1 (n_0_344), .A2 (n_0_182));
NOR3_X1 i_0_219 (.ZN (n_168), .A1 (n_0_63), .A2 (n_0_391), .A3 (n_0_123));
INV_X1 i_0_213 (.ZN (n_0_89), .A (n_0_126));
OAI222_X1 i_0_212 (.ZN (n_167), .A1 (n_0_28), .A2 (n_0_124), .B1 (n_0_60), .B2 (n_0_89)
    , .C1 (n_0_391), .C2 (n_0_150));
AOI22_X1 i_0_210 (.ZN (n_0_87), .A1 (\A_imm_2s_complement[22] ), .A2 (n_0_126), .B1 (n_0), .B2 (n_0_125));
OAI221_X1 i_0_209 (.ZN (n_166), .A (n_0_87), .B1 (n_0_28), .B2 (n_0_151), .C1 (n_0_60), .C2 (n_0_150));
AOI22_X1 i_0_208 (.ZN (n_0_86), .A1 (\A_imm_2s_complement[21] ), .A2 (n_0_126), .B1 (n_1), .B2 (n_0_125));
OAI221_X1 i_0_207 (.ZN (n_165), .A (n_0_86), .B1 (n_0_31), .B2 (n_0_151), .C1 (n_0_27), .C2 (n_0_150));
AOI22_X1 i_0_206 (.ZN (n_0_85), .A1 (\A_imm_2s_complement[20] ), .A2 (n_0_126), .B1 (n_2), .B2 (n_0_125));
OAI221_X1 i_0_205 (.ZN (n_164), .A (n_0_85), .B1 (n_0_365), .B2 (n_0_151), .C1 (n_0_388), .C2 (n_0_150));
AOI22_X1 i_0_204 (.ZN (n_0_84), .A1 (\A_imm_2s_complement[19] ), .A2 (n_0_126), .B1 (n_3), .B2 (n_0_125));
OAI221_X1 i_0_203 (.ZN (n_163), .A (n_0_84), .B1 (n_0_404), .B2 (n_0_151), .C1 (n_0_403), .C2 (n_0_150));
AOI22_X1 i_0_202 (.ZN (n_0_83), .A1 (\A_imm_2s_complement[18] ), .A2 (n_0_126), .B1 (n_4), .B2 (n_0_125));
OAI221_X1 i_0_201 (.ZN (n_162), .A (n_0_83), .B1 (n_0_363), .B2 (n_0_151), .C1 (n_0_386), .C2 (n_0_150));
AOI22_X1 i_0_200 (.ZN (n_0_82), .A1 (\A_imm_2s_complement[17] ), .A2 (n_0_126), .B1 (n_5), .B2 (n_0_125));
OAI221_X1 i_0_199 (.ZN (n_161), .A (n_0_82), .B1 (n_0_310), .B2 (n_0_151), .C1 (n_0_385), .C2 (n_0_150));
AOI22_X1 i_0_198 (.ZN (n_0_81), .A1 (\A_imm_2s_complement[16] ), .A2 (n_0_126), .B1 (n_6), .B2 (n_0_125));
OAI221_X1 i_0_197 (.ZN (n_160), .A (n_0_81), .B1 (n_0_361), .B2 (n_0_151), .C1 (n_0_384), .C2 (n_0_150));
AOI22_X1 i_0_196 (.ZN (n_0_80), .A1 (\A_imm_2s_complement[15] ), .A2 (n_0_126), .B1 (n_7), .B2 (n_0_125));
OAI221_X1 i_0_195 (.ZN (n_159), .A (n_0_80), .B1 (n_0_360), .B2 (n_0_151), .C1 (n_0_383), .C2 (n_0_150));
AOI22_X1 i_0_194 (.ZN (n_0_79), .A1 (\A_imm_2s_complement[14] ), .A2 (n_0_126), .B1 (n_8), .B2 (n_0_125));
OAI221_X1 i_0_193 (.ZN (n_158), .A (n_0_79), .B1 (n_0_359), .B2 (n_0_151), .C1 (n_0_382), .C2 (n_0_150));
AOI22_X1 i_0_192 (.ZN (n_0_78), .A1 (\A_imm_2s_complement[13] ), .A2 (n_0_126), .B1 (n_9), .B2 (n_0_125));
OAI221_X1 i_0_191 (.ZN (n_157), .A (n_0_78), .B1 (n_0_306), .B2 (n_0_151), .C1 (n_0_305), .C2 (n_0_150));
AOI22_X1 i_0_190 (.ZN (n_0_77), .A1 (\A_imm_2s_complement[12] ), .A2 (n_0_126), .B1 (n_10), .B2 (n_0_125));
OAI221_X1 i_0_189 (.ZN (n_156), .A (n_0_77), .B1 (n_0_357), .B2 (n_0_151), .C1 (n_0_380), .C2 (n_0_150));
AOI22_X1 i_0_188 (.ZN (n_0_76), .A1 (\A_imm_2s_complement[11] ), .A2 (n_0_126), .B1 (n_11), .B2 (n_0_125));
OAI221_X1 i_0_187 (.ZN (n_155), .A (n_0_76), .B1 (n_0_356), .B2 (n_0_151), .C1 (n_0_379), .C2 (n_0_150));
AOI22_X1 i_0_186 (.ZN (n_0_75), .A1 (\A_imm_2s_complement[10] ), .A2 (n_0_126), .B1 (n_12), .B2 (n_0_125));
OAI221_X1 i_0_185 (.ZN (n_154), .A (n_0_75), .B1 (n_0_355), .B2 (n_0_151), .C1 (n_0_378), .C2 (n_0_150));
AOI22_X1 i_0_184 (.ZN (n_0_74), .A1 (\A_imm_2s_complement[9] ), .A2 (n_0_126), .B1 (n_13), .B2 (n_0_125));
OAI221_X1 i_0_183 (.ZN (n_153), .A (n_0_74), .B1 (n_0_354), .B2 (n_0_151), .C1 (n_0_377), .C2 (n_0_150));
AOI22_X1 i_0_182 (.ZN (n_0_73), .A1 (\A_imm_2s_complement[8] ), .A2 (n_0_126), .B1 (n_14), .B2 (n_0_125));
OAI221_X1 i_0_181 (.ZN (n_152), .A (n_0_73), .B1 (n_0_353), .B2 (n_0_151), .C1 (n_0_376), .C2 (n_0_150));
AOI22_X1 i_0_180 (.ZN (n_0_72), .A1 (\A_imm_2s_complement[7] ), .A2 (n_0_126), .B1 (n_15), .B2 (n_0_125));
OAI221_X1 i_0_179 (.ZN (n_151), .A (n_0_72), .B1 (n_0_352), .B2 (n_0_151), .C1 (n_0_375), .C2 (n_0_150));
AOI22_X1 i_0_178 (.ZN (n_0_71), .A1 (\A_imm_2s_complement[6] ), .A2 (n_0_126), .B1 (n_16), .B2 (n_0_125));
OAI221_X1 i_0_177 (.ZN (n_150), .A (n_0_71), .B1 (n_0_351), .B2 (n_0_151), .C1 (n_0_374), .C2 (n_0_150));
AOI22_X1 i_0_176 (.ZN (n_0_70), .A1 (\A_imm_2s_complement[5] ), .A2 (n_0_126), .B1 (n_17), .B2 (n_0_125));
OAI221_X1 i_0_175 (.ZN (n_149), .A (n_0_70), .B1 (n_0_350), .B2 (n_0_151), .C1 (n_0_373), .C2 (n_0_150));
AOI22_X1 i_0_174 (.ZN (n_0_69), .A1 (\A_imm_2s_complement[4] ), .A2 (n_0_126), .B1 (n_18), .B2 (n_0_125));
OAI221_X1 i_0_173 (.ZN (n_148), .A (n_0_69), .B1 (n_0_349), .B2 (n_0_151), .C1 (n_0_372), .C2 (n_0_150));
AOI22_X1 i_0_172 (.ZN (n_0_68), .A1 (\A_imm_2s_complement[3] ), .A2 (n_0_126), .B1 (n_19), .B2 (n_0_125));
OAI221_X1 i_0_171 (.ZN (n_147), .A (n_0_68), .B1 (n_0_348), .B2 (n_0_151), .C1 (n_0_371), .C2 (n_0_150));
AOI22_X1 i_0_170 (.ZN (n_0_67), .A1 (\A_imm_2s_complement[2] ), .A2 (n_0_126), .B1 (n_20), .B2 (n_0_125));
OAI221_X1 i_0_169 (.ZN (n_146), .A (n_0_67), .B1 (n_0_347), .B2 (n_0_151), .C1 (n_0_370), .C2 (n_0_150));
AOI22_X1 i_0_168 (.ZN (n_0_66), .A1 (\A_imm_2s_complement[1] ), .A2 (n_0_126), .B1 (n_21), .B2 (n_0_125));
OAI221_X1 i_0_167 (.ZN (n_145), .A (n_0_66), .B1 (n_0_346), .B2 (n_0_151), .C1 (n_0_369), .C2 (n_0_150));
NOR2_X1 i_0_164 (.ZN (n_144), .A1 (n_0_344), .A2 (n_0_127));
NOR3_X1 i_0_106 (.ZN (n_143), .A1 (n_0_33), .A2 (n_0_391), .A3 (n_0_65));
INV_X1 i_0_105 (.ZN (n_0_58), .A (spc__n136));
OAI222_X1 i_0_104 (.ZN (n_142), .A1 (n_0_28), .A2 (n_0_88), .B1 (n_0_60), .B2 (n_0_58)
    , .C1 (n_0_391), .C2 (n_0_94));
AOI22_X1 i_0_153 (.ZN (n_0_56), .A1 (\A_imm_2s_complement[22] ), .A2 (spc__n136), .B1 (n_0), .B2 (n_0_90));
OAI221_X1 i_0_152 (.ZN (n_141), .A (n_0_56), .B1 (n_0_28), .B2 (n_0_96), .C1 (n_0_60), .C2 (n_0_94));
AOI22_X1 i_0_103 (.ZN (n_0_55), .A1 (\A_imm_2s_complement[21] ), .A2 (spc__n136), .B1 (n_1), .B2 (n_0_90));
OAI221_X1 i_0_102 (.ZN (n_140), .A (n_0_55), .B1 (n_0_31), .B2 (n_0_96), .C1 (n_0_27), .C2 (n_0_94));
AOI22_X1 i_0_149 (.ZN (n_0_54), .A1 (\A_imm_2s_complement[20] ), .A2 (spc__n136), .B1 (n_2), .B2 (n_0_90));
OAI221_X1 i_0_148 (.ZN (n_139), .A (n_0_54), .B1 (n_0_365), .B2 (n_0_96), .C1 (n_0_388), .C2 (n_0_94));
AOI22_X1 i_0_147 (.ZN (n_0_53), .A1 (\A_imm_2s_complement[19] ), .A2 (spc__n136), .B1 (n_3), .B2 (n_0_90));
OAI221_X1 i_0_146 (.ZN (n_138), .A (n_0_53), .B1 (n_0_404), .B2 (n_0_96), .C1 (n_0_403), .C2 (n_0_94));
AOI22_X1 i_0_145 (.ZN (n_0_52), .A1 (\A_imm_2s_complement[18] ), .A2 (spc__n136), .B1 (n_4), .B2 (n_0_90));
OAI221_X1 i_0_144 (.ZN (n_137), .A (n_0_52), .B1 (n_0_363), .B2 (n_0_96), .C1 (n_0_386), .C2 (n_0_94));
AOI22_X1 i_0_143 (.ZN (n_0_51), .A1 (\A_imm_2s_complement[17] ), .A2 (spc__n136), .B1 (n_5), .B2 (n_0_90));
OAI221_X1 i_0_142 (.ZN (n_136), .A (n_0_51), .B1 (n_0_310), .B2 (n_0_96), .C1 (n_0_385), .C2 (n_0_94));
AOI22_X1 i_0_141 (.ZN (n_0_50), .A1 (\A_imm_2s_complement[16] ), .A2 (spc__n136), .B1 (n_6), .B2 (n_0_90));
OAI221_X1 i_0_140 (.ZN (n_135), .A (n_0_50), .B1 (n_0_361), .B2 (n_0_96), .C1 (n_0_384), .C2 (n_0_94));
AOI22_X1 i_0_139 (.ZN (n_0_49), .A1 (\A_imm_2s_complement[15] ), .A2 (spc__n136), .B1 (n_7), .B2 (n_0_90));
OAI221_X1 i_0_138 (.ZN (n_134), .A (n_0_49), .B1 (n_0_360), .B2 (n_0_96), .C1 (n_0_383), .C2 (n_0_94));
AOI22_X1 i_0_137 (.ZN (n_0_48), .A1 (\A_imm_2s_complement[14] ), .A2 (spc__n136), .B1 (n_8), .B2 (n_0_90));
OAI221_X1 i_0_136 (.ZN (n_133), .A (n_0_48), .B1 (n_0_359), .B2 (n_0_96), .C1 (n_0_382), .C2 (n_0_94));
AOI22_X1 i_0_135 (.ZN (n_0_47), .A1 (\A_imm_2s_complement[13] ), .A2 (spc__n136), .B1 (n_9), .B2 (n_0_90));
OAI221_X1 i_0_134 (.ZN (n_132), .A (n_0_47), .B1 (n_0_306), .B2 (n_0_96), .C1 (n_0_305), .C2 (n_0_94));
AOI22_X1 i_0_133 (.ZN (n_0_46), .A1 (\A_imm_2s_complement[12] ), .A2 (spc__n136), .B1 (n_10), .B2 (n_0_90));
OAI221_X1 i_0_132 (.ZN (n_131), .A (n_0_46), .B1 (n_0_357), .B2 (n_0_96), .C1 (n_0_380), .C2 (n_0_94));
AOI22_X1 i_0_131 (.ZN (n_0_45), .A1 (\A_imm_2s_complement[11] ), .A2 (spc__n136), .B1 (n_11), .B2 (n_0_90));
OAI221_X1 i_0_130 (.ZN (n_130), .A (n_0_45), .B1 (n_0_356), .B2 (n_0_96), .C1 (n_0_379), .C2 (n_0_94));
AOI22_X1 i_0_129 (.ZN (n_0_44), .A1 (\A_imm_2s_complement[10] ), .A2 (spc__n136), .B1 (n_12), .B2 (n_0_90));
OAI221_X1 i_0_128 (.ZN (n_129), .A (n_0_44), .B1 (n_0_355), .B2 (n_0_96), .C1 (n_0_378), .C2 (n_0_94));
AOI22_X1 i_0_127 (.ZN (n_0_43), .A1 (\A_imm_2s_complement[9] ), .A2 (spc__n136), .B1 (n_13), .B2 (n_0_90));
OAI221_X1 i_0_126 (.ZN (n_128), .A (n_0_43), .B1 (n_0_354), .B2 (n_0_96), .C1 (n_0_377), .C2 (n_0_94));
AOI22_X1 i_0_125 (.ZN (n_0_42), .A1 (\A_imm_2s_complement[8] ), .A2 (spc__n136), .B1 (n_14), .B2 (n_0_90));
OAI221_X1 i_0_124 (.ZN (n_127), .A (n_0_42), .B1 (n_0_353), .B2 (n_0_96), .C1 (n_0_376), .C2 (n_0_94));
AOI22_X1 i_0_123 (.ZN (n_0_41), .A1 (\A_imm_2s_complement[7] ), .A2 (spc__n136), .B1 (n_15), .B2 (n_0_90));
OAI221_X1 i_0_122 (.ZN (n_126), .A (n_0_41), .B1 (n_0_352), .B2 (n_0_96), .C1 (n_0_375), .C2 (n_0_94));
AOI22_X1 i_0_121 (.ZN (n_0_40), .A1 (\A_imm_2s_complement[6] ), .A2 (spc__n136), .B1 (n_16), .B2 (n_0_90));
OAI221_X1 i_0_120 (.ZN (n_125), .A (n_0_40), .B1 (n_0_351), .B2 (n_0_96), .C1 (n_0_374), .C2 (n_0_94));
AOI22_X1 i_0_119 (.ZN (n_0_39), .A1 (\A_imm_2s_complement[5] ), .A2 (spc__n136), .B1 (n_17), .B2 (n_0_90));
OAI221_X1 i_0_118 (.ZN (n_124), .A (n_0_39), .B1 (n_0_350), .B2 (n_0_96), .C1 (n_0_373), .C2 (n_0_94));
AOI22_X1 i_0_117 (.ZN (n_0_38), .A1 (\A_imm_2s_complement[4] ), .A2 (spc__n136), .B1 (n_18), .B2 (n_0_90));
OAI221_X1 i_0_116 (.ZN (n_123), .A (n_0_38), .B1 (n_0_349), .B2 (n_0_96), .C1 (n_0_372), .C2 (n_0_94));
AOI22_X1 i_0_115 (.ZN (n_0_37), .A1 (\A_imm_2s_complement[3] ), .A2 (spc__n136), .B1 (n_19), .B2 (n_0_90));
OAI221_X1 i_0_114 (.ZN (n_122), .A (n_0_37), .B1 (n_0_348), .B2 (n_0_96), .C1 (n_0_371), .C2 (n_0_94));
AOI22_X1 i_0_113 (.ZN (n_0_36), .A1 (\A_imm_2s_complement[2] ), .A2 (spc__n136), .B1 (n_20), .B2 (n_0_90));
OAI221_X1 i_0_112 (.ZN (n_121), .A (n_0_36), .B1 (n_0_347), .B2 (n_0_96), .C1 (n_0_370), .C2 (n_0_94));
AOI22_X1 i_0_101 (.ZN (n_0_35), .A1 (\A_imm_2s_complement[1] ), .A2 (spc__n136), .B1 (n_21), .B2 (n_0_90));
OAI221_X1 i_0_100 (.ZN (n_120), .A (n_0_35), .B1 (n_0_346), .B2 (n_0_96), .C1 (n_0_369), .C2 (n_0_94));
NOR2_X1 i_0_107 (.ZN (n_119), .A1 (n_0_344), .A2 (n_0_93));
NAND2_X1 i_0_99 (.ZN (n_0_32), .A1 (\A_imm_2s_complement[27] ), .A2 (n_46));
NOR2_X1 i_0_98 (.ZN (n_118), .A1 (n_0_57), .A2 (n_0_32));
OAI22_X1 i_0_97 (.ZN (n_117), .A1 (n_0_60), .A2 (n_0_30), .B1 (n_0_32), .B2 (n_0_61));
INV_X1 i_0_96 (.ZN (n_0_26), .A (n_0_59));
OR2_X1 i_0_95 (.ZN (n_0_25), .A1 (n_46), .A2 (n_0_61));
AOI22_X1 i_0_94 (.ZN (n_0_24), .A1 (n_1), .A2 (n_0_26), .B1 (\A_imm_2s_complement[21] ), .B2 (n_0_29));
OAI221_X1 i_0_93 (.ZN (n_116), .A (n_0_24), .B1 (n_0_31), .B2 (n_0_25), .C1 (n_0_27), .C2 (n_0_62));
AOI22_X1 i_0_92 (.ZN (n_0_23), .A1 (n_2), .A2 (n_0_26), .B1 (\A_imm_2s_complement[20] ), .B2 (n_0_29));
OAI221_X1 i_0_91 (.ZN (n_115), .A (n_0_23), .B1 (n_0_365), .B2 (n_0_25), .C1 (n_0_388), .C2 (n_0_62));
AOI22_X1 i_0_90 (.ZN (n_0_22), .A1 (n_3), .A2 (n_0_26), .B1 (\A_imm_2s_complement[19] ), .B2 (n_0_29));
OAI221_X1 i_0_89 (.ZN (n_114), .A (n_0_22), .B1 (n_0_404), .B2 (n_0_25), .C1 (n_0_403), .C2 (n_0_62));
AOI22_X1 i_0_88 (.ZN (n_0_21), .A1 (n_4), .A2 (n_0_26), .B1 (\A_imm_2s_complement[18] ), .B2 (n_0_29));
OAI221_X1 i_0_87 (.ZN (n_113), .A (n_0_21), .B1 (n_0_363), .B2 (n_0_25), .C1 (n_0_386), .C2 (n_0_62));
AOI22_X1 i_0_86 (.ZN (n_0_20), .A1 (n_5), .A2 (n_0_26), .B1 (\A_imm_2s_complement[17] ), .B2 (n_0_29));
OAI221_X1 i_0_85 (.ZN (n_112), .A (n_0_20), .B1 (n_0_310), .B2 (n_0_25), .C1 (n_0_385), .C2 (n_0_62));
AOI22_X1 i_0_84 (.ZN (n_0_19), .A1 (n_6), .A2 (n_0_26), .B1 (\A_imm_2s_complement[16] ), .B2 (n_0_29));
OAI221_X1 i_0_83 (.ZN (n_111), .A (n_0_19), .B1 (n_0_361), .B2 (n_0_25), .C1 (n_0_384), .C2 (n_0_62));
AOI22_X1 i_0_82 (.ZN (n_0_18), .A1 (n_7), .A2 (n_0_26), .B1 (\A_imm_2s_complement[15] ), .B2 (n_0_29));
OAI221_X1 i_0_81 (.ZN (n_110), .A (n_0_18), .B1 (n_0_360), .B2 (n_0_25), .C1 (n_0_383), .C2 (n_0_62));
AOI22_X1 i_0_80 (.ZN (n_0_17), .A1 (n_8), .A2 (n_0_26), .B1 (\A_imm_2s_complement[14] ), .B2 (n_0_29));
OAI221_X1 i_0_79 (.ZN (n_109), .A (n_0_17), .B1 (n_0_359), .B2 (n_0_25), .C1 (n_0_382), .C2 (n_0_62));
AOI22_X1 i_0_78 (.ZN (n_0_16), .A1 (n_9), .A2 (n_0_26), .B1 (\A_imm_2s_complement[13] ), .B2 (n_0_29));
OAI221_X1 i_0_77 (.ZN (n_108), .A (n_0_16), .B1 (n_0_306), .B2 (n_0_25), .C1 (n_0_305), .C2 (n_0_62));
AOI22_X1 i_0_76 (.ZN (n_0_15), .A1 (n_10), .A2 (n_0_26), .B1 (\A_imm_2s_complement[12] ), .B2 (n_0_29));
OAI221_X1 i_0_75 (.ZN (n_107), .A (n_0_15), .B1 (n_0_357), .B2 (n_0_25), .C1 (n_0_380), .C2 (n_0_62));
AOI22_X1 i_0_74 (.ZN (n_0_14), .A1 (n_11), .A2 (n_0_26), .B1 (\A_imm_2s_complement[11] ), .B2 (n_0_29));
OAI221_X1 i_0_73 (.ZN (n_106), .A (n_0_14), .B1 (n_0_356), .B2 (n_0_25), .C1 (n_0_379), .C2 (n_0_62));
AOI22_X1 i_0_72 (.ZN (n_0_13), .A1 (n_12), .A2 (n_0_26), .B1 (\A_imm_2s_complement[10] ), .B2 (n_0_29));
OAI221_X1 i_0_71 (.ZN (n_105), .A (n_0_13), .B1 (n_0_355), .B2 (n_0_25), .C1 (n_0_378), .C2 (n_0_62));
AOI22_X1 i_0_70 (.ZN (n_0_12), .A1 (n_13), .A2 (n_0_26), .B1 (\A_imm_2s_complement[9] ), .B2 (n_0_29));
OAI221_X1 i_0_69 (.ZN (n_104), .A (n_0_12), .B1 (n_0_354), .B2 (n_0_25), .C1 (n_0_377), .C2 (n_0_62));
AOI22_X1 i_0_68 (.ZN (n_0_11), .A1 (n_14), .A2 (n_0_26), .B1 (\A_imm_2s_complement[8] ), .B2 (n_0_29));
OAI221_X1 i_0_67 (.ZN (n_103), .A (n_0_11), .B1 (n_0_353), .B2 (n_0_25), .C1 (n_0_376), .C2 (n_0_62));
AOI22_X1 i_0_66 (.ZN (n_0_10), .A1 (n_15), .A2 (n_0_26), .B1 (\A_imm_2s_complement[7] ), .B2 (n_0_29));
OAI221_X1 i_0_65 (.ZN (n_102), .A (n_0_10), .B1 (n_0_352), .B2 (n_0_25), .C1 (n_0_375), .C2 (n_0_62));
AOI22_X1 i_0_64 (.ZN (n_0_9), .A1 (n_16), .A2 (n_0_26), .B1 (\A_imm_2s_complement[6] ), .B2 (n_0_29));
OAI221_X1 i_0_63 (.ZN (n_101), .A (n_0_9), .B1 (n_0_351), .B2 (n_0_25), .C1 (n_0_374), .C2 (n_0_62));
AOI22_X1 i_0_62 (.ZN (n_0_8), .A1 (n_17), .A2 (n_0_26), .B1 (\A_imm_2s_complement[5] ), .B2 (n_0_29));
OAI221_X1 i_0_61 (.ZN (n_100), .A (n_0_8), .B1 (n_0_350), .B2 (n_0_25), .C1 (n_0_373), .C2 (n_0_62));
AOI22_X1 i_0_60 (.ZN (n_0_7), .A1 (n_18), .A2 (n_0_26), .B1 (\A_imm_2s_complement[4] ), .B2 (n_0_29));
OAI221_X1 i_0_59 (.ZN (n_99), .A (n_0_7), .B1 (n_0_349), .B2 (n_0_25), .C1 (n_0_372), .C2 (n_0_62));
AOI22_X1 i_0_58 (.ZN (n_0_6), .A1 (n_19), .A2 (n_0_26), .B1 (\A_imm_2s_complement[3] ), .B2 (n_0_29));
OAI221_X1 i_0_57 (.ZN (n_98), .A (n_0_6), .B1 (n_0_348), .B2 (n_0_25), .C1 (n_0_371), .C2 (n_0_62));
AOI22_X1 i_0_56 (.ZN (n_0_5), .A1 (n_20), .A2 (n_0_26), .B1 (\A_imm_2s_complement[2] ), .B2 (n_0_29));
OAI221_X1 i_0_55 (.ZN (n_97), .A (n_0_5), .B1 (n_0_347), .B2 (n_0_25), .C1 (n_0_370), .C2 (n_0_62));
AOI22_X1 i_0_54 (.ZN (n_0_4), .A1 (n_21), .A2 (n_0_26), .B1 (\A_imm_2s_complement[1] ), .B2 (n_0_29));
OAI221_X1 i_0_53 (.ZN (n_96), .A (n_0_4), .B1 (n_0_346), .B2 (n_0_25), .C1 (n_0_369), .C2 (n_0_62));
OAI21_X1 i_0_52 (.ZN (n_0_3), .A (n_22), .B1 (n_0_29), .B2 (n_0_26));
OAI221_X1 i_0_51 (.ZN (n_95), .A (n_0_3), .B1 (n_0_95), .B2 (n_0_25), .C1 (n_0_92), .C2 (n_0_62));
NOR2_X1 i_0_50 (.ZN (n_94), .A1 (n_0_344), .A2 (n_0_61));
NOR2_X1 i_0_49 (.ZN (n_93), .A1 (n_0_28), .A2 (n_0_31));
NOR2_X1 i_0_48 (.ZN (n_92), .A1 (n_0_28), .A2 (n_0_365));
NOR2_X1 i_0_47 (.ZN (n_91), .A1 (n_0_28), .A2 (n_0_404));
NOR2_X1 i_0_46 (.ZN (n_90), .A1 (n_0_28), .A2 (n_0_363));
NOR2_X1 i_0_45 (.ZN (n_89), .A1 (n_0_28), .A2 (n_0_310));
NOR2_X1 i_0_44 (.ZN (n_88), .A1 (n_0_28), .A2 (n_0_361));
NOR2_X1 i_0_43 (.ZN (n_87), .A1 (n_0_28), .A2 (n_0_360));
NOR2_X1 i_0_42 (.ZN (n_86), .A1 (n_0_28), .A2 (n_0_359));
NOR2_X1 i_0_41 (.ZN (n_85), .A1 (n_0_28), .A2 (n_0_306));
NOR2_X1 i_0_40 (.ZN (n_84), .A1 (n_0_28), .A2 (n_0_357));
NOR2_X1 i_0_39 (.ZN (n_83), .A1 (n_0_28), .A2 (n_0_356));
NOR2_X1 i_0_38 (.ZN (n_82), .A1 (n_0_28), .A2 (n_0_355));
NOR2_X1 i_0_37 (.ZN (n_81), .A1 (n_0_28), .A2 (n_0_354));
NOR2_X1 i_0_36 (.ZN (n_80), .A1 (n_0_28), .A2 (n_0_353));
NOR2_X1 i_0_35 (.ZN (n_79), .A1 (n_0_28), .A2 (n_0_352));
NOR2_X1 i_0_34 (.ZN (n_78), .A1 (n_0_28), .A2 (n_0_351));
NOR2_X1 i_0_33 (.ZN (n_77), .A1 (n_0_28), .A2 (n_0_350));
NOR2_X1 i_0_32 (.ZN (n_76), .A1 (n_0_28), .A2 (n_0_349));
NOR2_X1 i_0_31 (.ZN (n_75), .A1 (n_0_28), .A2 (n_0_348));
NOR2_X1 i_0_30 (.ZN (n_74), .A1 (n_0_28), .A2 (n_0_347));
NOR2_X1 i_0_29 (.ZN (n_73), .A1 (n_0_28), .A2 (n_0_346));
NOR2_X1 i_0_28 (.ZN (n_72), .A1 (n_0_28), .A2 (n_0_95));
NOR2_X1 i_0_27 (.ZN (n_71), .A1 (n_0_28), .A2 (n_0_344));
NOR2_X1 i_0_26 (.ZN (n_70), .A1 (n_0_407), .A2 (n_0_391));
OR2_X2 i_0_25 (.ZN (n_0_2), .A1 (n_0_407), .A2 (n_45));
NAND2_X1 i_0_24 (.ZN (n_0_1), .A1 (n_44), .A2 (n_45));
OAI22_X1 i_0_23 (.ZN (n_69), .A1 (n_0_60), .A2 (n_0_2), .B1 (n_0_391), .B2 (n_0_1));
NAND2_X2 i_0_22 (.ZN (n_0_0), .A1 (n_0_407), .A2 (n_45));
OAI222_X1 i_0_21 (.ZN (n_68), .A1 (n_0_28), .A2 (n_0_0), .B1 (n_0_27), .B2 (n_0_2)
    , .C1 (n_0_60), .C2 (n_0_1));
OAI222_X1 i_0_20 (.ZN (n_67), .A1 (n_0_31), .A2 (n_0_0), .B1 (n_0_388), .B2 (n_0_2)
    , .C1 (n_0_27), .C2 (n_0_1));
OAI222_X1 i_0_19 (.ZN (n_66), .A1 (n_0_365), .A2 (n_0_0), .B1 (n_0_403), .B2 (n_0_2)
    , .C1 (n_0_388), .C2 (n_0_1));
OAI222_X1 i_0_18 (.ZN (n_65), .A1 (n_0_404), .A2 (n_0_0), .B1 (n_0_386), .B2 (n_0_2)
    , .C1 (n_0_403), .C2 (n_0_1));
OAI222_X1 i_0_17 (.ZN (n_64), .A1 (n_0_363), .A2 (n_0_0), .B1 (n_0_385), .B2 (n_0_2)
    , .C1 (n_0_386), .C2 (n_0_1));
OAI222_X1 i_0_16 (.ZN (n_63), .A1 (n_0_310), .A2 (n_0_0), .B1 (n_0_384), .B2 (n_0_2)
    , .C1 (n_0_385), .C2 (n_0_1));
OAI222_X1 i_0_15 (.ZN (n_62), .A1 (n_0_361), .A2 (n_0_0), .B1 (n_0_383), .B2 (n_0_2)
    , .C1 (n_0_384), .C2 (n_0_1));
OAI222_X1 i_0_14 (.ZN (n_61), .A1 (n_0_360), .A2 (n_0_0), .B1 (n_0_382), .B2 (n_0_2)
    , .C1 (n_0_383), .C2 (n_0_1));
OAI222_X1 i_0_13 (.ZN (n_60), .A1 (n_0_359), .A2 (n_0_0), .B1 (n_0_305), .B2 (n_0_2)
    , .C1 (n_0_382), .C2 (n_0_1));
OAI222_X1 i_0_12 (.ZN (n_59), .A1 (n_0_306), .A2 (n_0_0), .B1 (n_0_380), .B2 (n_0_2)
    , .C1 (n_0_305), .C2 (n_0_1));
OAI222_X1 i_0_11 (.ZN (n_58), .A1 (n_0_357), .A2 (n_0_0), .B1 (n_0_379), .B2 (n_0_2)
    , .C1 (n_0_380), .C2 (n_0_1));
OAI222_X1 i_0_10 (.ZN (n_57), .A1 (n_0_356), .A2 (n_0_0), .B1 (n_0_378), .B2 (n_0_2)
    , .C1 (n_0_379), .C2 (n_0_1));
OAI222_X1 i_0_9 (.ZN (n_56), .A1 (n_0_355), .A2 (n_0_0), .B1 (n_0_377), .B2 (n_0_2)
    , .C1 (n_0_378), .C2 (n_0_1));
OAI222_X1 i_0_8 (.ZN (n_55), .A1 (n_0_354), .A2 (n_0_0), .B1 (n_0_376), .B2 (n_0_2)
    , .C1 (n_0_377), .C2 (n_0_1));
OAI222_X1 i_0_7 (.ZN (n_54), .A1 (n_0_353), .A2 (n_0_0), .B1 (n_0_375), .B2 (n_0_2)
    , .C1 (n_0_376), .C2 (n_0_1));
OAI222_X1 i_0_6 (.ZN (n_53), .A1 (n_0_352), .A2 (n_0_0), .B1 (n_0_374), .B2 (n_0_2)
    , .C1 (n_0_375), .C2 (n_0_1));
OAI222_X1 i_0_5 (.ZN (n_52), .A1 (n_0_351), .A2 (n_0_0), .B1 (n_0_373), .B2 (n_0_2)
    , .C1 (n_0_374), .C2 (n_0_1));
OAI222_X1 i_0_4 (.ZN (n_51), .A1 (n_0_350), .A2 (n_0_0), .B1 (n_0_372), .B2 (n_0_2)
    , .C1 (n_0_373), .C2 (n_0_1));
OAI222_X1 i_0_3 (.ZN (n_50), .A1 (n_0_349), .A2 (n_0_0), .B1 (n_0_371), .B2 (n_0_2)
    , .C1 (n_0_372), .C2 (n_0_1));
OAI222_X1 i_0_2 (.ZN (n_49), .A1 (n_0_348), .A2 (n_0_0), .B1 (n_0_370), .B2 (n_0_2)
    , .C1 (n_0_371), .C2 (n_0_1));
OAI222_X1 i_0_1 (.ZN (n_48), .A1 (n_0_347), .A2 (n_0_0), .B1 (n_0_369), .B2 (n_0_2)
    , .C1 (n_0_370), .C2 (n_0_1));
OAI222_X1 i_0_0 (.ZN (n_47), .A1 (n_0_346), .A2 (n_0_0), .B1 (n_0_92), .B2 (n_0_2)
    , .C1 (n_0_369), .C2 (n_0_1));
DLH_X1 \A_in_reg[23]  (.Q (n_46), .D (hfn_ipo_n29), .G (CTS_n38));
DLH_X1 \B_in_reg[0]  (.Q (n_45), .D (n_405), .G (CTS_n38));
DLH_X1 \B_in_reg[1]  (.Q (n_44), .D (n_406), .G (CTS_n38));
DLH_X1 \B_in_reg[2]  (.Q (n_43), .D (n_407), .G (CTS_n38));
DLH_X1 \B_in_reg[3]  (.Q (n_42), .D (n_408), .G (CTS_n38));
DLH_X1 \B_in_reg[4]  (.Q (n_41), .D (n_409), .G (CTS_n38));
DLH_X1 \B_in_reg[5]  (.Q (n_40), .D (n_410), .G (CTS_n38));
DLH_X1 \B_in_reg[6]  (.Q (n_39), .D (n_411), .G (CTS_n38));
DLH_X1 \B_in_reg[7]  (.Q (n_38), .D (n_412), .G (CTS_n38));
DLH_X1 \B_in_reg[8]  (.Q (n_37), .D (n_413), .G (CTS_n38));
DLH_X1 \B_in_reg[9]  (.Q (n_36), .D (n_414), .G (CTS_n38));
DLH_X1 \B_in_reg[10]  (.Q (n_35), .D (n_415), .G (CTS_n38));
DLH_X1 \B_in_reg[11]  (.Q (n_34), .D (n_416), .G (CTS_n38));
DLH_X1 \B_in_reg[12]  (.Q (n_33), .D (n_417), .G (CTS_n38));
DLH_X1 \B_in_reg[13]  (.Q (n_32), .D (n_418), .G (CTS_n38));
DLH_X1 \B_in_reg[14]  (.Q (n_31), .D (n_419), .G (CTS_n38));
DLH_X1 \B_in_reg[15]  (.Q (n_30), .D (n_420), .G (CTS_n38));
DLH_X1 \B_in_reg[16]  (.Q (n_29), .D (n_421), .G (CTS_n38));
DLH_X1 \B_in_reg[17]  (.Q (n_28), .D (n_422), .G (CTS_n38));
DLH_X1 \B_in_reg[18]  (.Q (n_27), .D (n_423), .G (CTS_n38));
DLH_X1 \B_in_reg[19]  (.Q (n_26), .D (n_424), .G (CTS_n38));
DLH_X1 \B_in_reg[20]  (.Q (n_25), .D (n_425), .G (CTS_n38));
DLH_X1 \B_in_reg[21]  (.Q (n_24), .D (n_426), .G (CTS_n38));
DLH_X1 \B_in_reg[22]  (.Q (n_23), .D (n_427), .G (CTS_n38));
DLH_X1 \A_in_reg[0]  (.Q (n_22), .D (n_429), .G (CTS_n38));
DLH_X1 \A_in_reg[1]  (.Q (n_21), .D (n_430), .G (CTS_n38));
DLH_X1 \A_in_reg[2]  (.Q (n_20), .D (n_431), .G (CTS_n38));
DLH_X1 \A_in_reg[3]  (.Q (n_19), .D (n_432), .G (CTS_n38));
DLH_X1 \A_in_reg[4]  (.Q (n_18), .D (n_433), .G (CTS_n38));
DLH_X1 \A_in_reg[5]  (.Q (n_17), .D (n_434), .G (CTS_n38));
DLH_X1 \A_in_reg[6]  (.Q (n_16), .D (n_435), .G (CTS_n38));
DLH_X1 \A_in_reg[7]  (.Q (n_15), .D (n_436), .G (CTS_n38));
DLH_X1 \A_in_reg[8]  (.Q (n_14), .D (n_437), .G (CTS_n38));
DLH_X1 \A_in_reg[9]  (.Q (n_13), .D (n_438), .G (CTS_n38));
DLH_X1 \A_in_reg[10]  (.Q (n_12), .D (n_439), .G (CTS_n38));
DLH_X1 \A_in_reg[11]  (.Q (n_11), .D (n_440), .G (CTS_n38));
DLH_X1 \A_in_reg[12]  (.Q (n_10), .D (n_441), .G (CTS_n38));
DLH_X1 \A_in_reg[13]  (.Q (n_9), .D (n_442), .G (CTS_n38));
DLH_X1 \A_in_reg[14]  (.Q (n_8), .D (n_443), .G (CTS_n38));
DLH_X1 \A_in_reg[15]  (.Q (n_7), .D (n_444), .G (CTS_n38));
DLH_X1 \A_in_reg[16]  (.Q (n_6), .D (n_445), .G (CTS_n38));
DLH_X1 \A_in_reg[17]  (.Q (n_5), .D (n_446), .G (CTS_n38));
DLH_X1 \A_in_reg[18]  (.Q (n_4), .D (n_447), .G (CTS_n38));
DLH_X1 \A_in_reg[19]  (.Q (n_3), .D (n_448), .G (CTS_n38));
DLH_X1 \A_in_reg[20]  (.Q (n_2), .D (n_449), .G (CTS_n38));
DLH_X1 \A_in_reg[21]  (.Q (n_1), .D (n_450), .G (CTS_n38));
DLH_X1 \A_in_reg[22]  (.Q (n_0), .D (n_451), .G (CTS_n38));
DLH_X1 \Res_reg[23]  (.Q (Res[23]), .D (n_380), .G (n_452));
DLH_X1 \Res_reg[24]  (.Q (Res[24]), .D (n_381), .G (n_452));
DLH_X1 \Res_reg[25]  (.Q (Res[25]), .D (n_382), .G (n_452));
DLH_X1 \Res_reg[26]  (.Q (Res[26]), .D (n_383), .G (n_452));
DLH_X1 \Res_reg[27]  (.Q (Res[27]), .D (n_384), .G (n_452));
DLH_X1 \Res_reg[28]  (.Q (Res[28]), .D (n_385), .G (n_452));
DLH_X1 \Res_reg[29]  (.Q (Res[29]), .D (n_386), .G (n_452));
DLH_X1 \Res_reg[30]  (.Q (Res[30]), .D (n_387), .G (n_452));
DLH_X1 \Res_reg[31]  (.Q (Res[31]), .D (n_388), .G (n_452));
DLH_X1 \Res_reg[32]  (.Q (Res[32]), .D (n_389), .G (n_452));
DLH_X1 \Res_reg[33]  (.Q (Res[33]), .D (n_390), .G (n_452));
DLH_X1 \Res_reg[34]  (.Q (Res[34]), .D (n_391), .G (n_452));
DLH_X1 \Res_reg[35]  (.Q (Res[35]), .D (n_392), .G (n_452));
DLH_X1 \Res_reg[36]  (.Q (Res[36]), .D (n_393), .G (n_452));
DLH_X1 \Res_reg[37]  (.Q (Res[37]), .D (n_394), .G (n_452));
DLH_X1 \Res_reg[38]  (.Q (Res[38]), .D (n_395), .G (n_452));
DLH_X1 \Res_reg[39]  (.Q (Res[39]), .D (n_396), .G (n_452));
DLH_X1 \Res_reg[40]  (.Q (Res[40]), .D (n_397), .G (n_452));
DLH_X1 \Res_reg[41]  (.Q (Res[41]), .D (n_398), .G (n_452));
DLH_X1 \Res_reg[42]  (.Q (Res[42]), .D (n_399), .G (n_452));
DLH_X1 \Res_reg[43]  (.Q (Res[43]), .D (n_400), .G (n_452));
DLH_X1 \Res_reg[44]  (.Q (Res[44]), .D (n_401), .G (n_452));
DLH_X1 \Res_reg[45]  (.Q (Res[45]), .D (n_402), .G (n_452));
DLH_X1 \Res_reg[46]  (.Q (Res[46]), .D (n_403), .G (n_452));
DLH_X1 \Res_reg[47]  (.Q (Res[47]), .D (n_404), .G (n_452));
datapath__0_67 i_53 (.\aggregated_res[14]  ({uc_514, uc_515, uc_516, uc_517, uc_518, 
    uc_519, uc_520, uc_521, uc_522, uc_523, uc_524, uc_525, uc_526, uc_527, uc_528, 
    uc_529, \aggregated_res[14][47] , \aggregated_res[14][46] , \aggregated_res[14][45] , 
    \aggregated_res[14][44] , \aggregated_res[14][43] , \aggregated_res[14][42] , 
    \aggregated_res[14][41] , \aggregated_res[14][40] , \aggregated_res[14][39] , 
    \aggregated_res[14][38] , \aggregated_res[14][37] , \aggregated_res[14][36] , 
    \aggregated_res[14][35] , \aggregated_res[14][34] , \aggregated_res[14][33] , 
    \aggregated_res[14][32] , \aggregated_res[14][31] , \aggregated_res[14][30] , 
    \aggregated_res[14][29] , \aggregated_res[14][28] , \aggregated_res[14][27] , 
    \aggregated_res[14][26] , \aggregated_res[14][25] , \aggregated_res[14][24] , 
    \aggregated_res[14][23] , uc_530, uc_531, uc_532, uc_533, uc_534, uc_535, uc_536, 
    uc_537, uc_538, uc_539, uc_540, uc_541, uc_542, uc_543, uc_544, uc_545, uc_546, 
    uc_547, uc_548, uc_549, uc_550, uc_551, uc_552}), .p_0 ({uc_16, uc_17, uc_18, 
    uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, 
    uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, 
    uc_41, uc_42, uc_43, uc_44, n_361, uc_45, uc_46, uc_47, uc_48, uc_49, uc_50, 
    uc_51, n_360, n_359, n_379, n_358, n_357, n_356, n_378, n_355, n_354, n_353, 
    n_352, n_351, n_350, n_349, n_348, n_347, n_346, n_345, n_344, n_343, n_342, 
    n_341, n_340, n_377, n_339, uc_52, uc_53}), .p_10 ({uc_396, uc_397, uc_398, uc_399, 
    uc_400, uc_401, uc_402, uc_403, uc_404, uc_405, uc_406, uc_407, uc_408, uc_409, 
    uc_410, uc_411, n_118, n_117, n_362, n_116, n_115, n_114, n_113, n_112, n_111, 
    n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, 
    n_99, n_98, n_97, n_96, n_95, n_94, uc_412, uc_413, uc_414, uc_415, uc_416, uc_417, 
    uc_418, uc_419, uc_420, uc_421, uc_422, uc_423, uc_424, uc_425, uc_426, uc_427, 
    uc_428, uc_429, uc_430, uc_431, uc_432, uc_433}), .p_11 ({uc_434, uc_435, uc_436, 
    uc_437, uc_438, uc_439, uc_440, uc_441, uc_442, uc_443, uc_444, uc_445, uc_446, 
    uc_447, uc_448, uc_449, n_46, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, 
    n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
    n_72, n_71, uc_450, uc_451, uc_452, uc_453, uc_454, uc_455, uc_456, uc_457, uc_458, 
    uc_459, uc_460, uc_461, uc_462, uc_463, uc_464, uc_465, uc_466, uc_467, uc_468, 
    uc_469, uc_470, uc_471, uc_472, uc_473}), .p_15 ({uc_474, uc_475, uc_476, uc_477, 
    uc_478, uc_479, uc_480, uc_481, uc_482, uc_483, uc_484, uc_485, uc_486, uc_487, 
    uc_488, uc_489, uc_490, uc_491, uc_492, uc_493, uc_494, uc_495, uc_496, uc_497, 
    uc_498, uc_499, uc_500, uc_501, uc_502, uc_503, uc_504, n_70, uc_505, uc_506, 
    uc_507, uc_508, uc_509, uc_510, uc_511, n_69, n_68, n_67, n_66, n_65, n_64, n_63, 
    n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, 
    n_49, n_48, n_47, uc_512, uc_513}), .p_1 ({uc_54, uc_55, uc_56, uc_57, uc_58, 
    uc_59, uc_60, uc_61, uc_62, uc_63, uc_64, uc_65, uc_66, uc_67, uc_68, uc_69, 
    uc_70, uc_71, uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, uc_79, uc_80, 
    n_338, uc_81, uc_82, uc_83, uc_84, uc_85, uc_86, uc_87, n_337, n_376, n_336, 
    n_335, n_375, n_334, n_333, n_332, n_331, n_330, n_329, n_328, n_327, n_326, 
    n_325, n_324, n_323, n_322, n_321, n_320, n_319, n_318, n_317, n_374, n_316, 
    uc_88, uc_89, uc_90, uc_91}), .p_2 ({uc_92, uc_93, uc_94, uc_95, uc_96, uc_97, 
    uc_98, uc_99, uc_100, uc_101, uc_102, uc_103, uc_104, uc_105, uc_106, uc_107, 
    uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, uc_114, uc_115, uc_116, n_315, 
    uc_117, uc_118, uc_119, uc_120, uc_121, uc_122, uc_123, n_314, n_313, n_312, 
    n_311, n_310, n_309, n_373, n_308, n_307, n_306, n_305, n_304, n_303, n_302, 
    n_301, n_300, n_299, n_298, n_297, n_296, n_295, n_294, n_293, n_372, n_292, 
    uc_124, uc_125, uc_126, uc_127, uc_128, uc_129}), .p_3 ({uc_130, uc_131, uc_132, 
    uc_133, uc_134, uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, uc_141, uc_142, 
    uc_143, uc_144, uc_145, uc_146, uc_147, uc_148, uc_149, uc_150, uc_151, uc_152, 
    n_291, uc_153, uc_154, uc_155, uc_156, uc_157, uc_158, uc_159, n_290, n_289, 
    n_288, n_287, n_286, n_285, n_284, n_283, n_282, n_281, n_280, n_279, n_278, 
    n_277, n_276, n_275, n_274, n_273, n_272, n_271, n_270, n_269, n_268, n_371, 
    n_267, uc_160, uc_161, uc_162, uc_163, uc_164, uc_165, uc_166, uc_167}), .p_4 ({
    uc_168, uc_169, uc_170, uc_171, uc_172, uc_173, uc_174, uc_175, uc_176, uc_177, 
    uc_178, uc_179, uc_180, uc_181, uc_182, uc_183, uc_184, uc_185, uc_186, uc_187, 
    uc_188, n_266, uc_189, uc_190, uc_191, uc_192, uc_193, uc_194, uc_195, n_265, 
    n_264, n_263, n_262, n_261, n_260, n_370, n_259, n_258, n_257, n_369, n_256, 
    n_255, n_254, n_253, n_252, n_251, n_250, n_249, n_248, n_247, n_246, n_245, 
    n_368, n_244, uc_196, uc_197, uc_198, uc_199, uc_200, uc_201, uc_202, uc_203, 
    uc_204, uc_205}), .p_5 ({uc_206, uc_207, uc_208, uc_209, uc_210, uc_211, uc_212, 
    uc_213, uc_214, uc_215, uc_216, uc_217, uc_218, uc_219, uc_220, uc_221, uc_222, 
    uc_223, uc_224, uc_225, n_243, uc_226, uc_227, uc_228, uc_229, uc_230, uc_231, 
    n_242, n_241, n_240, n_239, n_238, n_237, n_236, n_235, n_234, n_233, n_232, 
    n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, n_222, n_221, 
    n_220, n_367, n_219, uc_232, uc_233, uc_234, uc_235, uc_236, uc_237, uc_238, 
    uc_239, uc_240, uc_241, uc_242, uc_243}), .p_6 ({uc_244, uc_245, uc_246, uc_247, 
    uc_248, uc_249, uc_250, uc_251, uc_252, uc_253, uc_254, uc_255, uc_256, uc_257, 
    uc_258, uc_259, uc_260, uc_261, n_218, uc_262, uc_263, uc_264, uc_265, uc_266, 
    uc_267, n_217, n_216, n_215, n_214, n_213, n_212, n_211, n_210, n_209, n_208, 
    n_207, n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, n_197, 
    n_196, n_195, n_366, n_194, uc_268, uc_269, uc_270, uc_271, uc_272, uc_273, uc_274, 
    uc_275, uc_276, uc_277, uc_278, uc_279, uc_280, uc_281}), .p_7 ({uc_282, uc_283, 
    uc_284, uc_285, uc_286, uc_287, uc_288, uc_289, uc_290, uc_291, uc_292, uc_293, 
    uc_294, uc_295, uc_296, uc_297, uc_298, uc_299, n_193, uc_300, uc_301, uc_302, 
    uc_303, n_192, n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, 
    n_182, n_181, n_180, n_179, n_178, n_177, n_176, n_175, n_174, n_173, n_172, 
    n_171, n_170, n_365, n_169, uc_304, uc_305, uc_306, uc_307, uc_308, uc_309, uc_310, 
    uc_311, uc_312, uc_313, uc_314, uc_315, uc_316, uc_317, uc_318, uc_319}), .p_8 ({
    uc_320, uc_321, uc_322, uc_323, uc_324, uc_325, uc_326, uc_327, uc_328, uc_329, 
    uc_330, uc_331, uc_332, uc_333, uc_334, uc_335, uc_336, uc_337, n_168, uc_338, 
    uc_339, n_167, n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, 
    n_157, n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, n_147, 
    n_146, n_145, n_364, n_144, uc_340, uc_341, uc_342, uc_343, uc_344, uc_345, uc_346, 
    uc_347, uc_348, uc_349, uc_350, uc_351, uc_352, uc_353, uc_354, uc_355, uc_356, 
    uc_357}), .p_9 ({uc_358, uc_359, uc_360, uc_361, uc_362, uc_363, uc_364, uc_365, 
    uc_366, uc_367, uc_368, uc_369, uc_370, uc_371, uc_372, uc_373, uc_374, uc_375, 
    n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, 
    n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, 
    n_121, n_120, n_363, n_119, uc_376, uc_377, uc_378, uc_379, uc_380, uc_381, uc_382, 
    uc_383, uc_384, uc_385, uc_386, uc_387, uc_388, uc_389, uc_390, uc_391, uc_392, 
    uc_393, uc_394, uc_395}));
datapath__0_0 i_2 (.A_imm_2s_complement ({uc_8, uc_9, uc_10, uc_11, \A_imm_2s_complement[27] , 
    uc_12, uc_13, uc_14, \A_imm_2s_complement[23] , \A_imm_2s_complement[22] , \A_imm_2s_complement[21] , 
    \A_imm_2s_complement[20] , \A_imm_2s_complement[19] , \A_imm_2s_complement[18] , 
    \A_imm_2s_complement[17] , \A_imm_2s_complement[16] , \A_imm_2s_complement[15] , 
    \A_imm_2s_complement[14] , \A_imm_2s_complement[13] , \A_imm_2s_complement[12] , 
    \A_imm_2s_complement[11] , \A_imm_2s_complement[10] , \A_imm_2s_complement[9] , 
    \A_imm_2s_complement[8] , \A_imm_2s_complement[7] , \A_imm_2s_complement[6] , 
    \A_imm_2s_complement[5] , \A_imm_2s_complement[4] , \A_imm_2s_complement[3] , 
    \A_imm_2s_complement[2] , \A_imm_2s_complement[1] , uc_15}), .A_imm ({uc_0, uc_1, 
    uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, n_46, n_0, n_1, n_2, n_3, n_4, n_5, n_6, 
    n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, 
    n_21, n_22}));
BUF_X4 hfn_ipo_c28 (.Z (hfn_ipo_n28), .A (n_1_0__1));
CLKBUF_X3 hfn_ipo_c29 (.Z (hfn_ipo_n29), .A (n_1_0__1));
BUF_X8 spc__L1_c91 (.Z (spc__n136), .A (n_0_91));
BUF_X8 spc__L1_c89 (.Z (spc__n134), .A (n_0_218));
CLKBUF_X1 CTS_L1_c_tid1_57 (.Z (CTS_n_tid1_52), .A (clk_CTS_1_PP_9));
CLKBUF_X1 CTS_L1_c_tid1_56 (.Z (clk_CTS_1_PP_1), .A (clk_CTS_1_PP_9));
BUF_X4 spc__L1_c86 (.Z (spc__n131), .A (n_0_251));
CLKBUF_X2 drc_ipo_c32 (.Z (drc_ipo_n32), .A (n_0_311));
CLKBUF_X2 drc_ipo_c31 (.Z (drc_ipo_n31), .A (n_0_154));
CLKBUF_X2 drc_ipo_c30 (.Z (drc_ipo_n30), .A (n_0_187));

endmodule //boothAlgoR4

module FPU_boothAlgoR4 (Res, A, B, clk, reset, enable);

output [31:0] Res;
input [31:0] A;
input [31:0] B;
input clk;
input enable;
input reset;
wire CLOCK_slh__n154;
wire CLOCK_slh_n153;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire \M_resultTruncated[22] ;
wire \M_resultTruncated[21] ;
wire \M_resultTruncated[20] ;
wire \M_resultTruncated[19] ;
wire \M_resultTruncated[18] ;
wire \M_resultTruncated[17] ;
wire \M_resultTruncated[16] ;
wire \M_resultTruncated[15] ;
wire \M_resultTruncated[14] ;
wire \M_resultTruncated[13] ;
wire \M_resultTruncated[12] ;
wire \M_resultTruncated[11] ;
wire \M_resultTruncated[10] ;
wire \M_resultTruncated[9] ;
wire \M_resultTruncated[8] ;
wire \M_resultTruncated[7] ;
wire \M_resultTruncated[6] ;
wire \M_resultTruncated[5] ;
wire \M_resultTruncated[4] ;
wire \M_resultTruncated[3] ;
wire \M_resultTruncated[2] ;
wire \M_resultTruncated[1] ;
wire \M_resultTruncated[0] ;
wire \EA[7] ;
wire \EA[6] ;
wire \EA[5] ;
wire \EA[4] ;
wire \EA[3] ;
wire \EA[2] ;
wire \EA[1] ;
wire \EA[0] ;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire \EB[7] ;
wire \EB[6] ;
wire \EB[5] ;
wire \EB[4] ;
wire \EB[3] ;
wire \EB[2] ;
wire \EB[1] ;
wire \EB[0] ;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire A_reg;
wire B_reg;
wire n_0_1_2;
wire n_0_1_3;
wire n_0_1_4;
wire n_0_1_5;
wire n_0_1_6;
wire n_0_1_7;
wire n_0_1_8;
wire n_0_1_9;
wire n_0_1_10;
wire n_0_1_11;
wire n_0_1_12;
wire n_0_1_13;
wire n_0_1_14;
wire n_0_1_15;
wire n_0_1_22;
wire n_0_1_16;
wire n_0_1_23;
wire n_0_1_17;
wire n_0_1_24;
wire n_0_1_18;
wire n_0_1_25;
wire n_0_1_19;
wire n_0_1_26;
wire n_0_1_20;
wire n_0_1_27;
wire n_0_1_21;
wire n_0_1_0;
wire n_0_1_1;
wire n_0_72;
wire n_0_1_32;
wire n_0_73;
wire n_0_1_33;
wire n_0_74;
wire n_0_1_34;
wire n_0_75;
wire n_0_1_35;
wire n_0_76;
wire n_0_1_36;
wire n_0_77;
wire n_0_1_37;
wire n_0_78;
wire n_0_1_38;
wire n_0_79;
wire n_0_1_39;
wire n_0_80;
wire n_0_1_40;
wire n_0_81;
wire n_0_1_41;
wire n_0_82;
wire n_0_1_42;
wire n_0_83;
wire n_0_1_43;
wire n_0_84;
wire n_0_1_44;
wire n_0_85;
wire n_0_1_45;
wire n_0_86;
wire n_0_1_46;
wire n_0_87;
wire n_0_1_47;
wire n_0_88;
wire n_0_1_48;
wire n_0_89;
wire n_0_1_49;
wire n_0_90;
wire n_0_1_50;
wire n_0_91;
wire n_0_1_51;
wire n_0_92;
wire n_0_1_52;
wire n_0_93;
wire n_0_1_53;
wire n_0_1_54;
wire n_0_1_55;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_1_56;
wire n_0_1_57;
wire n_0_1_58;
wire n_0_1_59;
wire n_0_1_60;
wire n_0_1_62;
wire n_0_1_64;
wire n_0_103;
wire CTS_n_tid1_15;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_1_105;
wire n_0_1_106;
wire n_0_1_107;
wire n_0_1_108;
wire n_0_1_109;
wire n_0_1_110;
wire n_0_1_111;
wire n_0_1_112;
wire n_0_1_28;
wire n_0_1_29;
wire n_0_71;
wire n_0_1_30;
wire n_0_1_31;
wire n_0_1_61;
wire n_0_1_63;
wire n_0_1_65;
wire n_0_1_66;
wire n_0_1_67;
wire n_0_1_68;
wire n_0_1_69;
wire n_0_1_70;
wire n_0_1_71;
wire n_0_1_72;
wire n_0_1_73;
wire n_0_1_74;
wire n_0_1_75;
wire n_0_1_76;
wire n_0_1_77;
wire n_0_1_78;
wire n_0_1_79;
wire n_0_1_80;
wire n_0_1_81;
wire n_0_1_82;
wire n_0_1_83;
wire n_0_1_84;
wire n_0_1_85;
wire n_0_1_86;
wire n_0_1_87;
wire n_0_1_88;
wire n_0_1_89;
wire n_0_1_90;
wire n_0_1_91;
wire n_0_1_92;
wire n_0_1_93;
wire n_0_1_94;
wire n_0_1_95;
wire n_0_1_96;
wire n_0_1_97;
wire n_0_1_98;
wire n_0_1_99;
wire n_0_1_100;
wire n_0_1_101;
wire n_0_1_102;
wire CTS_n_tid1_97;
wire n_0_102;
wire n_0_1_104;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire uc_28;
wire uc_29;
wire uc_30;
wire uc_31;
wire uc_32;
wire uc_33;
wire uc_34;
wire uc_35;
wire uc_36;
wire uc_37;
wire uc_38;
wire uc_39;
wire uc_40;
wire uc_41;
wire uc_42;
wire uc_43;
wire uc_44;
wire uc_45;
wire uc_46;
wire uc_47;
wire uc_48;
wire uc_49;
wire uc_50;
wire uc_51;
wire uc_52;
wire uc_53;
wire uc_54;
wire uc_55;
wire uc_56;
wire hfn_ipo_n10;
wire CTS_n_tid1_16;
wire CLOCK_slh__n156;
wire CLOCK_slh__n155;
wire CLOCK_slh__n162;
wire CLOCK_slh__n163;
wire CLOCK_slh__n164;
wire CLOCK_slh__n170;
wire CLOCK_slh__n171;
wire CLOCK_slh__n172;
wire CLOCK_slh__n178;
wire CLOCK_slh__n179;
wire CLOCK_slh__n180;
wire CLOCK_slh__n186;
wire CLOCK_slh__n187;
wire CLOCK_slh__n188;
wire CLOCK_slh__n192;
wire CLOCK_slh__n193;
wire CLOCK_slh__n194;
wire CLOCK_slh__n198;
wire CLOCK_slh__n199;
wire CLOCK_slh__n200;
wire CLOCK_slh__n204;
wire CLOCK_slh__n205;
wire CLOCK_slh__n206;
wire sph__n235;
wire sph__n236;


NOR2_X1 i_0_1_196 (.ZN (n_0_1_104), .A1 (B_reg), .A2 (A_reg));
AOI211_X1 i_0_1_124 (.ZN (n_0_102), .A (reset), .B (n_0_1_104), .C1 (B_reg), .C2 (A_reg));
CLKBUF_X1 CLOCK_slh__c99 (.Z (CLOCK_slh__n155), .A (CLOCK_slh__n154));
AND4_X1 i_0_1_122 (.ZN (n_0_1_102), .A1 (\EB[5] ), .A2 (\EB[4] ), .A3 (\EB[3] ), .A4 (\EB[0] ));
AND3_X1 i_0_1_121 (.ZN (n_0_1_101), .A1 (\EB[2] ), .A2 (\EB[1] ), .A3 (n_0_1_102));
NAND3_X1 i_0_1_120 (.ZN (n_0_1_100), .A1 (\EB[7] ), .A2 (n_0_1_101), .A3 (\EB[6] ));
AND4_X1 i_0_1_119 (.ZN (n_0_1_99), .A1 (\EA[5] ), .A2 (\EA[4] ), .A3 (\EA[3] ), .A4 (\EA[0] ));
AND3_X1 i_0_1_118 (.ZN (n_0_1_98), .A1 (\EA[2] ), .A2 (\EA[1] ), .A3 (n_0_1_99));
NAND3_X1 i_0_1_117 (.ZN (n_0_1_97), .A1 (\EA[7] ), .A2 (n_0_1_98), .A3 (\EA[6] ));
OR4_X1 i_0_1_116 (.ZN (n_0_1_96), .A1 (\EA[3] ), .A2 (\EA[2] ), .A3 (\EA[1] ), .A4 (\EA[0] ));
OR2_X1 i_0_1_115 (.ZN (n_0_1_95), .A1 (\EA[7] ), .A2 (\EA[6] ));
OR4_X1 i_0_1_114 (.ZN (n_0_1_94), .A1 (n_0_1_96), .A2 (n_0_1_95), .A3 (\EA[5] ), .A4 (\EA[4] ));
OR4_X1 i_0_1_113 (.ZN (n_0_1_93), .A1 (\EB[3] ), .A2 (\EB[2] ), .A3 (\EB[1] ), .A4 (\EB[0] ));
OR2_X1 i_0_1_112 (.ZN (n_0_1_92), .A1 (\EB[7] ), .A2 (\EB[6] ));
OR4_X1 i_0_1_111 (.ZN (n_0_1_91), .A1 (n_0_1_93), .A2 (n_0_1_92), .A3 (\EB[5] ), .A4 (\EB[4] ));
OAI22_X1 i_0_1_110 (.ZN (n_0_1_90), .A1 (n_0_1_100), .A2 (n_0_1_94), .B1 (n_0_1_97), .B2 (n_0_1_91));
INV_X1 i_0_1_109 (.ZN (n_0_1_89), .A (n_0_1_90));
NOR4_X1 i_0_1_108 (.ZN (n_0_1_88), .A1 (n_0_52), .A2 (n_0_53), .A3 (n_0_54), .A4 (n_0_55));
NOR4_X1 i_0_1_107 (.ZN (n_0_1_87), .A1 (n_0_48), .A2 (n_0_49), .A3 (n_0_50), .A4 (n_0_51));
NOR4_X1 i_0_1_106 (.ZN (n_0_1_86), .A1 (n_0_61), .A2 (n_0_62), .A3 (n_0_56), .A4 (n_0_59));
NOR3_X1 i_0_1_105 (.ZN (n_0_1_85), .A1 (n_0_65), .A2 (n_0_66), .A3 (n_0_69));
NOR4_X1 i_0_1_104 (.ZN (n_0_1_84), .A1 (n_0_60), .A2 (n_0_63), .A3 (n_0_57), .A4 (n_0_58));
NOR4_X1 i_0_1_103 (.ZN (n_0_1_83), .A1 (n_0_68), .A2 (n_0_70), .A3 (n_0_64), .A4 (n_0_67));
AND4_X1 i_0_1_102 (.ZN (n_0_1_82), .A1 (n_0_1_88), .A2 (n_0_1_87), .A3 (n_0_1_84), .A4 (n_0_1_83));
NAND3_X1 i_0_1_101 (.ZN (n_0_1_81), .A1 (n_0_1_86), .A2 (n_0_1_85), .A3 (n_0_1_82));
NOR4_X1 i_0_1_100 (.ZN (n_0_1_80), .A1 (n_0_29), .A2 (n_0_30), .A3 (n_0_31), .A4 (n_0_32));
NOR4_X1 i_0_1_99 (.ZN (n_0_1_79), .A1 (n_0_25), .A2 (n_0_26), .A3 (n_0_27), .A4 (n_0_28));
NOR4_X1 i_0_1_98 (.ZN (n_0_1_78), .A1 (n_0_38), .A2 (n_0_39), .A3 (n_0_33), .A4 (n_0_36));
NOR3_X1 i_0_1_97 (.ZN (n_0_1_77), .A1 (n_0_42), .A2 (n_0_43), .A3 (n_0_46));
NOR4_X1 i_0_1_96 (.ZN (n_0_1_76), .A1 (n_0_37), .A2 (n_0_40), .A3 (n_0_34), .A4 (n_0_35));
NOR4_X1 i_0_1_95 (.ZN (n_0_1_75), .A1 (n_0_45), .A2 (n_0_47), .A3 (n_0_41), .A4 (n_0_44));
AND4_X1 i_0_1_94 (.ZN (n_0_1_74), .A1 (n_0_1_80), .A2 (n_0_1_79), .A3 (n_0_1_76), .A4 (n_0_1_75));
NAND3_X1 i_0_1_93 (.ZN (n_0_1_73), .A1 (n_0_1_78), .A2 (n_0_1_77), .A3 (n_0_1_74));
NOR4_X1 i_0_1_92 (.ZN (n_0_1_72), .A1 (reset), .A2 (n_0_1_73), .A3 (n_0_1_81), .A4 (n_0_1_89));
INV_X1 i_0_1_91 (.ZN (n_0_1_71), .A (n_0_1_72));
OAI22_X1 i_0_1_90 (.ZN (n_0_1_70), .A1 (n_0_1_91), .A2 (n_0_1_81), .B1 (n_0_1_94), .B2 (n_0_1_73));
NOR2_X1 i_0_1_89 (.ZN (n_0_1_69), .A1 (reset), .A2 (n_0_1_70));
AND2_X1 i_0_1_88 (.ZN (n_0_1_68), .A1 (\EA[7] ), .A2 (\EB[7] ));
OAI221_X1 i_0_1_87 (.ZN (n_0_1_67), .A (n_0_1_68), .B1 (\EA[6] ), .B2 (n_0_1_98), .C1 (\EB[6] ), .C2 (n_0_1_101));
OR4_X1 i_0_1_86 (.ZN (n_0_1_66), .A1 (n_0_1_101), .A2 (n_0_1_98), .A3 (n_0_1_92), .A4 (n_0_1_95));
AOI22_X1 i_0_1_85 (.ZN (n_0_1_65), .A1 (n_0_1_29), .A2 (n_0_0), .B1 (n_0_24), .B2 (\M_resultTruncated[0] ));
NAND2_X1 i_0_1_84 (.ZN (n_0_1_63), .A1 (n_0_1_67), .A2 (n_0_1_66));
OAI211_X1 i_0_1_83 (.ZN (n_0_1_61), .A (n_0_1_100), .B (n_0_1_97), .C1 (n_0_1_65), .C2 (n_0_1_63));
INV_X1 i_0_1_82 (.ZN (n_0_1_31), .A (n_0_1_61));
OAI221_X1 i_0_1_81 (.ZN (n_0_1_30), .A (n_0_1_69), .B1 (n_0_1_100), .B2 (n_0_1_81)
    , .C1 (n_0_1_97), .C2 (n_0_1_73));
OAI21_X1 i_0_1_80 (.ZN (n_0_71), .A (n_0_1_71), .B1 (n_0_1_31), .B2 (n_0_1_30));
INV_X1 i_0_1_79 (.ZN (n_0_1_29), .A (n_0_24));
INV_X1 i_0_1_198 (.ZN (n_0_1_28), .A (enable));
INV_X1 i_0_1_78 (.ZN (n_0_1_112), .A (reset));
INV_X1 i_0_1_66 (.ZN (n_0_1_111), .A (n_0_1_14));
INV_X1 i_0_1_195 (.ZN (n_0_1_110), .A (n_0_1_22));
INV_X1 i_0_1_194 (.ZN (n_0_1_109), .A (n_0_1_23));
INV_X1 i_0_1_193 (.ZN (n_0_1_108), .A (n_0_1_24));
INV_X1 i_0_1_192 (.ZN (n_0_1_107), .A (n_0_1_25));
INV_X1 i_0_1_191 (.ZN (n_0_1_106), .A (n_0_1_26));
INV_X1 i_0_1_190 (.ZN (n_0_1_105), .A (n_0_1_27));
OR2_X2 i_0_1_189 (.ZN (n_0_168), .A1 (CTS_n_tid1_97), .A2 (reset));
AND2_X1 i_0_1_188 (.ZN (n_0_167), .A1 (hfn_ipo_n10), .A2 (B[30]));
AND2_X1 i_0_1_187 (.ZN (n_0_166), .A1 (hfn_ipo_n10), .A2 (B[29]));
AND2_X1 i_0_1_186 (.ZN (n_0_165), .A1 (hfn_ipo_n10), .A2 (B[28]));
AND2_X1 i_0_1_185 (.ZN (n_0_164), .A1 (hfn_ipo_n10), .A2 (B[27]));
AND2_X1 i_0_1_184 (.ZN (n_0_163), .A1 (hfn_ipo_n10), .A2 (B[26]));
AND2_X1 i_0_1_183 (.ZN (n_0_162), .A1 (hfn_ipo_n10), .A2 (B[25]));
AND2_X1 i_0_1_182 (.ZN (n_0_161), .A1 (hfn_ipo_n10), .A2 (B[24]));
AND2_X1 i_0_1_181 (.ZN (n_0_160), .A1 (hfn_ipo_n10), .A2 (B[23]));
AND2_X1 i_0_1_180 (.ZN (n_0_159), .A1 (n_0_1_112), .A2 (B[22]));
AND2_X1 i_0_1_179 (.ZN (n_0_158), .A1 (n_0_1_112), .A2 (B[21]));
AND2_X1 i_0_1_178 (.ZN (n_0_157), .A1 (n_0_1_112), .A2 (B[20]));
AND2_X1 i_0_1_177 (.ZN (n_0_156), .A1 (n_0_1_112), .A2 (B[19]));
AND2_X1 i_0_1_176 (.ZN (n_0_155), .A1 (n_0_1_112), .A2 (B[18]));
AND2_X1 i_0_1_175 (.ZN (n_0_154), .A1 (n_0_1_112), .A2 (B[17]));
AND2_X1 i_0_1_174 (.ZN (n_0_153), .A1 (n_0_1_112), .A2 (B[16]));
AND2_X1 i_0_1_173 (.ZN (n_0_152), .A1 (n_0_1_112), .A2 (B[15]));
AND2_X1 i_0_1_172 (.ZN (n_0_151), .A1 (n_0_1_112), .A2 (B[14]));
AND2_X1 i_0_1_171 (.ZN (n_0_150), .A1 (n_0_1_112), .A2 (B[13]));
AND2_X1 i_0_1_170 (.ZN (n_0_149), .A1 (n_0_1_112), .A2 (B[12]));
AND2_X1 i_0_1_169 (.ZN (n_0_148), .A1 (n_0_1_112), .A2 (B[11]));
AND2_X1 i_0_1_168 (.ZN (n_0_147), .A1 (n_0_1_112), .A2 (B[10]));
AND2_X1 i_0_1_167 (.ZN (n_0_146), .A1 (n_0_1_112), .A2 (B[9]));
AND2_X1 i_0_1_166 (.ZN (n_0_145), .A1 (n_0_1_112), .A2 (B[8]));
AND2_X1 i_0_1_165 (.ZN (n_0_144), .A1 (n_0_1_112), .A2 (B[7]));
AND2_X1 i_0_1_164 (.ZN (n_0_143), .A1 (n_0_1_112), .A2 (B[6]));
AND2_X1 i_0_1_163 (.ZN (n_0_142), .A1 (n_0_1_112), .A2 (B[5]));
AND2_X1 i_0_1_162 (.ZN (n_0_141), .A1 (n_0_1_112), .A2 (B[4]));
AND2_X1 i_0_1_161 (.ZN (n_0_140), .A1 (n_0_1_112), .A2 (B[3]));
AND2_X1 i_0_1_160 (.ZN (n_0_139), .A1 (n_0_1_112), .A2 (B[2]));
AND2_X1 i_0_1_159 (.ZN (n_0_138), .A1 (n_0_1_112), .A2 (B[1]));
AND2_X1 i_0_1_158 (.ZN (n_0_137), .A1 (n_0_1_112), .A2 (B[0]));
AND2_X1 i_0_1_157 (.ZN (n_0_136), .A1 (hfn_ipo_n10), .A2 (A[30]));
AND2_X1 i_0_1_156 (.ZN (n_0_135), .A1 (hfn_ipo_n10), .A2 (A[29]));
AND2_X1 i_0_1_155 (.ZN (n_0_134), .A1 (hfn_ipo_n10), .A2 (A[28]));
AND2_X1 i_0_1_154 (.ZN (n_0_133), .A1 (hfn_ipo_n10), .A2 (A[27]));
AND2_X1 i_0_1_153 (.ZN (n_0_132), .A1 (hfn_ipo_n10), .A2 (A[26]));
AND2_X1 i_0_1_152 (.ZN (n_0_131), .A1 (hfn_ipo_n10), .A2 (A[25]));
AND2_X1 i_0_1_151 (.ZN (n_0_130), .A1 (hfn_ipo_n10), .A2 (A[24]));
AND2_X1 i_0_1_150 (.ZN (n_0_129), .A1 (hfn_ipo_n10), .A2 (A[23]));
AND2_X1 i_0_1_149 (.ZN (n_0_128), .A1 (hfn_ipo_n10), .A2 (A[22]));
AND2_X1 i_0_1_148 (.ZN (n_0_127), .A1 (hfn_ipo_n10), .A2 (A[21]));
AND2_X1 i_0_1_147 (.ZN (n_0_126), .A1 (hfn_ipo_n10), .A2 (A[20]));
AND2_X1 i_0_1_146 (.ZN (n_0_125), .A1 (hfn_ipo_n10), .A2 (A[19]));
AND2_X1 i_0_1_145 (.ZN (n_0_124), .A1 (hfn_ipo_n10), .A2 (A[18]));
AND2_X1 i_0_1_144 (.ZN (n_0_123), .A1 (hfn_ipo_n10), .A2 (A[17]));
AND2_X1 i_0_1_143 (.ZN (n_0_122), .A1 (hfn_ipo_n10), .A2 (A[16]));
AND2_X1 i_0_1_142 (.ZN (n_0_121), .A1 (hfn_ipo_n10), .A2 (A[15]));
AND2_X1 i_0_1_141 (.ZN (n_0_120), .A1 (hfn_ipo_n10), .A2 (A[14]));
AND2_X1 i_0_1_140 (.ZN (n_0_119), .A1 (hfn_ipo_n10), .A2 (A[13]));
AND2_X1 i_0_1_139 (.ZN (n_0_118), .A1 (hfn_ipo_n10), .A2 (A[12]));
AND2_X1 i_0_1_138 (.ZN (n_0_117), .A1 (hfn_ipo_n10), .A2 (A[11]));
AND2_X1 i_0_1_137 (.ZN (n_0_116), .A1 (hfn_ipo_n10), .A2 (A[10]));
AND2_X1 i_0_1_136 (.ZN (n_0_115), .A1 (hfn_ipo_n10), .A2 (A[9]));
AND2_X1 i_0_1_135 (.ZN (n_0_114), .A1 (hfn_ipo_n10), .A2 (A[8]));
AND2_X1 i_0_1_134 (.ZN (n_0_113), .A1 (hfn_ipo_n10), .A2 (A[7]));
AND2_X1 i_0_1_133 (.ZN (n_0_112), .A1 (hfn_ipo_n10), .A2 (A[6]));
AND2_X1 i_0_1_132 (.ZN (n_0_111), .A1 (hfn_ipo_n10), .A2 (A[5]));
AND2_X1 i_0_1_131 (.ZN (n_0_110), .A1 (hfn_ipo_n10), .A2 (A[4]));
AND2_X1 i_0_1_130 (.ZN (n_0_109), .A1 (hfn_ipo_n10), .A2 (A[3]));
AND2_X1 i_0_1_129 (.ZN (n_0_108), .A1 (hfn_ipo_n10), .A2 (A[2]));
AND2_X1 i_0_1_128 (.ZN (n_0_107), .A1 (hfn_ipo_n10), .A2 (A[1]));
AND2_X1 i_0_1_127 (.ZN (n_0_106), .A1 (hfn_ipo_n10), .A2 (A[0]));
AND2_X1 i_0_1_126 (.ZN (n_0_105), .A1 (n_0_1_112), .A2 (B[31]));
OAI21_X4 i_0_1_125 (.ZN (CTS_n_tid1_16), .A (hfn_ipo_n10), .B1 (n_0_1_28), .B2 (clk));
AND2_X1 i_0_1_65 (.ZN (n_0_103), .A1 (n_0_1_112), .A2 (A[31]));
NAND3_X1 i_0_1_64 (.ZN (n_0_1_64), .A1 (n_0_1_100), .A2 (n_0_1_97), .A3 (n_0_1_67));
AOI21_X1 i_0_1_21 (.ZN (n_0_1_62), .A (n_0_1_72), .B1 (n_0_1_69), .B2 (n_0_1_64));
NAND2_X1 i_0_1_20 (.ZN (n_0_1_60), .A1 (n_0_1_69), .A2 (n_0_1_66));
NOR2_X1 i_0_1_77 (.ZN (n_0_1_59), .A1 (\EB[7] ), .A2 (\EA[7] ));
NOR2_X1 i_0_1_76 (.ZN (n_0_1_58), .A1 (n_0_1_68), .A2 (n_0_1_59));
XNOR2_X1 i_0_1_75 (.ZN (n_0_1_57), .A (n_0_1_13), .B (n_0_1_21));
XNOR2_X1 i_0_1_74 (.ZN (n_0_1_56), .A (n_0_1_58), .B (n_0_1_57));
OAI21_X1 i_0_1_73 (.ZN (n_0_101), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_56));
OAI21_X1 i_0_1_72 (.ZN (n_0_100), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_105));
OAI21_X1 i_0_1_71 (.ZN (n_0_99), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_106));
OAI21_X1 i_0_1_70 (.ZN (n_0_98), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_107));
OAI21_X1 i_0_1_69 (.ZN (n_0_97), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_108));
OAI21_X1 i_0_1_68 (.ZN (n_0_96), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_109));
OAI21_X1 i_0_1_67 (.ZN (n_0_95), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_110));
OAI21_X1 i_0_1_19 (.ZN (n_0_94), .A (n_0_1_62), .B1 (n_0_1_60), .B2 (n_0_1_111));
NOR3_X4 i_0_1_18 (.ZN (n_0_1_55), .A1 (n_0_1_29), .A2 (n_0_1_64), .A3 (n_0_1_60));
NOR3_X4 i_0_1_17 (.ZN (n_0_1_54), .A1 (n_0_1_60), .A2 (n_0_24), .A3 (n_0_1_64));
AOI22_X1 i_0_1_63 (.ZN (n_0_1_53), .A1 (\M_resultTruncated[22] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_22));
INV_X1 i_0_1_62 (.ZN (n_0_93), .A (n_0_1_53));
AOI22_X1 i_0_1_61 (.ZN (n_0_1_52), .A1 (\M_resultTruncated[21] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_21));
INV_X1 i_0_1_60 (.ZN (n_0_92), .A (n_0_1_52));
AOI22_X1 i_0_1_59 (.ZN (n_0_1_51), .A1 (\M_resultTruncated[20] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_20));
INV_X1 i_0_1_58 (.ZN (n_0_91), .A (n_0_1_51));
AOI22_X1 i_0_1_57 (.ZN (n_0_1_50), .A1 (\M_resultTruncated[19] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_19));
INV_X1 i_0_1_56 (.ZN (n_0_90), .A (n_0_1_50));
AOI22_X1 i_0_1_55 (.ZN (n_0_1_49), .A1 (\M_resultTruncated[18] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_18));
INV_X1 i_0_1_54 (.ZN (n_0_89), .A (n_0_1_49));
AOI22_X1 i_0_1_53 (.ZN (n_0_1_48), .A1 (\M_resultTruncated[17] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_17));
INV_X1 i_0_1_52 (.ZN (n_0_88), .A (n_0_1_48));
AOI22_X1 i_0_1_51 (.ZN (n_0_1_47), .A1 (\M_resultTruncated[16] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_16));
INV_X1 i_0_1_50 (.ZN (n_0_87), .A (n_0_1_47));
AOI22_X1 i_0_1_49 (.ZN (n_0_1_46), .A1 (\M_resultTruncated[15] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_15));
INV_X1 i_0_1_48 (.ZN (n_0_86), .A (n_0_1_46));
AOI22_X1 i_0_1_47 (.ZN (n_0_1_45), .A1 (\M_resultTruncated[14] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_14));
INV_X1 i_0_1_46 (.ZN (n_0_85), .A (n_0_1_45));
AOI22_X1 i_0_1_45 (.ZN (n_0_1_44), .A1 (\M_resultTruncated[13] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_13));
INV_X1 i_0_1_44 (.ZN (n_0_84), .A (n_0_1_44));
AOI22_X1 i_0_1_43 (.ZN (n_0_1_43), .A1 (\M_resultTruncated[12] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_12));
INV_X1 i_0_1_42 (.ZN (n_0_83), .A (n_0_1_43));
AOI22_X1 i_0_1_41 (.ZN (n_0_1_42), .A1 (\M_resultTruncated[11] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_11));
INV_X1 i_0_1_40 (.ZN (n_0_82), .A (n_0_1_42));
AOI22_X1 i_0_1_39 (.ZN (n_0_1_41), .A1 (\M_resultTruncated[10] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_10));
INV_X1 i_0_1_38 (.ZN (n_0_81), .A (n_0_1_41));
AOI22_X1 i_0_1_37 (.ZN (n_0_1_40), .A1 (\M_resultTruncated[9] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_9));
INV_X1 i_0_1_36 (.ZN (n_0_80), .A (n_0_1_40));
AOI22_X1 i_0_1_35 (.ZN (n_0_1_39), .A1 (\M_resultTruncated[8] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_8));
INV_X1 i_0_1_34 (.ZN (n_0_79), .A (n_0_1_39));
AOI22_X1 i_0_1_33 (.ZN (n_0_1_38), .A1 (\M_resultTruncated[7] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_7));
INV_X1 i_0_1_32 (.ZN (n_0_78), .A (n_0_1_38));
AOI22_X1 i_0_1_31 (.ZN (n_0_1_37), .A1 (\M_resultTruncated[6] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_6));
INV_X1 i_0_1_30 (.ZN (n_0_77), .A (n_0_1_37));
AOI22_X1 i_0_1_29 (.ZN (n_0_1_36), .A1 (\M_resultTruncated[5] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_5));
INV_X1 i_0_1_28 (.ZN (n_0_76), .A (n_0_1_36));
AOI22_X1 i_0_1_27 (.ZN (n_0_1_35), .A1 (\M_resultTruncated[4] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_4));
INV_X1 i_0_1_26 (.ZN (n_0_75), .A (n_0_1_35));
AOI22_X1 i_0_1_25 (.ZN (n_0_1_34), .A1 (\M_resultTruncated[3] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_3));
INV_X1 i_0_1_24 (.ZN (n_0_74), .A (n_0_1_34));
AOI22_X1 i_0_1_23 (.ZN (n_0_1_33), .A1 (\M_resultTruncated[2] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_2));
INV_X1 i_0_1_22 (.ZN (n_0_73), .A (n_0_1_33));
AOI22_X1 i_0_1_16 (.ZN (n_0_1_32), .A1 (\M_resultTruncated[1] ), .A2 (n_0_1_55), .B1 (n_0_1_54), .B2 (n_0_1));
INV_X1 i_0_1_15 (.ZN (n_0_72), .A (n_0_1_32));
OR2_X1 i_0_1_14 (.ZN (n_0_1_1), .A1 (\EB[0] ), .A2 (n_0_24));
XNOR2_X1 i_0_1_13 (.ZN (n_0_1_0), .A (\EB[0] ), .B (n_0_24));
FA_X1 i_0_1_12 (.CO (n_0_1_21), .S (n_0_1_27), .A (n_0_1_11), .B (n_0_1_12), .CI (n_0_1_20));
FA_X1 i_0_1_11 (.CO (n_0_1_20), .S (n_0_1_26), .A (n_0_1_9), .B (n_0_1_10), .CI (n_0_1_19));
FA_X1 i_0_1_10 (.CO (n_0_1_19), .S (n_0_1_25), .A (n_0_1_7), .B (n_0_1_8), .CI (n_0_1_18));
FA_X1 i_0_1_9 (.CO (n_0_1_18), .S (n_0_1_24), .A (n_0_1_5), .B (n_0_1_6), .CI (n_0_1_17));
FA_X1 i_0_1_8 (.CO (n_0_1_17), .S (n_0_1_23), .A (n_0_1_3), .B (n_0_1_4), .CI (n_0_1_16));
FA_X1 i_0_1_7 (.CO (n_0_1_16), .S (n_0_1_22), .A (n_0_1_1), .B (n_0_1_2), .CI (n_0_1_15));
HA_X1 i_0_1_6 (.CO (n_0_1_15), .S (n_0_1_14), .A (\EA[0] ), .B (n_0_1_0));
HA_X1 i_0_1_5 (.CO (n_0_1_13), .S (n_0_1_12), .A (\EB[6] ), .B (\EA[6] ));
HA_X1 i_0_1_4 (.CO (n_0_1_11), .S (n_0_1_10), .A (\EB[5] ), .B (\EA[5] ));
HA_X1 i_0_1_3 (.CO (n_0_1_9), .S (n_0_1_8), .A (\EB[4] ), .B (\EA[4] ));
HA_X1 i_0_1_2 (.CO (n_0_1_7), .S (n_0_1_6), .A (\EB[3] ), .B (\EA[3] ));
HA_X1 i_0_1_1 (.CO (n_0_1_5), .S (n_0_1_4), .A (\EB[2] ), .B (\EA[2] ));
HA_X1 i_0_1_0 (.CO (n_0_1_3), .S (n_0_1_2), .A (\EB[1] ), .B (\EA[1] ));
DLH_X1 \B_reg_reg[31]  (.Q (B_reg), .D (n_0_105), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[31]  (.Q (A_reg), .D (n_0_103), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[0]  (.Q (n_0_70), .D (n_0_137), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[1]  (.Q (n_0_69), .D (n_0_138), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[2]  (.Q (n_0_68), .D (n_0_139), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[3]  (.Q (n_0_67), .D (n_0_140), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[4]  (.Q (n_0_66), .D (n_0_141), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[5]  (.Q (n_0_65), .D (n_0_142), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[6]  (.Q (n_0_64), .D (n_0_143), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[7]  (.Q (n_0_63), .D (n_0_144), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[8]  (.Q (n_0_62), .D (n_0_145), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[9]  (.Q (n_0_61), .D (n_0_146), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[10]  (.Q (n_0_60), .D (n_0_147), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[11]  (.Q (n_0_59), .D (n_0_148), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[12]  (.Q (n_0_58), .D (n_0_149), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[13]  (.Q (n_0_57), .D (n_0_150), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[14]  (.Q (n_0_56), .D (n_0_151), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[15]  (.Q (n_0_55), .D (n_0_152), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[16]  (.Q (n_0_54), .D (n_0_153), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[17]  (.Q (n_0_53), .D (n_0_154), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[18]  (.Q (n_0_52), .D (n_0_155), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[19]  (.Q (n_0_51), .D (n_0_156), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[20]  (.Q (n_0_50), .D (n_0_157), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[21]  (.Q (n_0_49), .D (n_0_158), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[22]  (.Q (n_0_48), .D (n_0_159), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[23]  (.Q (\EB[0] ), .D (n_0_160), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[24]  (.Q (\EB[1] ), .D (n_0_161), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[25]  (.Q (\EB[2] ), .D (n_0_162), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[26]  (.Q (\EB[3] ), .D (n_0_163), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[27]  (.Q (\EB[4] ), .D (n_0_164), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[28]  (.Q (\EB[5] ), .D (n_0_165), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[29]  (.Q (\EB[6] ), .D (n_0_166), .G (CTS_n_tid1_15));
DLH_X1 \B_reg_reg[30]  (.Q (\EB[7] ), .D (n_0_167), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[0]  (.Q (n_0_47), .D (n_0_106), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[1]  (.Q (n_0_46), .D (n_0_107), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[2]  (.Q (n_0_45), .D (n_0_108), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[3]  (.Q (n_0_44), .D (n_0_109), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[4]  (.Q (n_0_43), .D (n_0_110), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[5]  (.Q (n_0_42), .D (n_0_111), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[6]  (.Q (n_0_41), .D (n_0_112), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[7]  (.Q (n_0_40), .D (n_0_113), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[8]  (.Q (n_0_39), .D (n_0_114), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[9]  (.Q (n_0_38), .D (n_0_115), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[10]  (.Q (n_0_37), .D (n_0_116), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[11]  (.Q (n_0_36), .D (n_0_117), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[12]  (.Q (n_0_35), .D (n_0_118), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[13]  (.Q (n_0_34), .D (n_0_119), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[14]  (.Q (n_0_33), .D (n_0_120), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[15]  (.Q (n_0_32), .D (n_0_121), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[16]  (.Q (n_0_31), .D (n_0_122), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[17]  (.Q (n_0_30), .D (n_0_123), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[18]  (.Q (n_0_29), .D (n_0_124), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[19]  (.Q (n_0_28), .D (n_0_125), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[20]  (.Q (n_0_27), .D (n_0_126), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[21]  (.Q (n_0_26), .D (n_0_127), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[22]  (.Q (n_0_25), .D (n_0_128), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[23]  (.Q (\EA[0] ), .D (n_0_129), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[24]  (.Q (\EA[1] ), .D (n_0_130), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[25]  (.Q (\EA[2] ), .D (n_0_131), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[26]  (.Q (\EA[3] ), .D (n_0_132), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[27]  (.Q (\EA[4] ), .D (n_0_133), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[28]  (.Q (\EA[5] ), .D (n_0_134), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[29]  (.Q (\EA[6] ), .D (n_0_135), .G (CTS_n_tid1_15));
DLH_X1 \A_reg_reg[30]  (.Q (\EA[7] ), .D (n_0_136), .G (CTS_n_tid1_15));
DLH_X1 \Res_reg[0]  (.Q (Res[0]), .D (n_0_71), .G (n_0_168));
DLH_X1 \Res_reg[1]  (.Q (Res[1]), .D (n_0_72), .G (n_0_168));
DLH_X1 \Res_reg[2]  (.Q (Res[2]), .D (n_0_73), .G (n_0_168));
DLH_X1 \Res_reg[3]  (.Q (Res[3]), .D (n_0_74), .G (n_0_168));
DLH_X1 \Res_reg[4]  (.Q (Res[4]), .D (n_0_75), .G (n_0_168));
DLH_X1 \Res_reg[5]  (.Q (Res[5]), .D (n_0_76), .G (n_0_168));
DLH_X1 \Res_reg[6]  (.Q (Res[6]), .D (n_0_77), .G (n_0_168));
DLH_X1 \Res_reg[7]  (.Q (Res[7]), .D (n_0_78), .G (n_0_168));
DLH_X1 \Res_reg[8]  (.Q (Res[8]), .D (n_0_79), .G (n_0_168));
DLH_X1 \Res_reg[9]  (.Q (Res[9]), .D (n_0_80), .G (n_0_168));
DLH_X1 \Res_reg[10]  (.Q (Res[10]), .D (n_0_81), .G (n_0_168));
DLH_X1 \Res_reg[11]  (.Q (Res[11]), .D (n_0_82), .G (n_0_168));
DLH_X1 \Res_reg[12]  (.Q (Res[12]), .D (n_0_83), .G (n_0_168));
DLH_X1 \Res_reg[13]  (.Q (Res[13]), .D (n_0_84), .G (n_0_168));
DLH_X1 \Res_reg[14]  (.Q (Res[14]), .D (n_0_85), .G (n_0_168));
DLH_X1 \Res_reg[15]  (.Q (Res[15]), .D (n_0_86), .G (n_0_168));
DLH_X1 \Res_reg[16]  (.Q (Res[16]), .D (n_0_87), .G (n_0_168));
DLH_X1 \Res_reg[17]  (.Q (Res[17]), .D (n_0_88), .G (n_0_168));
DLH_X1 \Res_reg[18]  (.Q (Res[18]), .D (n_0_89), .G (n_0_168));
DLH_X1 \Res_reg[19]  (.Q (Res[19]), .D (n_0_90), .G (n_0_168));
DLH_X1 \Res_reg[20]  (.Q (Res[20]), .D (n_0_91), .G (n_0_168));
DLH_X1 \Res_reg[21]  (.Q (Res[21]), .D (n_0_92), .G (n_0_168));
DLH_X1 \Res_reg[22]  (.Q (Res[22]), .D (n_0_93), .G (n_0_168));
DLH_X1 \Res_reg[23]  (.Q (Res[23]), .D (n_0_94), .G (n_0_168));
DLH_X1 \Res_reg[24]  (.Q (Res[24]), .D (n_0_95), .G (n_0_168));
DLH_X1 \Res_reg[25]  (.Q (Res[25]), .D (n_0_96), .G (n_0_168));
DLH_X1 \Res_reg[26]  (.Q (Res[26]), .D (n_0_97), .G (n_0_168));
DLH_X1 \Res_reg[27]  (.Q (Res[27]), .D (n_0_98), .G (n_0_168));
DLH_X1 \Res_reg[28]  (.Q (Res[28]), .D (n_0_99), .G (n_0_168));
DLH_X1 \Res_reg[29]  (.Q (Res[29]), .D (n_0_100), .G (n_0_168));
DLH_X1 \Res_reg[30]  (.Q (Res[30]), .D (n_0_101), .G (n_0_168));
DLH_X1 \Res_reg[31]  (.Q (Res[31]), .D (n_0_102), .G (n_0_168));
datapath__0_78 i_0_0 (.M_resultTruncated ({\M_resultTruncated[22] , \M_resultTruncated[21] , 
    \M_resultTruncated[20] , \M_resultTruncated[19] , \M_resultTruncated[18] , \M_resultTruncated[17] , 
    \M_resultTruncated[16] , \M_resultTruncated[15] , \M_resultTruncated[14] , \M_resultTruncated[13] , 
    \M_resultTruncated[12] , \M_resultTruncated[11] , \M_resultTruncated[10] , \M_resultTruncated[9] , 
    \M_resultTruncated[8] , \M_resultTruncated[7] , \M_resultTruncated[6] , \M_resultTruncated[5] , 
    \M_resultTruncated[4] , \M_resultTruncated[3] , \M_resultTruncated[2] , \M_resultTruncated[1] , 
    \M_resultTruncated[0] }), .M_multiplied (n_0_0), .p_0 ({n_0_23, n_0_22, n_0_21, 
    n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, 
    n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1}));
boothAlgoR4 multiplier (.Res ({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, 
    uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, n_0_24, n_0_23, n_0_22, n_0_21, 
    n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, 
    n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, 
    uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, 
    uc_27, uc_28, uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, 
    uc_38}), .clk_CTS_1_PP_1 (CTS_n_tid1_97), .A ({uc_39, uc_40, uc_41, uc_42, uc_43, 
    uc_44, uc_45, uc_46, uc_47, n_0_25, n_0_26, n_0_27, n_0_28, n_0_29, n_0_30, n_0_31, 
    n_0_32, n_0_33, n_0_34, n_0_35, n_0_36, n_0_37, n_0_38, n_0_39, n_0_40, n_0_41, 
    n_0_42, n_0_43, n_0_44, n_0_45, n_0_46, n_0_47}), .B ({uc_48, uc_49, uc_50, uc_51, 
    uc_52, uc_53, uc_54, uc_55, uc_56, n_0_48, n_0_49, n_0_50, n_0_51, n_0_52, n_0_53, 
    n_0_54, n_0_55, n_0_56, n_0_57, n_0_58, n_0_59, n_0_60, n_0_61, n_0_62, n_0_63, 
    n_0_64, n_0_65, n_0_66, n_0_67, n_0_68, n_0_69, n_0_70}), .enable (CLOCK_slh_n153)
    , .reset (reset), .clk_CTS_1_PP_9 (clk));
BUF_X4 hfn_ipo_c10 (.Z (hfn_ipo_n10), .A (n_0_1_112));
CLKBUF_X3 CTS_L2_c_tid1_17 (.Z (CTS_n_tid1_15), .A (CTS_n_tid1_16));
CLKBUF_X1 CLOCK_slh__c95 (.Z (CLOCK_slh__n154), .A (enable));
CLKBUF_X1 CLOCK_slh__c100 (.Z (CLOCK_slh__n156), .A (CLOCK_slh__n155));
CLKBUF_X1 CLOCK_slh__c101 (.Z (CLOCK_slh__n162), .A (CLOCK_slh__n156));
CLKBUF_X1 CLOCK_slh__c107 (.Z (CLOCK_slh__n163), .A (CLOCK_slh__n162));
CLKBUF_X1 CLOCK_slh__c108 (.Z (CLOCK_slh__n164), .A (CLOCK_slh__n163));
CLKBUF_X1 CLOCK_slh__c109 (.Z (CLOCK_slh__n170), .A (CLOCK_slh__n164));
CLKBUF_X1 CLOCK_slh__c115 (.Z (CLOCK_slh__n171), .A (CLOCK_slh__n170));
CLKBUF_X1 CLOCK_slh__c116 (.Z (CLOCK_slh__n172), .A (CLOCK_slh__n171));
CLKBUF_X1 CLOCK_slh__c117 (.Z (CLOCK_slh__n178), .A (CLOCK_slh__n172));
CLKBUF_X1 CLOCK_slh__c123 (.Z (CLOCK_slh__n179), .A (CLOCK_slh__n178));
CLKBUF_X1 CLOCK_slh__c124 (.Z (CLOCK_slh__n180), .A (CLOCK_slh__n179));
CLKBUF_X1 CLOCK_slh__c125 (.Z (CLOCK_slh__n186), .A (CLOCK_slh__n180));
CLKBUF_X1 CLOCK_slh__c131 (.Z (CLOCK_slh__n187), .A (CLOCK_slh__n186));
CLKBUF_X1 CLOCK_slh__c132 (.Z (CLOCK_slh__n188), .A (CLOCK_slh__n187));
CLKBUF_X1 CLOCK_slh__c133 (.Z (CLOCK_slh__n192), .A (CLOCK_slh__n188));
CLKBUF_X1 CLOCK_slh__c137 (.Z (CLOCK_slh__n193), .A (CLOCK_slh__n192));
CLKBUF_X1 CLOCK_slh__c138 (.Z (CLOCK_slh__n194), .A (CLOCK_slh__n193));
CLKBUF_X1 CLOCK_slh__c139 (.Z (CLOCK_slh__n198), .A (CLOCK_slh__n194));
CLKBUF_X1 CLOCK_slh__c143 (.Z (CLOCK_slh__n199), .A (CLOCK_slh__n198));
CLKBUF_X1 CLOCK_slh__c144 (.Z (CLOCK_slh__n200), .A (CLOCK_slh__n199));
CLKBUF_X1 CLOCK_slh__c145 (.Z (CLOCK_slh__n204), .A (CLOCK_slh__n200));
CLKBUF_X1 CLOCK_slh__c149 (.Z (CLOCK_slh__n205), .A (CLOCK_slh__n204));
CLKBUF_X1 CLOCK_slh__c150 (.Z (CLOCK_slh__n206), .A (CLOCK_slh__n205));
CLKBUF_X1 CLOCK_slh__c151 (.Z (sph__n235), .A (CLOCK_slh__n206));
CLKBUF_X1 sph__c180 (.Z (sph__n236), .A (sph__n235));
CLKBUF_X1 sph__c181 (.Z (CLOCK_slh_n153), .A (sph__n236));

endmodule //FPU_boothAlgoR4


